//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n464), .A2(KEYINPUT66), .A3(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(KEYINPUT3), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G137), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n480), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n481), .A2(new_n475), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n469), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT67), .Z(G160));
  AOI21_X1  g059(.A(new_n476), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n478), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n475), .A2(G138), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n474), .A2(new_n477), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  OR2_X1    g074(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n480), .A2(new_n497), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n496), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n485), .A2(KEYINPUT68), .A3(G126), .A4(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n474), .A2(G126), .A3(G2105), .A4(new_n477), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(new_n515), .B1(new_n512), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(G651), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n519), .A2(new_n521), .B1(new_n518), .B2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n520), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n527), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XOR2_X1   g107(.A(new_n532), .B(KEYINPUT7), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n513), .A2(new_n515), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n512), .A2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n519), .A2(new_n521), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n518), .A2(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n533), .B1(new_n540), .B2(G89), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n543));
  INV_X1    g118(.A(G51), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n525), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n541), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n545), .A2(new_n542), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(G168));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  INV_X1    g124(.A(G52), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n523), .A2(new_n549), .B1(new_n525), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n520), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n551), .A2(new_n553), .ZN(G171));
  XNOR2_X1  g129(.A(KEYINPUT73), .B(G81), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n540), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n539), .A2(new_n514), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G43), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n520), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT74), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n561), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n563), .A2(new_n556), .A3(new_n564), .A4(new_n558), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n523), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n516), .A2(new_n522), .A3(KEYINPUT76), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(G91), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n516), .A2(G65), .ZN(new_n577));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n520), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  XNOR2_X1  g157(.A(KEYINPUT75), .B(KEYINPUT9), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n522), .A2(G53), .A3(G543), .A4(new_n583), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n522), .A2(G53), .A3(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n582), .A2(new_n587), .ZN(G299));
  INV_X1    g163(.A(G171), .ZN(G301));
  INV_X1    g164(.A(G168), .ZN(G286));
  AND3_X1   g165(.A1(new_n516), .A2(new_n522), .A3(KEYINPUT76), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT76), .B1(new_n516), .B2(new_n522), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G87), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n516), .A2(G74), .ZN(new_n595));
  AOI22_X1  g170(.A1(G651), .A2(new_n595), .B1(new_n557), .B2(G49), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(G288));
  NAND2_X1  g172(.A1(new_n516), .A2(G61), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n520), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g175(.A1(G48), .A2(G543), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n522), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n593), .A2(G86), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(G85), .A2(new_n540), .B1(new_n557), .B2(G47), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n520), .B2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n593), .A2(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n536), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(new_n557), .B2(G54), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n608), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n608), .B1(new_n617), .B2(G868), .ZN(G321));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(G299), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G168), .B2(new_n620), .ZN(G280));
  XNOR2_X1  g197(.A(G280), .B(KEYINPUT77), .ZN(G297));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n566), .A2(new_n620), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n616), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n620), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g204(.A(G123), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n475), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI22_X1  g207(.A1(new_n486), .A2(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(G135), .B2(new_n478), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT78), .Z(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n464), .A2(new_n480), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT13), .B(G2100), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT81), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n645), .B(new_n651), .Z(new_n652));
  XOR2_X1   g227(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT80), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(G401));
  XOR2_X1   g235(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  INV_X1    g243(.A(new_n661), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n668), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2096), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n679), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n681), .B(new_n684), .C1(new_n676), .C2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G229));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G22), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G166), .B2(new_n693), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G1971), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n693), .A2(G6), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G305), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n695), .A2(G1971), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n696), .A2(new_n701), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n594), .A2(new_n596), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(new_n693), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n693), .B2(G23), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT87), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT33), .B(G1976), .Z(new_n709));
  AOI21_X1  g284(.A(new_n704), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n707), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n709), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n710), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  MUX2_X1   g291(.A(G24), .B(G290), .S(G16), .Z(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT85), .B(G1986), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n478), .A2(G131), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n475), .A2(G107), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n722));
  INV_X1    g297(.A(G119), .ZN(new_n723));
  OAI221_X1 g298(.A(new_n720), .B1(new_n721), .B2(new_n722), .C1(new_n723), .C2(new_n486), .ZN(new_n724));
  MUX2_X1   g299(.A(G25), .B(new_n724), .S(G29), .Z(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n725), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n719), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n716), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n711), .B1(new_n710), .B2(new_n715), .ZN(new_n731));
  OAI21_X1  g306(.A(KEYINPUT36), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n710), .A2(new_n715), .ZN(new_n733));
  INV_X1    g308(.A(new_n711), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n735), .A2(new_n736), .A3(new_n716), .A4(new_n729), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n567), .A2(new_n693), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n693), .B2(G19), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G1341), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(G1341), .ZN(new_n743));
  INV_X1    g318(.A(G29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G35), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G162), .B2(new_n744), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT29), .Z(new_n747));
  INV_X1    g322(.A(G2090), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n742), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n617), .A2(new_n693), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G4), .B2(new_n693), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT95), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G16), .B2(G21), .ZN(new_n756));
  NAND2_X1  g331(.A1(G168), .A2(G16), .ZN(new_n757));
  MUX2_X1   g332(.A(new_n755), .B(new_n756), .S(new_n757), .Z(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n754), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n693), .A2(G20), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT23), .ZN(new_n763));
  INV_X1    g338(.A(G299), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n693), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n752), .B2(new_n753), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n744), .A2(G32), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n464), .A2(G105), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n487), .A2(G129), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n773), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n478), .A2(G141), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT92), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n770), .B1(new_n781), .B2(new_n744), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT27), .B(G1996), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(new_n784), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n744), .A2(G26), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n487), .A2(G128), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n478), .A2(G140), .ZN(new_n792));
  OR2_X1    g367(.A1(G104), .A2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n790), .B1(new_n796), .B2(new_n744), .ZN(new_n797));
  INV_X1    g372(.A(G2067), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n635), .A2(new_n744), .ZN(new_n800));
  INV_X1    g375(.A(G28), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT30), .ZN(new_n802));
  AOI21_X1  g377(.A(G29), .B1(new_n801), .B2(KEYINPUT30), .ZN(new_n803));
  OR2_X1    g378(.A1(KEYINPUT31), .A2(G11), .ZN(new_n804));
  NAND2_X1  g379(.A1(KEYINPUT31), .A2(G11), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n787), .A2(new_n799), .A3(new_n800), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n747), .A2(new_n748), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT24), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(G34), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(G34), .ZN(new_n812));
  AOI21_X1  g387(.A(G29), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G160), .B2(new_n744), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT90), .B(G2084), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n744), .A2(G33), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT89), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT25), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n478), .A2(G139), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(new_n475), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n819), .B1(new_n826), .B2(G29), .ZN(new_n827));
  INV_X1    g402(.A(G2072), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT91), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n815), .A2(new_n817), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n808), .A2(new_n818), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n744), .A2(G27), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G164), .B2(new_n744), .ZN(new_n834));
  INV_X1    g409(.A(G2078), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n693), .A2(G5), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G171), .B2(new_n693), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(G1961), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n828), .B2(new_n827), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(G1961), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n807), .A2(new_n832), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n758), .A2(new_n759), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT96), .Z(new_n845));
  AND4_X1   g420(.A1(new_n750), .A2(new_n769), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n738), .A2(KEYINPUT97), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT97), .B1(new_n738), .B2(new_n846), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(G311));
  NAND2_X1  g424(.A1(new_n738), .A2(new_n846), .ZN(G150));
  NAND2_X1  g425(.A1(new_n617), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n523), .A2(new_n853), .B1(new_n525), .B2(new_n854), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(new_n520), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n562), .A2(new_n565), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n563), .A2(new_n558), .A3(new_n556), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(new_n858), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n562), .A2(new_n565), .A3(new_n859), .A4(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n852), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n868));
  AOI21_X1  g443(.A(G860), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n868), .B2(new_n867), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n859), .A2(G860), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT37), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(G145));
  INV_X1    g448(.A(new_n781), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n795), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n781), .A2(new_n796), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n509), .ZN(new_n878));
  INV_X1    g453(.A(new_n826), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n879), .A2(KEYINPUT99), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n875), .A2(G164), .A3(new_n876), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(KEYINPUT99), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n724), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n878), .A2(new_n880), .A3(new_n881), .A4(new_n884), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n478), .A2(G142), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n891));
  INV_X1    g466(.A(G118), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n890), .A2(new_n891), .B1(new_n892), .B2(G2105), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n891), .B2(new_n890), .ZN(new_n894));
  INV_X1    g469(.A(G130), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n889), .B(new_n894), .C1(new_n895), .C2(new_n486), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n638), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n888), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n886), .A2(new_n897), .A3(new_n887), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n635), .B(G160), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(G162), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  INV_X1    g481(.A(new_n904), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n899), .A2(new_n900), .A3(new_n907), .A4(new_n901), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g485(.A(new_n627), .B(new_n866), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n616), .A2(new_n764), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n611), .A2(G299), .A3(new_n615), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  INV_X1    g492(.A(new_n913), .ZN(new_n918));
  AOI21_X1  g493(.A(G299), .B1(new_n611), .B2(new_n615), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n912), .A2(KEYINPUT41), .A3(new_n913), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT102), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n914), .A2(new_n923), .A3(new_n917), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n911), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n916), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(G305), .B(G290), .ZN(new_n927));
  XNOR2_X1  g502(.A(G288), .B(G303), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n927), .B(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT42), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n930), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(new_n916), .A3(new_n925), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n933), .A3(G868), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n859), .B2(new_n620), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n931), .A2(new_n933), .A3(new_n935), .A4(G868), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(G295));
  NAND2_X1  g515(.A1(new_n939), .A2(KEYINPUT104), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n937), .A2(new_n942), .A3(new_n938), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(G331));
  NAND3_X1  g519(.A1(new_n864), .A2(G301), .A3(new_n865), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G301), .B1(new_n864), .B2(new_n865), .ZN(new_n947));
  OAI21_X1  g522(.A(G286), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(G168), .A3(new_n945), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n922), .A2(new_n948), .A3(new_n924), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G168), .B1(new_n949), .B2(new_n945), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n946), .A2(G286), .A3(new_n947), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n914), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n954), .A3(new_n929), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n906), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n929), .B1(new_n951), .B2(new_n954), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT43), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n920), .A2(new_n921), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n948), .A3(new_n950), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n929), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n955), .A3(new_n964), .A4(new_n906), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n958), .A2(new_n959), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT43), .B1(new_n956), .B2(new_n962), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT105), .B(KEYINPUT43), .C1(new_n956), .C2(new_n962), .ZN(new_n970));
  OR3_X1    g545(.A1(new_n956), .A2(KEYINPUT43), .A3(new_n957), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n966), .B1(new_n972), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n499), .A2(new_n502), .ZN(new_n975));
  INV_X1    g550(.A(new_n496), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n505), .B(KEYINPUT68), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n503), .B2(new_n508), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT108), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n979), .A2(new_n986), .A3(KEYINPUT50), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT109), .B1(new_n983), .B2(new_n982), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n469), .A2(G40), .A3(new_n479), .A4(new_n482), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(G2090), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(KEYINPUT45), .B2(new_n983), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n979), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT107), .B(G1971), .Z(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(G303), .A2(G8), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT55), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(G8), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1981), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n602), .A2(new_n603), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n516), .A2(new_n522), .A3(G86), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n522), .A2(new_n601), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(new_n600), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1006), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1005), .B1(new_n1012), .B2(new_n1004), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT49), .B(new_n1005), .C1(new_n1012), .C2(new_n1004), .ZN(new_n1016));
  INV_X1    g591(.A(new_n990), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n981), .A2(new_n1017), .A3(new_n984), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .A4(G8), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n705), .A2(G1976), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(G8), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT52), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1018), .A2(G8), .A3(new_n1020), .A4(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1019), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1005), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G288), .A2(G1976), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1019), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1018), .A2(G8), .ZN(new_n1030));
  OAI22_X1  g605(.A1(new_n1003), .A2(new_n1026), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT45), .B1(new_n981), .B2(new_n984), .ZN(new_n1032));
  INV_X1    g607(.A(new_n993), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n759), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n990), .A2(G2084), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n985), .A2(new_n989), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(G168), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G8), .ZN(new_n1038));
  AOI21_X1  g613(.A(G168), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT51), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT62), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1042), .A3(G8), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1041), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n509), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT111), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n509), .A2(new_n1051), .A3(new_n1048), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n990), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT108), .B1(new_n509), .B2(new_n974), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n980), .B(G1384), .C1(new_n503), .C2(new_n508), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT50), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n748), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1047), .B1(new_n1057), .B2(new_n998), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1003), .B1(new_n1002), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT124), .B1(new_n1059), .B2(new_n1026), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n985), .A2(new_n989), .A3(new_n1017), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT122), .B(G1961), .Z(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n996), .B2(G2078), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(G2078), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n993), .B(new_n1066), .C1(new_n1067), .C2(KEYINPUT45), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1063), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G171), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1058), .A2(new_n1002), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1026), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1003), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1060), .A2(new_n1071), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1031), .B1(new_n1046), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n982), .B1(new_n981), .B2(new_n984), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1051), .B1(new_n509), .B2(new_n1048), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1048), .ZN(new_n1080));
  AOI211_X1 g655(.A(KEYINPUT111), .B(new_n1080), .C1(new_n503), .C2(new_n508), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1017), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n766), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n581), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n576), .A2(new_n580), .A3(KEYINPUT115), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n587), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n576), .A2(new_n587), .A3(new_n580), .A4(KEYINPUT57), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1090), .B(KEYINPUT116), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n993), .A2(new_n995), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1083), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1061), .A2(new_n753), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1018), .A2(G2067), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n616), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1092), .B1(new_n1083), .B2(new_n1094), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1095), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT61), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1104));
  AOI21_X1  g679(.A(G1956), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1094), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(KEYINPUT120), .A3(new_n1095), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1067), .A2(new_n982), .B1(new_n988), .B2(new_n987), .ZN(new_n1111));
  AOI21_X1  g686(.A(G1348), .B1(new_n1111), .B2(new_n1017), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1110), .B1(new_n1112), .B2(new_n1097), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1096), .A2(KEYINPUT60), .A3(new_n1098), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1114), .A3(new_n617), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1095), .A2(KEYINPUT121), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1083), .A2(new_n1117), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1116), .A2(KEYINPUT61), .A3(new_n1107), .A4(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1109), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1018), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1018), .A2(KEYINPUT118), .A3(new_n1121), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n996), .B2(G1996), .ZN(new_n1127));
  INV_X1    g702(.A(G1996), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n993), .A2(KEYINPUT117), .A3(new_n1128), .A4(new_n995), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1130), .A2(new_n1131), .A3(KEYINPUT59), .A4(new_n567), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1096), .A2(KEYINPUT60), .A3(new_n616), .A4(new_n1098), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1125), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT118), .B1(new_n1018), .B2(new_n1121), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n566), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1139));
  OAI211_X1 g714(.A(new_n1132), .B(new_n1133), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1101), .B1(new_n1120), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n993), .A2(new_n995), .A3(new_n1066), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1063), .A2(KEYINPUT123), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1065), .B(new_n1142), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1070), .B1(new_n1146), .B2(G171), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1060), .A2(new_n1075), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1146), .A2(G171), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1069), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1148), .B1(new_n1152), .B2(G301), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1151), .A2(new_n1153), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1141), .A2(new_n1149), .A3(new_n1150), .A4(new_n1154), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1047), .B(new_n1001), .C1(new_n992), .C2(new_n998), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(G8), .A3(G168), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT113), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n999), .A2(G8), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1001), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n1074), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1002), .B1(new_n999), .B2(G8), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1165), .A2(new_n1026), .A3(KEYINPUT113), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1160), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT114), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT114), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1160), .B(new_n1169), .C1(new_n1164), .C2(new_n1166), .ZN(new_n1170));
  XNOR2_X1  g745(.A(KEYINPUT112), .B(KEYINPUT63), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1072), .A2(new_n1074), .A3(new_n1003), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1171), .B1(new_n1172), .B2(new_n1158), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1168), .A2(new_n1170), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1077), .A2(new_n1155), .A3(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n995), .A2(new_n990), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT106), .B1(new_n1177), .B2(G1996), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT106), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1176), .A2(new_n1179), .A3(new_n1128), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1181), .A2(new_n874), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n795), .B(G2067), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1183), .B1(new_n874), .B2(G1996), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1184), .A2(new_n1177), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n724), .B(new_n726), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1177), .A2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1182), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(G290), .B(G1986), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1176), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1175), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n724), .A2(new_n727), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT125), .ZN(new_n1195));
  OAI221_X1 g770(.A(new_n1195), .B1(new_n1177), .B2(new_n1184), .C1(new_n1181), .C2(new_n874), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n796), .A2(new_n798), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1177), .A2(G1986), .A3(G290), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1199), .B(KEYINPUT48), .Z(new_n1200));
  AOI22_X1  g775(.A1(new_n1198), .A2(new_n1176), .B1(new_n1188), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1176), .B1(new_n1183), .B2(new_n874), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1178), .A2(KEYINPUT46), .A3(new_n1180), .ZN(new_n1203));
  AOI21_X1  g778(.A(KEYINPUT46), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT47), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1201), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1208), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1193), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1212), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1214), .A2(KEYINPUT127), .A3(new_n1210), .A4(new_n1201), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1192), .A2(new_n1216), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g792(.A1(new_n958), .A2(new_n965), .ZN(new_n1219));
  NOR4_X1   g793(.A1(G229), .A2(new_n459), .A3(new_n659), .A4(G227), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n1219), .A2(new_n909), .A3(new_n1220), .ZN(G225));
  INV_X1    g795(.A(G225), .ZN(G308));
endmodule


