//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n550,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n578, new_n579, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G137), .ZN(new_n462));
  NAND2_X1  g037(.A1(G101), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n464), .B1(new_n468), .B2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n461), .A2(G2105), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT68), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n461), .A2(new_n467), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n469), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n482), .A2(G136), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n470), .A2(new_n472), .A3(G138), .A4(new_n467), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n461), .A2(KEYINPUT4), .A3(G138), .A4(new_n467), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n470), .A2(new_n472), .A3(G126), .A4(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(G2105), .B1(KEYINPUT69), .B2(G114), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT69), .A2(G114), .ZN(new_n496));
  OAI211_X1 g071(.A(G2104), .B(new_n494), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n500), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(G88), .B1(G62), .B2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(G166));
  NAND2_X1  g091(.A1(G63), .A2(G651), .ZN(new_n517));
  OR3_X1    g092(.A1(new_n514), .A2(KEYINPUT71), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT71), .B1(new_n514), .B2(new_n517), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(new_n514), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n506), .A2(new_n523), .A3(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n506), .A2(G51), .A3(G543), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n520), .A2(new_n522), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(G168));
  NAND2_X1  g102(.A1(G77), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G64), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n514), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n506), .A2(new_n523), .A3(G90), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n506), .A2(G52), .A3(G543), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(G171));
  NAND2_X1  g110(.A1(new_n506), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n514), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n537), .A2(G43), .B1(G651), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n506), .A2(new_n523), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G81), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  XOR2_X1   g124(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n550));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G188));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n554));
  INV_X1    g129(.A(G91), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n542), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n506), .A2(new_n523), .A3(KEYINPUT74), .A4(G91), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(KEYINPUT73), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(KEYINPUT73), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n561), .B(new_n562), .C1(new_n536), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n537), .A2(G53), .A3(new_n560), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  INV_X1    g141(.A(G78), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n514), .A2(new_n566), .B1(new_n567), .B2(new_n508), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT75), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  OAI221_X1 g145(.A(new_n570), .B1(new_n567), .B2(new_n508), .C1(new_n514), .C2(new_n566), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(G651), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n558), .A2(new_n564), .A3(new_n565), .A4(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(G299));
  OR2_X1    g152(.A1(new_n534), .A2(KEYINPUT77), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n534), .A2(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G301));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n526), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n526), .A2(new_n581), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G286));
  INV_X1    g161(.A(G166), .ZN(G303));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n500), .B1(new_n514), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT79), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n543), .A2(G87), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n537), .A2(G49), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  AOI22_X1  g168(.A1(new_n506), .A2(G48), .B1(G73), .B2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(G61), .A2(G651), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n506), .B2(G86), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n594), .A2(new_n508), .B1(new_n597), .B2(new_n514), .ZN(G305));
  NAND2_X1  g173(.A1(new_n543), .A2(G85), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n537), .A2(G47), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n500), .C2(new_n601), .ZN(G290));
  NAND3_X1  g177(.A1(new_n543), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n542), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n537), .A2(G54), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(new_n500), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G301), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(new_n612), .ZN(G284));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(new_n612), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(G299), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G280));
  INV_X1    g195(.A(G860), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n611), .B1(G559), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT80), .ZN(G148));
  NOR2_X1   g198(.A1(new_n611), .A2(G559), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(new_n612), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n546), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT81), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(KEYINPUT81), .B2(new_n625), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n479), .A2(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n482), .A2(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(new_n467), .B2(G111), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NOR2_X1   g211(.A1(new_n469), .A2(G2105), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n461), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT13), .B(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n636), .A2(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  OAI21_X1  g222(.A(KEYINPUT14), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT84), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT16), .Z(new_n652));
  XOR2_X1   g227(.A(G2443), .B(G2446), .Z(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n652), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(G14), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT85), .Z(G401));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT86), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n664), .B(KEYINPUT17), .Z(new_n669));
  OAI211_X1 g244(.A(new_n666), .B(new_n668), .C1(new_n663), .C2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT87), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n669), .A2(new_n667), .A3(new_n663), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT88), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n667), .A2(new_n662), .A3(new_n664), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2100), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT89), .B(G2096), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n681), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  AOI22_X1  g262(.A1(new_n685), .A2(KEYINPUT20), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n687), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n689), .A2(new_n681), .A3(new_n684), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n688), .B(new_n690), .C1(KEYINPUT20), .C2(new_n685), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1986), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1981), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1991), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(G229));
  XNOR2_X1  g272(.A(KEYINPUT90), .B(G29), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT30), .B(G28), .Z(new_n700));
  OAI22_X1  g275(.A1(new_n635), .A2(new_n699), .B1(G29), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G5), .A2(G16), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G171), .B2(G16), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n701), .B1(G1961), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G21), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G168), .B2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(G1966), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT31), .B(G11), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n704), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT100), .Z(new_n712));
  OR2_X1    g287(.A1(G29), .A2(G32), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT27), .B(G1996), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n479), .A2(G129), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT99), .ZN(new_n716));
  INV_X1    g291(.A(G141), .ZN(new_n717));
  OR3_X1    g292(.A1(new_n481), .A2(KEYINPUT98), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(KEYINPUT98), .B1(new_n481), .B2(new_n717), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n718), .A2(new_n719), .B1(G105), .B2(new_n637), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT26), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n713), .B(new_n714), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n703), .A2(G1961), .ZN(new_n727));
  NAND2_X1  g302(.A1(G160), .A2(G29), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT24), .B(G34), .Z(new_n729));
  OAI21_X1  g304(.A(KEYINPUT97), .B1(new_n729), .B2(new_n698), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n729), .A2(KEYINPUT97), .A3(new_n698), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G2084), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n726), .A2(new_n727), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(KEYINPUT101), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT101), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n726), .A2(new_n737), .A3(new_n727), .A4(new_n734), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n712), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n705), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n618), .B2(new_n705), .ZN(new_n743));
  INV_X1    g318(.A(G1956), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n699), .A2(G35), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n699), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT29), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G2090), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n725), .A2(G33), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT96), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT25), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n482), .A2(G139), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n753), .B(new_n754), .C1(new_n467), .C2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n750), .B1(new_n756), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(G2072), .ZN(new_n758));
  OAI22_X1  g333(.A1(new_n757), .A2(new_n758), .B1(new_n732), .B2(new_n733), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n749), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n713), .B1(new_n724), .B2(new_n725), .ZN(new_n761));
  INV_X1    g336(.A(new_n714), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n761), .A2(new_n762), .B1(G2090), .B2(new_n748), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n757), .A2(new_n758), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n760), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n699), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT95), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT28), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n479), .A2(G128), .B1(G140), .B2(new_n482), .ZN(new_n769));
  OR2_X1    g344(.A1(G104), .A2(G2105), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n770), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT93), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n774), .A2(KEYINPUT94), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(KEYINPUT94), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n768), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n705), .A2(G4), .ZN(new_n780));
  INV_X1    g355(.A(new_n611), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n705), .ZN(new_n782));
  INV_X1    g357(.A(G1348), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n546), .A2(new_n705), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n705), .B2(G19), .ZN(new_n786));
  INV_X1    g361(.A(G1341), .ZN(new_n787));
  INV_X1    g362(.A(G2078), .ZN(new_n788));
  NOR2_X1   g363(.A1(G164), .A2(new_n699), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G27), .B2(new_n699), .ZN(new_n790));
  OAI22_X1  g365(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n787), .B2(new_n786), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n779), .A2(new_n784), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n765), .A2(new_n793), .ZN(new_n794));
  AND3_X1   g369(.A1(new_n739), .A2(new_n745), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n790), .A2(new_n788), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n705), .A2(G23), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G288), .B2(G16), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT33), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G1976), .ZN(new_n803));
  INV_X1    g378(.A(G1976), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n800), .A2(new_n804), .A3(new_n801), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n705), .A2(G22), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n705), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT92), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(G1971), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n705), .A2(G6), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n503), .A2(G651), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n500), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n813));
  AOI21_X1  g388(.A(KEYINPUT70), .B1(new_n500), .B2(KEYINPUT6), .ZN(new_n814));
  OAI211_X1 g389(.A(G48), .B(new_n812), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(G73), .A2(G651), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n508), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g392(.A(G86), .B(new_n812), .C1(new_n813), .C2(new_n814), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n514), .B1(new_n818), .B2(new_n595), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n811), .B1(new_n820), .B2(new_n705), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT32), .B(G1981), .Z(new_n822));
  XOR2_X1   g397(.A(new_n821), .B(new_n822), .Z(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n809), .B2(G1971), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n806), .A2(new_n810), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT34), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n479), .A2(G119), .ZN(new_n827));
  OR2_X1    g402(.A1(G95), .A2(G2105), .ZN(new_n828));
  INV_X1    g403(.A(G107), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n469), .B1(new_n829), .B2(G2105), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n482), .A2(G131), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  MUX2_X1   g407(.A(G25), .B(new_n832), .S(new_n698), .Z(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT35), .B(G1991), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n833), .B(new_n834), .Z(new_n835));
  INV_X1    g410(.A(KEYINPUT34), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n806), .A2(new_n836), .A3(new_n810), .A4(new_n824), .ZN(new_n837));
  NOR2_X1   g412(.A1(G16), .A2(G24), .ZN(new_n838));
  XOR2_X1   g413(.A(G290), .B(KEYINPUT91), .Z(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(G16), .ZN(new_n840));
  INV_X1    g415(.A(G1986), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n826), .A2(new_n835), .A3(new_n837), .A4(new_n842), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(KEYINPUT36), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n795), .B(new_n796), .C1(new_n844), .C2(new_n845), .ZN(G150));
  NAND2_X1  g421(.A1(G150), .A2(KEYINPUT103), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n848), .A2(new_n849), .A3(new_n796), .A4(new_n795), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(G311));
  NAND2_X1  g426(.A1(new_n781), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT39), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(G80), .A2(G543), .ZN(new_n856));
  INV_X1    g431(.A(G67), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n514), .B2(new_n857), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n543), .A2(G93), .B1(G651), .B2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT104), .B(G55), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n537), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n546), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n545), .A2(new_n859), .A3(new_n861), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n855), .B(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n621), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT106), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n862), .A2(G860), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT107), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(G145));
  NAND2_X1  g447(.A1(new_n479), .A2(G130), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n482), .A2(G142), .ZN(new_n874));
  NOR2_X1   g449(.A1(G106), .A2(G2105), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(new_n467), .B2(G118), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n724), .B(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n756), .B(new_n832), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT108), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n498), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n497), .A2(new_n493), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n883), .A2(KEYINPUT108), .A3(new_n491), .A4(new_n492), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n640), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n879), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n878), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n635), .B(new_n487), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n773), .B(G160), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n888), .B(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g470(.A(G290), .B(G166), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n896), .A2(new_n820), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n820), .ZN(new_n898));
  OR3_X1    g473(.A1(new_n897), .A2(new_n898), .A3(G288), .ZN(new_n899));
  OAI21_X1  g474(.A(G288), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(KEYINPUT42), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n865), .B(new_n624), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n565), .A2(new_n572), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n904), .A2(KEYINPUT76), .A3(new_n564), .A4(new_n558), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n573), .A2(new_n574), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n905), .A2(new_n906), .A3(new_n611), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n611), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT41), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n781), .B1(new_n575), .B2(new_n576), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n905), .A2(new_n906), .A3(new_n611), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n912), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n903), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n916), .B2(new_n903), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n902), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n902), .A2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(G868), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n862), .A2(new_n612), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(G295));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n923), .ZN(G331));
  NAND2_X1  g500(.A1(G168), .A2(KEYINPUT78), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n534), .B1(new_n926), .B2(new_n582), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n526), .B1(new_n578), .B2(new_n579), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n865), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(G171), .B1(new_n583), .B2(new_n584), .ZN(new_n930));
  INV_X1    g505(.A(new_n928), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n930), .A2(new_n931), .A3(new_n863), .A4(new_n864), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n915), .A2(new_n917), .A3(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n929), .A2(new_n932), .ZN(new_n935));
  INV_X1    g510(.A(new_n916), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(KEYINPUT110), .A3(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n929), .A2(new_n932), .A3(new_n910), .A4(new_n912), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n934), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n901), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n934), .A2(new_n901), .A3(new_n940), .A4(new_n937), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n893), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT43), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT111), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n935), .A2(new_n948), .A3(new_n936), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n938), .A2(KEYINPUT112), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n935), .B1(new_n909), .B2(new_n913), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n942), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT113), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n942), .B(KEYINPUT113), .C1(new_n951), .C2(new_n952), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  INV_X1    g533(.A(new_n945), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n961), .B(KEYINPUT43), .C1(new_n943), .C2(new_n945), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n947), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n957), .A2(KEYINPUT43), .A3(new_n959), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n958), .B1(new_n943), .B2(new_n945), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT44), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n965), .A2(new_n969), .ZN(G397));
  AOI21_X1  g545(.A(G1384), .B1(new_n881), .B2(new_n884), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n971), .A2(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n462), .A2(new_n463), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n467), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT67), .B1(new_n475), .B2(G2105), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n465), .B(new_n467), .C1(new_n473), .C2(new_n474), .ZN(new_n976));
  OAI211_X1 g551(.A(G40), .B(new_n974), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n972), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n979), .A2(G1986), .A3(G290), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT48), .Z(new_n981));
  XNOR2_X1  g556(.A(new_n773), .B(G2067), .ZN(new_n982));
  INV_X1    g557(.A(G1996), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n724), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n721), .A2(G1996), .A3(new_n723), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n832), .A2(new_n834), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n832), .A2(new_n834), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n981), .B1(new_n990), .B2(new_n979), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n978), .B1(new_n724), .B2(new_n982), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n979), .B2(G1996), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n978), .A2(KEYINPUT46), .A3(new_n983), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT47), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n986), .A2(new_n989), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n773), .A2(G2067), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n978), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n991), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT126), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT121), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n1005));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n491), .A2(new_n492), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n882), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT50), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n498), .A2(new_n1010), .A3(new_n1006), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1005), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1010), .B1(new_n498), .B2(new_n1006), .ZN(new_n1013));
  OAI211_X1 g588(.A(G40), .B(G160), .C1(new_n1013), .C2(KEYINPUT114), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1004), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1961), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n977), .B1(new_n1009), .B2(new_n1005), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n498), .A2(new_n1010), .A3(new_n1006), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT114), .B1(new_n1018), .B2(new_n1013), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1019), .A3(KEYINPUT121), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(new_n1016), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n971), .A2(KEYINPUT45), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT45), .B1(new_n498), .B2(new_n1006), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n977), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1022), .B1(new_n1026), .B2(G2078), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n1006), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1022), .A2(G2078), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1021), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1031), .A2(new_n614), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n974), .A2(G40), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n971), .B2(KEYINPUT45), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n475), .A2(G2105), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n972), .A2(new_n1034), .A3(new_n1035), .A4(new_n1029), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1021), .A2(new_n1027), .A3(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(new_n614), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1003), .B1(new_n1032), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT125), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n526), .A2(G8), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT124), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1966), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1045), .B2(new_n733), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1040), .B(new_n1043), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1017), .A2(new_n1019), .A3(new_n733), .ZN(new_n1049));
  INV_X1    g624(.A(new_n977), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1024), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(new_n1028), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n708), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1047), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT125), .B1(new_n1054), .B2(new_n1042), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1048), .A2(new_n1055), .A3(KEYINPUT51), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1046), .A2(new_n1043), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n1058));
  OAI211_X1 g633(.A(KEYINPUT125), .B(new_n1058), .C1(new_n1054), .C2(new_n1042), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1039), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1037), .A2(G171), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1021), .A2(new_n1027), .A3(G301), .A4(new_n1030), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(KEYINPUT54), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G305), .A2(G1981), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT116), .B(G1981), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n820), .B2(new_n1068), .ZN(new_n1069));
  NOR4_X1   g644(.A1(new_n817), .A2(new_n819), .A3(KEYINPUT117), .A4(new_n1067), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT49), .B(new_n1065), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1065), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT49), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT117), .B1(G305), .B2(new_n1067), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n820), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(KEYINPUT118), .A3(KEYINPUT49), .A4(new_n1065), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n977), .A2(new_n1008), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(new_n1047), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1073), .A2(new_n1076), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1082), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G288), .A2(new_n804), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT52), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n804), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1082), .B(new_n1087), .C1(new_n804), .C2(G288), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1083), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G303), .A2(G8), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1971), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1026), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n1095));
  INV_X1    g670(.A(G2090), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1017), .A2(new_n1019), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1045), .B2(new_n1096), .ZN(new_n1099));
  OAI211_X1 g674(.A(G8), .B(new_n1092), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1092), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1971), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1050), .A2(new_n1011), .A3(new_n1009), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(G2090), .ZN(new_n1104));
  OAI21_X1  g679(.A(G8), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1064), .A2(new_n1089), .A3(new_n1100), .A4(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1002), .B1(new_n1061), .B2(new_n1107), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1062), .A2(KEYINPUT54), .A3(new_n1063), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1089), .A2(new_n1100), .A3(new_n1106), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1111), .A2(KEYINPUT126), .A3(new_n1039), .A4(new_n1060), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1015), .A2(new_n783), .A3(new_n1020), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1081), .A2(new_n778), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1023), .A2(new_n1025), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1103), .A2(new_n744), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n573), .A2(KEYINPUT57), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n573), .A2(KEYINPUT57), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1115), .A2(new_n781), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n1114), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT123), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1113), .A2(new_n1129), .A3(KEYINPUT60), .A4(new_n1114), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n781), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1115), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1127), .A2(KEYINPUT123), .A3(new_n611), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT58), .B(G1341), .ZN(new_n1136));
  OAI22_X1  g711(.A1(new_n1026), .A2(G1996), .B1(new_n1081), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n546), .ZN(new_n1138));
  NOR2_X1   g713(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1125), .A2(new_n1121), .A3(KEYINPUT61), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AND2_X1   g717(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1138), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT61), .B1(new_n1125), .B2(new_n1121), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1126), .B1(new_n1135), .B2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1108), .A2(new_n1112), .B1(new_n1122), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1046), .A2(new_n1047), .A3(G286), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1106), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1100), .ZN(new_n1152));
  OAI21_X1  g727(.A(G8), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n1101), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(new_n1089), .A3(new_n1150), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1089), .A2(new_n1152), .B1(new_n1155), .B2(KEYINPUT63), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1079), .B(KEYINPUT119), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1083), .A2(new_n804), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1157), .B1(new_n1158), .B2(G288), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT120), .Z(new_n1160));
  OAI21_X1  g735(.A(new_n1156), .B1(new_n1160), .B2(new_n1084), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1060), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1056), .A2(KEYINPUT62), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1032), .A2(new_n1089), .A3(new_n1100), .A4(new_n1106), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT127), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1169), .B(new_n1166), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1170));
  NOR4_X1   g745(.A1(new_n1148), .A2(new_n1161), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(G290), .B(new_n841), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n979), .B1(new_n990), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1001), .B1(new_n1171), .B2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g749(.A1(G229), .A2(new_n459), .ZN(new_n1176));
  OR2_X1    g750(.A1(new_n660), .A2(G227), .ZN(new_n1177));
  AOI21_X1  g751(.A(new_n1177), .B1(new_n892), .B2(new_n893), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n963), .A2(new_n1176), .A3(new_n1178), .ZN(G225));
  INV_X1    g753(.A(G225), .ZN(G308));
endmodule


