//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n449, new_n451, new_n452, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n569, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n639,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND2_X1  g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  INV_X1    g017(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(G234));
  NAND2_X1  g028(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n456), .A2(new_n460), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT67), .Z(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT68), .Z(G319));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(G101), .A3(new_n469), .ZN(new_n470));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n473), .A2(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT70), .ZN(G160));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(new_n468), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  MUX2_X1   g063(.A(G100), .B(G112), .S(G2105), .Z(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n486), .A2(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(G136), .B2(new_n492), .ZN(G162));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n471), .B2(new_n472), .ZN(new_n495));
  AND2_X1   g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT4), .A2(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n471), .B2(new_n472), .ZN(new_n499));
  NAND2_X1  g074(.A1(G102), .A2(G2104), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n468), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n468), .C1(new_n484), .C2(new_n485), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n497), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT71), .A3(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n513), .A2(G50), .A3(G543), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT72), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n510), .A2(new_n512), .B1(KEYINPUT6), .B2(new_n509), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n517), .A2(new_n518), .A3(G50), .A4(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT5), .B(G543), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n511), .A2(KEYINPUT71), .A3(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(KEYINPUT71), .B1(new_n511), .B2(G651), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n521), .B(new_n514), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT73), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n517), .A2(new_n526), .A3(new_n521), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n525), .A2(G88), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n521), .A2(G62), .ZN(new_n529));
  NAND2_X1  g104(.A1(G75), .A2(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n509), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n520), .A2(new_n528), .A3(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND3_X1  g109(.A1(new_n513), .A2(G543), .A3(new_n514), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n517), .A2(new_n537), .A3(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G51), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n525), .A2(G89), .A3(new_n527), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n540), .A2(new_n545), .A3(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  AND4_X1   g123(.A1(new_n537), .A2(new_n513), .A3(G543), .A4(new_n514), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n537), .B1(new_n517), .B2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(G52), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n525), .A2(G90), .A3(new_n527), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n509), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n551), .A2(new_n552), .A3(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  NAND3_X1  g132(.A1(new_n525), .A2(G81), .A3(new_n527), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(new_n521), .ZN(new_n560));
  INV_X1    g135(.A(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n549), .A2(new_n550), .ZN(new_n564));
  INV_X1    g139(.A(G43), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n558), .B(new_n563), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G188));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT9), .B1(new_n535), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n517), .A2(new_n576), .A3(G53), .A4(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(G65), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(G65), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n560), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g157(.A1(G78), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n525), .A2(G91), .A3(new_n527), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n578), .A2(new_n584), .A3(new_n585), .ZN(G299));
  OAI21_X1  g161(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n587));
  INV_X1    g162(.A(G49), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n535), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n525), .A2(new_n527), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(G87), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(new_n590), .A2(G86), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n509), .ZN(new_n595));
  INV_X1    g170(.A(new_n535), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G48), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(G305));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n525), .A2(G85), .A3(new_n527), .ZN(new_n600));
  AND2_X1   g175(.A1(G72), .A2(G543), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n521), .B2(G60), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT77), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n604));
  INV_X1    g179(.A(G60), .ZN(new_n605));
  OR2_X1    g180(.A1(KEYINPUT5), .A2(G543), .ZN(new_n606));
  NAND2_X1  g181(.A1(KEYINPUT5), .A2(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n604), .B1(new_n608), .B2(new_n601), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n603), .A2(G651), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n600), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G47), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n536), .B2(new_n538), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n599), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n539), .A2(G47), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n615), .A2(KEYINPUT78), .A3(new_n600), .A4(new_n610), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G301), .A2(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n560), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n539), .A2(G54), .B1(G651), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n525), .A2(new_n527), .ZN(new_n625));
  INV_X1    g200(.A(G92), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g202(.A1(new_n525), .A2(G92), .A3(new_n527), .A4(new_n623), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n622), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT80), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n631));
  NAND4_X1  g206(.A1(new_n622), .A2(new_n627), .A3(new_n631), .A4(new_n628), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n618), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n618), .B1(new_n634), .B2(G868), .ZN(G321));
  MUX2_X1   g211(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g212(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n634), .B1(new_n639), .B2(G860), .ZN(G148));
  NAND3_X1  g215(.A1(new_n630), .A2(new_n639), .A3(new_n632), .ZN(new_n641));
  MUX2_X1   g216(.A(new_n566), .B(new_n641), .S(G868), .Z(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g218(.A1(new_n467), .A2(new_n469), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(new_n473), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(G2100), .ZN(new_n650));
  MUX2_X1   g225(.A(G99), .B(G111), .S(G2105), .Z(new_n651));
  AOI22_X1  g226(.A1(new_n492), .A2(G135), .B1(G2104), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n487), .A2(KEYINPUT81), .A3(G123), .ZN(new_n653));
  AOI21_X1  g228(.A(KEYINPUT81), .B1(new_n487), .B2(G123), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(G2096), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n649), .A2(new_n650), .A3(new_n657), .ZN(G156));
  XOR2_X1   g233(.A(KEYINPUT15), .B(G2435), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2427), .ZN(new_n661));
  INV_X1    g236(.A(G2430), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(KEYINPUT14), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT83), .ZN(new_n666));
  XOR2_X1   g241(.A(G1341), .B(G1348), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2451), .B(G2454), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT82), .ZN(new_n671));
  XOR2_X1   g246(.A(G2443), .B(G2446), .Z(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  OR2_X1    g248(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n668), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(G14), .A3(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G401));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2072), .B(G2078), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT18), .Z(new_n682));
  INV_X1    g257(.A(new_n679), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n684), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n678), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n680), .B(KEYINPUT17), .Z(new_n689));
  OAI211_X1 g264(.A(new_n687), .B(new_n688), .C1(new_n689), .C2(new_n683), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n689), .A2(new_n683), .A3(new_n678), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n682), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(new_n656), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G2100), .ZN(G227));
  XOR2_X1   g269(.A(G1971), .B(G1976), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT19), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1956), .B(G2474), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1961), .B(G1966), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT20), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n696), .A2(new_n699), .A3(new_n702), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT85), .ZN(new_n709));
  XOR2_X1   g284(.A(G1981), .B(G1986), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n707), .B(new_n711), .ZN(G229));
  NAND2_X1  g287(.A1(new_n492), .A2(G139), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT91), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT25), .ZN(new_n716));
  NAND2_X1  g291(.A1(G115), .A2(G2104), .ZN(new_n717));
  INV_X1    g292(.A(G127), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n486), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n716), .B1(G2105), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  MUX2_X1   g297(.A(G33), .B(new_n722), .S(G29), .Z(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G2072), .Z(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G5), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G171), .B2(new_n725), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n724), .B1(G1961), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n729), .A2(G32), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n644), .A2(G105), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n732));
  NAND3_X1  g307(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n731), .B(new_n734), .C1(G141), .C2(new_n492), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n487), .A2(G129), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT93), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n730), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  NAND2_X1  g317(.A1(G164), .A2(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G27), .B2(G29), .ZN(new_n744));
  INV_X1    g319(.A(G2078), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  NOR4_X1   g322(.A1(new_n741), .A2(new_n742), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(G160), .A2(G29), .ZN(new_n749));
  AND2_X1   g324(.A1(KEYINPUT24), .A2(G34), .ZN(new_n750));
  NOR2_X1   g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n729), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2084), .ZN(new_n754));
  NOR2_X1   g329(.A1(G29), .A2(G35), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G162), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT29), .ZN(new_n757));
  INV_X1    g332(.A(G2090), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n729), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  MUX2_X1   g337(.A(G104), .B(G116), .S(G2105), .Z(new_n763));
  AOI22_X1  g338(.A1(new_n487), .A2(G128), .B1(G2104), .B2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G140), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n474), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n762), .B1(new_n770), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2067), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n748), .A2(new_n754), .A3(new_n759), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n725), .A2(G20), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT23), .Z(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G299), .B2(G16), .ZN(new_n776));
  INV_X1    g351(.A(G1956), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G16), .A2(G19), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n567), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1341), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n728), .A2(new_n773), .A3(new_n778), .A4(new_n781), .ZN(new_n782));
  AND2_X1   g357(.A1(KEYINPUT30), .A2(G28), .ZN(new_n783));
  NOR2_X1   g358(.A1(KEYINPUT30), .A2(G28), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n729), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT31), .B(G11), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n785), .B(new_n786), .C1(new_n655), .C2(new_n729), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n725), .A2(G21), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G168), .B2(new_n725), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1966), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n787), .B(new_n790), .C1(G1961), .C2(new_n727), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n725), .A2(G4), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n634), .B2(new_n725), .ZN(new_n794));
  INV_X1    g369(.A(G1348), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n782), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G6), .B(G305), .S(G16), .Z(new_n798));
  XOR2_X1   g373(.A(KEYINPUT32), .B(G1981), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n725), .A2(G23), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n591), .B2(new_n725), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT33), .B(G1976), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT88), .ZN(new_n806));
  NOR2_X1   g381(.A1(G16), .A2(G22), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G166), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1971), .ZN(new_n809));
  OR3_X1    g384(.A1(new_n805), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n806), .B1(new_n805), .B2(new_n809), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G25), .A2(G29), .ZN(new_n815));
  MUX2_X1   g390(.A(G95), .B(G107), .S(G2105), .Z(new_n816));
  AOI22_X1  g391(.A1(new_n487), .A2(G119), .B1(G2104), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n492), .A2(G131), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT86), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(KEYINPUT86), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n815), .B1(new_n822), .B2(G29), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT87), .Z(new_n824));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G1991), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G290), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G16), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G16), .B2(G24), .ZN(new_n829));
  INV_X1    g404(.A(G1986), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n826), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n810), .A2(KEYINPUT34), .A3(new_n811), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n814), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(KEYINPUT36), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(KEYINPUT36), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n797), .B1(new_n838), .B2(new_n839), .ZN(G311));
  INV_X1    g415(.A(new_n797), .ZN(new_n841));
  INV_X1    g416(.A(new_n839), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n837), .ZN(G150));
  NAND3_X1  g418(.A1(new_n525), .A2(G93), .A3(new_n527), .ZN(new_n844));
  NAND2_X1  g419(.A1(G80), .A2(G543), .ZN(new_n845));
  INV_X1    g420(.A(G67), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n560), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G651), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n844), .B(new_n848), .C1(new_n564), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  AOI22_X1  g427(.A1(new_n539), .A2(G43), .B1(G651), .B2(new_n562), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n539), .A2(G55), .B1(G651), .B2(new_n847), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n853), .A2(new_n854), .A3(new_n558), .A4(new_n844), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n566), .A2(new_n850), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n634), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G860), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n864), .B(new_n865), .C1(new_n861), .C2(new_n860), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n862), .A2(new_n863), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n852), .B1(new_n866), .B2(new_n867), .ZN(G145));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n770), .A2(new_n506), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n770), .A2(new_n506), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n738), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  INV_X1    g449(.A(new_n738), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n874), .A2(new_n875), .A3(new_n870), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n722), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n875), .B1(new_n874), .B2(new_n870), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n871), .A2(new_n738), .A3(new_n872), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n878), .A2(new_n879), .A3(new_n714), .A4(new_n720), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n820), .A2(KEYINPUT99), .A3(new_n821), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT99), .B1(new_n820), .B2(new_n821), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(KEYINPUT100), .A3(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n492), .A2(G142), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(KEYINPUT98), .Z(new_n891));
  MUX2_X1   g466(.A(G106), .B(G118), .S(G2105), .Z(new_n892));
  AOI22_X1  g467(.A1(new_n487), .A2(G130), .B1(G2104), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n646), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n886), .A2(new_n888), .A3(new_n895), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n869), .B1(new_n881), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G160), .B(KEYINPUT97), .ZN(new_n901));
  XNOR2_X1  g476(.A(G162), .B(new_n655), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n881), .B2(new_n899), .ZN(new_n904));
  INV_X1    g479(.A(new_n899), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n905), .A2(KEYINPUT101), .A3(new_n877), .A4(new_n880), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n900), .A2(new_n904), .A3(new_n906), .A4(KEYINPUT102), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n881), .A2(new_n899), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n881), .A2(new_n899), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n903), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n911), .B2(new_n916), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(G395));
  NOR2_X1   g495(.A1(new_n850), .A2(G868), .ZN(new_n921));
  INV_X1    g496(.A(G299), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n922), .A2(new_n628), .A3(new_n627), .A4(new_n622), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n629), .A2(G299), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT105), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT105), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n641), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n857), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n630), .A2(KEYINPUT104), .A3(new_n639), .A4(new_n632), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n930), .B1(new_n929), .B2(new_n931), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n927), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT106), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n937), .B(new_n927), .C1(new_n933), .C2(new_n934), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  INV_X1    g514(.A(new_n924), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n629), .A2(G299), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT41), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OR3_X1    g519(.A1(new_n933), .A2(new_n934), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n936), .A2(new_n938), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT42), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT42), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n936), .A2(new_n948), .A3(new_n945), .A4(new_n938), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(G166), .A2(new_n593), .A3(new_n597), .ZN(new_n951));
  NAND2_X1  g526(.A1(G305), .A2(G303), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n614), .A2(new_n591), .A3(new_n616), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n591), .B1(new_n614), .B2(new_n616), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT107), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n953), .B(new_n958), .C1(new_n954), .C2(new_n955), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n955), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n614), .A2(new_n591), .A3(new_n616), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(new_n953), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n950), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n957), .B2(new_n959), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n947), .A2(new_n968), .A3(new_n949), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n921), .B1(new_n970), .B2(G868), .ZN(G295));
  AOI21_X1  g546(.A(new_n921), .B1(new_n970), .B2(G868), .ZN(G331));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n554), .B1(new_n539), .B2(G52), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT109), .B1(new_n974), .B2(new_n552), .ZN(new_n975));
  AND4_X1   g550(.A1(KEYINPUT109), .A2(new_n551), .A3(new_n552), .A4(new_n555), .ZN(new_n976));
  OAI21_X1  g551(.A(G168), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  NAND2_X1  g553(.A1(G301), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n974), .A2(KEYINPUT109), .A3(new_n552), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n980), .A3(G286), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n977), .A2(new_n857), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n857), .B1(new_n977), .B2(new_n981), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n942), .B(new_n943), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n984), .A2(KEYINPUT110), .B1(new_n985), .B2(new_n927), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n942), .A2(new_n943), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n977), .A2(new_n981), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n930), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n977), .A2(new_n857), .A3(new_n981), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n987), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n966), .B1(new_n986), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n989), .A2(new_n924), .A3(new_n923), .A4(new_n990), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n984), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n915), .B1(new_n996), .B2(new_n968), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT43), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n984), .A2(new_n995), .ZN(new_n999));
  AOI21_X1  g574(.A(G37), .B1(new_n999), .B2(new_n966), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n968), .ZN(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n973), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1002), .B1(new_n994), .B2(new_n997), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1002), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1000), .A2(new_n1001), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT44), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1004), .A2(new_n1008), .A3(KEYINPUT111), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n984), .A2(KEYINPUT110), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n985), .A2(new_n927), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n993), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n968), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1011), .B1(new_n1015), .B2(new_n1000), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n966), .A2(new_n984), .A3(new_n995), .ZN(new_n1017));
  AND4_X1   g592(.A1(new_n915), .A2(new_n1017), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT44), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1006), .B1(new_n1015), .B2(new_n1000), .ZN(new_n1020));
  AND4_X1   g595(.A1(new_n915), .A2(new_n1017), .A3(new_n1001), .A4(new_n1006), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n973), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1010), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1009), .A2(new_n1023), .ZN(G397));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n506), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n477), .A2(G40), .A3(new_n481), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n738), .A2(G1996), .A3(new_n1030), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n1032), .B(KEYINPUT112), .Z(new_n1033));
  NAND2_X1  g608(.A1(new_n770), .A2(G2067), .ZN(new_n1034));
  INV_X1    g609(.A(G2067), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n768), .A2(new_n1035), .A3(new_n769), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1031), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n738), .A2(new_n1031), .A3(G1996), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1033), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n822), .A2(new_n825), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1031), .B1(new_n1041), .B2(new_n1036), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1042), .A2(KEYINPUT125), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1031), .A2(G1996), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT46), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1044), .A2(KEYINPUT46), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1034), .A2(new_n875), .A3(new_n1036), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1045), .B(new_n1046), .C1(new_n1047), .C2(new_n1031), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1049));
  XNOR2_X1  g624(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n1042), .B2(KEYINPUT125), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n822), .A2(new_n825), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1030), .B1(new_n1040), .B2(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1039), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n830), .A3(new_n1030), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT127), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT48), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1054), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1043), .A2(new_n1051), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(G8), .B1(KEYINPUT114), .B2(KEYINPUT55), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1065), .B1(G303), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n531), .B1(new_n516), .B2(new_n519), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1066), .B(new_n1064), .C1(new_n1069), .C2(new_n528), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n498), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n484), .B2(new_n485), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n500), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1074), .A2(new_n468), .B1(new_n504), .B2(new_n503), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1384), .B1(new_n1075), .B2(new_n497), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT45), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n468), .B1(new_n478), .B2(new_n479), .ZN(new_n1078));
  INV_X1    g653(.A(G40), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n476), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1028), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1971), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n506), .A2(new_n1084), .A3(new_n1025), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1085), .A2(KEYINPUT118), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1029), .B1(KEYINPUT50), .B2(new_n1026), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(KEYINPUT118), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1083), .B1(new_n1089), .B2(G2090), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1071), .B1(new_n1090), .B2(G8), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n1093));
  OAI21_X1  g668(.A(G1981), .B1(new_n595), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n593), .A2(new_n597), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n593), .B2(new_n597), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1092), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1094), .ZN(new_n1099));
  NAND2_X1  g674(.A1(G305), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(KEYINPUT49), .A3(new_n1095), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1029), .A2(new_n1026), .ZN(new_n1102));
  INV_X1    g677(.A(G8), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1098), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n591), .A2(G1976), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT52), .ZN(new_n1108));
  INV_X1    g683(.A(G1976), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT52), .B1(G288), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1105), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1113), .A2(new_n758), .A3(new_n1080), .A4(new_n1085), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT113), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1087), .A2(new_n1116), .A3(new_n758), .A4(new_n1085), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1083), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1120));
  NAND2_X1  g695(.A1(G303), .A2(new_n1067), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1064), .ZN(new_n1122));
  NAND3_X1  g697(.A1(G303), .A2(new_n1067), .A3(new_n1065), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(KEYINPUT115), .A3(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1118), .A2(G8), .A3(new_n1120), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT116), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1124), .A2(new_n1120), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(G8), .A4(new_n1118), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n1091), .B(new_n1112), .C1(new_n1126), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n1131));
  INV_X1    g706(.A(G1966), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1080), .B1(new_n1076), .B2(KEYINPUT45), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1081), .A2(KEYINPUT119), .A3(new_n1132), .ZN(new_n1138));
  INV_X1    g713(.A(G2084), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1087), .A2(new_n1139), .A3(new_n1085), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1131), .B1(new_n1141), .B2(G286), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1137), .A2(G168), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(G8), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1131), .B1(new_n1143), .B2(G8), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT62), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(KEYINPUT51), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1148), .B(new_n1149), .C1(new_n1144), .C2(new_n1142), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1077), .A2(new_n1028), .A3(new_n745), .A4(new_n1080), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1151), .A2(new_n1152), .A3(KEYINPUT53), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT53), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1087), .A2(new_n1085), .ZN(new_n1156));
  INV_X1    g731(.A(G1961), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(G301), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1130), .A2(new_n1147), .A3(new_n1150), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT124), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1159), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1141), .A2(G286), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT51), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1144), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1146), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1162), .B1(new_n1166), .B2(new_n1149), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(new_n1130), .A4(new_n1147), .ZN(new_n1169));
  XOR2_X1   g744(.A(G299), .B(KEYINPUT57), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n1089), .A2(new_n777), .ZN(new_n1171));
  XOR2_X1   g746(.A(KEYINPUT56), .B(G2072), .Z(new_n1172));
  OR2_X1    g747(.A1(new_n1081), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1170), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1156), .A2(new_n795), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1102), .A2(new_n1035), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n629), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1171), .A2(new_n1173), .A3(new_n1170), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1174), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1178), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n1181), .B2(new_n1174), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1170), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1185), .A2(KEYINPUT61), .A3(new_n1178), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1182), .A2(new_n1186), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1175), .A2(new_n629), .A3(new_n1176), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT60), .B1(new_n1188), .B2(new_n1177), .ZN(new_n1189));
  XNOR2_X1  g764(.A(KEYINPUT58), .B(G1341), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n1081), .A2(G1996), .B1(new_n1102), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n567), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT59), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1191), .A2(new_n1194), .A3(new_n567), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n629), .A2(KEYINPUT60), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1175), .A2(new_n1176), .A3(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1189), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1179), .B1(new_n1187), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT54), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1158), .A2(KEYINPUT123), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1156), .A2(new_n1204), .A3(new_n1157), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1203), .B(new_n1205), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1202), .B1(new_n1206), .B2(G171), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1155), .A2(G301), .A3(new_n1158), .ZN(new_n1208));
  AOI22_X1  g783(.A1(new_n1201), .A2(new_n1148), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1210));
  NOR2_X1   g785(.A1(new_n1206), .A2(G171), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1210), .B1(new_n1211), .B2(new_n1159), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1200), .A2(new_n1209), .A3(new_n1130), .A4(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1161), .A2(new_n1169), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1215));
  OR2_X1    g790(.A1(new_n1215), .A2(new_n1112), .ZN(new_n1216));
  AND3_X1   g791(.A1(new_n1105), .A2(new_n1109), .A3(new_n591), .ZN(new_n1217));
  NOR2_X1   g792(.A1(G305), .A2(G1981), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1104), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1220), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1141), .A2(G8), .A3(G168), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g798(.A(KEYINPUT63), .B1(new_n1130), .B2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1112), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1071), .B1(new_n1118), .B2(G8), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT63), .ZN(new_n1227));
  NOR3_X1   g802(.A1(new_n1222), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AND2_X1   g803(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g804(.A(new_n1221), .B(KEYINPUT120), .C1(new_n1224), .C2(new_n1229), .ZN(new_n1230));
  INV_X1    g805(.A(KEYINPUT120), .ZN(new_n1231));
  INV_X1    g806(.A(new_n1091), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1225), .A2(new_n1232), .A3(new_n1223), .ZN(new_n1233));
  AOI22_X1  g808(.A1(new_n1233), .A2(new_n1227), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1234));
  OAI21_X1  g809(.A(new_n1231), .B1(new_n1234), .B2(new_n1220), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1214), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g811(.A(G290), .B(new_n830), .ZN(new_n1237));
  OAI21_X1  g812(.A(new_n1054), .B1(new_n1031), .B2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g813(.A(new_n1061), .B1(new_n1236), .B2(new_n1238), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g814(.A(new_n463), .ZN(new_n1241));
  NOR3_X1   g815(.A1(G229), .A2(new_n1241), .A3(G227), .ZN(new_n1242));
  NAND2_X1  g816(.A1(new_n676), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g817(.A(new_n1243), .B1(new_n911), .B2(new_n916), .ZN(new_n1244));
  NOR2_X1   g818(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1245));
  AND2_X1   g819(.A1(new_n1244), .A2(new_n1245), .ZN(G308));
  NAND2_X1  g820(.A1(new_n1244), .A2(new_n1245), .ZN(G225));
endmodule


