//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT69), .B(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n207), .B2(KEYINPUT22), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT24), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n217), .A2(new_n218), .A3(G183gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n211), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n218), .ZN(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(KEYINPUT64), .A2(G190gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n213), .A2(new_n215), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(KEYINPUT65), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT23), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n220), .A2(new_n226), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n220), .A2(new_n234), .A3(KEYINPUT66), .A4(new_n226), .ZN(new_n238));
  INV_X1    g037(.A(G190gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n216), .B1(new_n222), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n233), .B1(new_n240), .B2(new_n232), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n217), .A2(new_n218), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT27), .B(G183gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT28), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n212), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(KEYINPUT26), .B2(new_n227), .ZN(new_n249));
  INV_X1    g048(.A(new_n229), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n227), .A2(KEYINPUT26), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n247), .B(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n242), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT70), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT29), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n242), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G226gat), .A2(G233gat), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n258), .A2(KEYINPUT71), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n261));
  INV_X1    g060(.A(new_n259), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n253), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(new_n258), .B2(new_n259), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n202), .B(new_n210), .C1(new_n260), .C2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n210), .ZN(new_n266));
  INV_X1    g065(.A(new_n263), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n242), .A2(new_n252), .A3(new_n256), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n256), .B1(new_n242), .B2(new_n252), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT29), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n267), .B1(new_n270), .B2(new_n262), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n258), .A2(KEYINPUT71), .A3(new_n259), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n266), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n257), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n262), .A2(KEYINPUT29), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n274), .A2(new_n262), .B1(new_n253), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT72), .B1(new_n276), .B2(new_n210), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n265), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  NAND2_X1  g080(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n278), .A2(KEYINPUT73), .A3(new_n281), .ZN(new_n285));
  INV_X1    g084(.A(G155gat), .ZN(new_n286));
  INV_X1    g085(.A(G162gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G141gat), .B(G148gat), .Z(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT74), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(KEYINPUT2), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n293), .B(KEYINPUT75), .Z(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT77), .B(G148gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G141gat), .ZN(new_n298));
  INV_X1    g097(.A(G148gat), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT76), .B1(new_n299), .B2(G141gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n301));
  INV_X1    g100(.A(G141gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(G148gat), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n298), .A2(KEYINPUT78), .A3(new_n300), .A4(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT78), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(KEYINPUT77), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G148gat), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n306), .A2(new_n308), .A3(G141gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n300), .A2(new_n303), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n290), .A2(KEYINPUT79), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n290), .A2(KEYINPUT79), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n313), .A2(new_n314), .B1(KEYINPUT2), .B2(new_n289), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(new_n315), .A3(KEYINPUT80), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT80), .B1(new_n312), .B2(new_n315), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n296), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n321), .B(new_n296), .C1(new_n317), .C2(new_n318), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(G113gat), .B2(G120gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n324), .B1(G113gat), .B2(G120gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI22_X1  g126(.A1(KEYINPUT68), .A2(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(KEYINPUT68), .B2(KEYINPUT1), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT67), .B(G120gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G113gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n331), .A3(new_n326), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT81), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n322), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n333), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n296), .B(new_n338), .C1(new_n317), .C2(new_n318), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n312), .A2(new_n315), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n295), .B1(new_n344), .B2(new_n316), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n336), .A2(new_n337), .A3(new_n341), .A4(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n339), .B1(new_n345), .B2(new_n334), .ZN(new_n348));
  INV_X1    g147(.A(new_n337), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT5), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(G1gat), .B(G29gat), .Z(new_n353));
  XNOR2_X1  g152(.A(G57gat), .B(G85gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n346), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n359), .A2(KEYINPUT5), .A3(new_n337), .A4(new_n336), .ZN(new_n360));
  AND4_X1   g159(.A1(KEYINPUT6), .A2(new_n352), .A3(new_n357), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n352), .A2(new_n360), .ZN(new_n362));
  INV_X1    g161(.A(new_n357), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT6), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n352), .A2(new_n360), .A3(new_n357), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n284), .A2(new_n285), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT37), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n271), .A2(new_n266), .A3(new_n272), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n369), .A2(KEYINPUT86), .B1(new_n210), .B2(new_n276), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT86), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n271), .A2(new_n272), .A3(new_n371), .A4(new_n266), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n368), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n210), .B1(new_n260), .B2(new_n264), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n274), .A2(new_n262), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n253), .A2(new_n275), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n202), .B1(new_n377), .B2(new_n266), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT37), .B1(new_n379), .B2(new_n265), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n281), .A2(KEYINPUT38), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n373), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT87), .B1(new_n367), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n281), .ZN(new_n384));
  AOI211_X1 g183(.A(new_n283), .B(new_n384), .C1(new_n379), .C2(new_n265), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT73), .B1(new_n278), .B2(new_n281), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n381), .B1(new_n278), .B2(new_n368), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n370), .A2(new_n372), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(new_n368), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n387), .A2(new_n390), .A3(new_n391), .A4(new_n366), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n379), .A2(KEYINPUT37), .A3(new_n265), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(KEYINPUT88), .A3(new_n384), .ZN(new_n394));
  INV_X1    g193(.A(new_n380), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT88), .B1(new_n393), .B2(new_n384), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT38), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT29), .B1(new_n345), .B2(new_n321), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(new_n266), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT3), .B1(new_n266), .B2(new_n255), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(new_n345), .ZN(new_n403));
  INV_X1    g202(.A(G228gat), .ZN(new_n404));
  INV_X1    g203(.A(G233gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n401), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n407), .B1(new_n401), .B2(new_n403), .ZN(new_n410));
  INV_X1    g209(.A(G22gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT85), .ZN(new_n413));
  XOR2_X1   g212(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G50gat), .ZN(new_n415));
  XOR2_X1   g214(.A(G78gat), .B(G106gat), .Z(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n410), .ZN(new_n418));
  OAI21_X1  g217(.A(G22gat), .B1(new_n418), .B2(new_n408), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n413), .A2(new_n417), .B1(new_n419), .B2(new_n412), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n421));
  AND4_X1   g220(.A1(new_n421), .A2(new_n412), .A3(new_n419), .A4(new_n417), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n284), .A2(new_n424), .A3(new_n285), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n278), .A2(KEYINPUT30), .A3(new_n281), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n379), .A2(new_n384), .A3(new_n265), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n336), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n349), .B1(new_n430), .B2(new_n358), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(KEYINPUT39), .C1(new_n349), .C2(new_n348), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(new_n363), .C1(KEYINPUT39), .C2(new_n431), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT40), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n365), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n434), .B2(new_n433), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n423), .B1(new_n429), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n399), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n399), .A2(new_n437), .A3(KEYINPUT89), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n253), .B(new_n333), .ZN(new_n442));
  NAND2_X1  g241(.A1(G227gat), .A2(G233gat), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT34), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT34), .ZN(new_n446));
  INV_X1    g245(.A(new_n253), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(new_n333), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n253), .A2(new_n338), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n446), .B(new_n443), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G43gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(G71gat), .B(G99gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n442), .A2(new_n444), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n457), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(KEYINPUT32), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n458), .A2(KEYINPUT32), .A3(new_n455), .A4(new_n459), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT36), .ZN(new_n465));
  INV_X1    g264(.A(new_n361), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n364), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n365), .B1(new_n364), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(new_n425), .A3(new_n428), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n465), .B1(new_n471), .B2(new_n423), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n440), .A2(new_n441), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n366), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n425), .A2(new_n428), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT90), .ZN(new_n476));
  INV_X1    g275(.A(new_n423), .ZN(new_n477));
  INV_X1    g276(.A(new_n464), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT91), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(KEYINPUT35), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n480), .A2(KEYINPUT35), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n429), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n485), .A2(new_n470), .A3(new_n477), .A4(new_n478), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT35), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(G71gat), .A2(G78gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(KEYINPUT9), .ZN(new_n491));
  INV_X1    g290(.A(G64gat), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n492), .A2(G57gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(G57gat), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(G71gat), .A2(G78gat), .ZN(new_n496));
  OAI22_X1  g295(.A1(new_n491), .A2(KEYINPUT99), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n495), .B(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT21), .ZN(new_n499));
  NAND2_X1  g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G127gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(G183gat), .B(G211gat), .Z(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT16), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n507), .B2(G1gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(G1gat), .B2(new_n506), .ZN(new_n509));
  INV_X1    g308(.A(G8gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n512), .B1(KEYINPUT21), .B2(new_n498), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT100), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G155gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n514), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n505), .B(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521));
  INV_X1    g320(.A(G85gat), .ZN(new_n522));
  INV_X1    g321(.A(G92gat), .ZN(new_n523));
  AOI22_X1  g322(.A1(KEYINPUT8), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G99gat), .B(G106gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(new_n498), .ZN(new_n528));
  NAND2_X1  g327(.A1(G230gat), .A2(G233gat), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(KEYINPUT103), .Z(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT104), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n527), .A2(new_n498), .A3(KEYINPUT10), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(new_n528), .B2(KEYINPUT10), .ZN(new_n534));
  INV_X1    g333(.A(new_n530), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G120gat), .B(G148gat), .Z(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT105), .ZN(new_n539));
  XNOR2_X1  g338(.A(G176gat), .B(G204gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n539), .B(new_n540), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n532), .A2(new_n541), .A3(new_n536), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(G29gat), .ZN(new_n546));
  INV_X1    g345(.A(G36gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G43gat), .B(G50gat), .Z(new_n549));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR3_X1   g350(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n554));
  AOI211_X1 g353(.A(new_n548), .B(new_n551), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n549), .A2(new_n550), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT95), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT96), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n552), .B(KEYINPUT93), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n560), .A2(new_n554), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n548), .B1(new_n561), .B2(KEYINPUT94), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(KEYINPUT94), .B2(new_n561), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n551), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT17), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT97), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n565), .A2(KEYINPUT17), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(new_n527), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n565), .ZN(new_n571));
  AND2_X1   g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n571), .A2(new_n527), .B1(KEYINPUT41), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n574), .B(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n578));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n574), .B(new_n575), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n580), .B(KEYINPUT101), .Z(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n584), .A3(KEYINPUT102), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT102), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n586), .A3(new_n583), .ZN(new_n587));
  AOI211_X1 g386(.A(new_n518), .B(new_n545), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G169gat), .B(G197gat), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT12), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n565), .A2(new_n511), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n568), .A2(new_n512), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n567), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT18), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT98), .B1(new_n565), .B2(new_n511), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(new_n596), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n565), .A2(KEYINPUT98), .A3(new_n511), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n599), .B(KEYINPUT13), .Z(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n600), .A2(new_n601), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n595), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n612), .A2(new_n608), .A3(new_n602), .A4(new_n594), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n588), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n489), .A2(KEYINPUT106), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT106), .B1(new_n489), .B2(new_n615), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n470), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g421(.A(new_n510), .B1(new_n619), .B2(new_n429), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT16), .B(G8gat), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n618), .A2(new_n485), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT42), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(KEYINPUT42), .B2(new_n625), .ZN(G1325gat));
  OR3_X1    g426(.A1(new_n618), .A2(G15gat), .A3(new_n464), .ZN(new_n628));
  INV_X1    g427(.A(new_n465), .ZN(new_n629));
  OAI21_X1  g428(.A(G15gat), .B1(new_n618), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(G1326gat));
  NOR2_X1   g430(.A1(new_n618), .A2(new_n477), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT43), .B(G22gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(G1327gat));
  NAND2_X1  g433(.A1(new_n585), .A2(new_n587), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n635), .B1(new_n473), .B2(new_n488), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n545), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n614), .A2(new_n518), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n546), .A3(new_n620), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT45), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT108), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n399), .A2(KEYINPUT89), .A3(new_n437), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT89), .B1(new_n399), .B2(new_n437), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n471), .A2(new_n423), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n476), .A2(new_n483), .B1(new_n486), .B2(KEYINPUT35), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n643), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n473), .A2(new_n488), .A3(KEYINPUT108), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n635), .A2(KEYINPUT44), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n645), .A2(new_n647), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n649), .B1(new_n654), .B2(new_n441), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT44), .B1(new_n655), .B2(new_n635), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n639), .B(KEYINPUT107), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(G29gat), .B1(new_n659), .B2(new_n470), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n660), .ZN(G1328gat));
  NAND3_X1  g460(.A1(new_n640), .A2(new_n547), .A3(new_n429), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT46), .Z(new_n663));
  OAI21_X1  g462(.A(G36gat), .B1(new_n659), .B2(new_n485), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(G1329gat));
  NAND3_X1  g464(.A1(new_n657), .A2(new_n465), .A3(new_n658), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(G43gat), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n585), .A2(new_n587), .ZN(new_n668));
  INV_X1    g467(.A(new_n639), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n464), .A2(G43gat), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n489), .A2(new_n668), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT109), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT109), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n636), .A2(new_n673), .A3(new_n669), .A4(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n667), .A2(KEYINPUT47), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n672), .A2(new_n677), .A3(new_n674), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n672), .B2(new_n674), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI211_X1 g479(.A(KEYINPUT111), .B(KEYINPUT47), .C1(new_n680), .C2(new_n667), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT111), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n675), .A2(KEYINPUT110), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n672), .A2(new_n677), .A3(new_n674), .ZN(new_n684));
  INV_X1    g483(.A(new_n658), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n629), .B(new_n685), .C1(new_n653), .C2(new_n656), .ZN(new_n686));
  INV_X1    g485(.A(G43gat), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n683), .B(new_n684), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT47), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n682), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n676), .B1(new_n681), .B2(new_n690), .ZN(G1330gat));
  NAND2_X1  g490(.A1(new_n423), .A2(G50gat), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n637), .A2(new_n477), .A3(new_n639), .ZN(new_n693));
  OAI22_X1  g492(.A1(new_n659), .A2(new_n692), .B1(G50gat), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g494(.A1(new_n668), .A2(new_n614), .A3(new_n518), .A4(new_n638), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n650), .A2(new_n651), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n620), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT112), .B(G57gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1332gat));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n429), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT49), .B(G64gat), .Z(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n701), .B2(new_n703), .ZN(G1333gat));
  INV_X1    g503(.A(G71gat), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n697), .A2(new_n705), .A3(new_n478), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n697), .A2(new_n465), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g508(.A1(new_n697), .A2(new_n423), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g510(.A1(new_n620), .A2(new_n522), .A3(new_n545), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT115), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n611), .A2(new_n613), .A3(new_n518), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT113), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n636), .A2(KEYINPUT51), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT51), .B1(new_n636), .B2(new_n715), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n545), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n653), .B2(new_n656), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT114), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n721), .A2(new_n722), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n724), .A2(new_n725), .A3(new_n470), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n719), .B1(new_n726), .B2(new_n522), .ZN(G1336gat));
  NAND2_X1  g526(.A1(new_n636), .A2(new_n715), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n638), .B1(new_n730), .B2(new_n716), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n731), .A2(new_n523), .A3(new_n429), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n523), .B1(new_n721), .B2(new_n429), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n732), .A2(KEYINPUT52), .A3(new_n733), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n653), .A2(new_n656), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT114), .B1(new_n735), .B2(new_n720), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n429), .A3(new_n723), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n732), .B1(new_n737), .B2(G92gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(G1337gat));
  AOI21_X1  g539(.A(G99gat), .B1(new_n731), .B2(new_n478), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n724), .A2(new_n725), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n465), .A2(G99gat), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(G1338gat));
  NAND2_X1  g543(.A1(new_n721), .A2(new_n423), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G106gat), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n477), .A2(G106gat), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n545), .B(new_n749), .C1(new_n717), .C2(new_n718), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n748), .ZN(new_n752));
  INV_X1    g551(.A(G106gat), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n721), .B2(new_n423), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT116), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n750), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n736), .A2(new_n423), .A3(new_n723), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(new_n758), .B2(G106gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n756), .B1(new_n759), .B2(new_n748), .ZN(G1339gat));
  INV_X1    g559(.A(new_n518), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n534), .A2(new_n535), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT117), .Z(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(KEYINPUT54), .A3(new_n536), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n764), .B(new_n542), .C1(KEYINPUT54), .C2(new_n536), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n544), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n766), .B2(new_n765), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n606), .A2(new_n607), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n599), .B2(new_n598), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n593), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n613), .A2(new_n768), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n761), .B1(new_n668), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n614), .A2(new_n768), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n613), .A2(new_n545), .A3(new_n774), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n635), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n614), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n776), .A2(new_n779), .B1(new_n780), .B2(new_n588), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n470), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n479), .A2(new_n429), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n614), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G113gat), .ZN(G1340gat));
  NOR2_X1   g586(.A1(new_n784), .A2(new_n638), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n330), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(G120gat), .B2(new_n788), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT119), .ZN(G1341gat));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n761), .ZN(new_n792));
  OR3_X1    g591(.A1(new_n792), .A2(KEYINPUT120), .A3(new_n502), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT120), .B1(new_n792), .B2(new_n502), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n502), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(G1342gat));
  NAND2_X1  g595(.A1(new_n785), .A2(new_n668), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT121), .B1(new_n797), .B2(KEYINPUT56), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n784), .A2(new_n635), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT121), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(G134gat), .B1(new_n797), .B2(KEYINPUT56), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n798), .A2(new_n804), .A3(new_n802), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1343gat));
  OR2_X1    g607(.A1(new_n782), .A2(KEYINPUT124), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n782), .A2(KEYINPUT124), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n465), .A2(new_n477), .A3(new_n429), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n780), .A2(G141gat), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n776), .A2(new_n779), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n588), .A2(new_n780), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(KEYINPUT57), .A3(new_n423), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n781), .B2(new_n477), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n817), .A2(new_n819), .A3(KEYINPUT123), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n465), .A2(new_n470), .A3(new_n429), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT122), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n822), .B1(new_n819), .B2(KEYINPUT123), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n820), .A2(new_n823), .A3(new_n780), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n813), .B1(new_n824), .B2(new_n302), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT58), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n827), .B(new_n813), .C1(new_n824), .C2(new_n302), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1344gat));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n820), .A2(new_n823), .A3(new_n638), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n297), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n545), .A2(new_n297), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n781), .A2(new_n477), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n818), .B1(new_n477), .B2(KEYINPUT125), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n545), .B(new_n822), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n830), .A2(new_n299), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n833), .A2(new_n834), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n832), .A2(new_n841), .ZN(G1345gat));
  NAND3_X1  g641(.A1(new_n833), .A2(new_n286), .A3(new_n761), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n820), .A2(new_n823), .A3(new_n518), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n286), .ZN(G1346gat));
  AOI21_X1  g644(.A(G162gat), .B1(new_n833), .B2(new_n668), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n820), .A2(new_n823), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n635), .A2(new_n287), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(G1347gat));
  NOR2_X1   g648(.A1(new_n781), .A2(new_n620), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n479), .A2(new_n485), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n614), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n545), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(G176gat), .ZN(G1349gat));
  OAI21_X1  g656(.A(new_n222), .B1(new_n852), .B2(new_n518), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n853), .A2(new_n761), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n244), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n860), .B(new_n861), .ZN(G1350gat));
  NOR2_X1   g661(.A1(new_n852), .A2(new_n635), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n239), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT61), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n243), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(KEYINPUT61), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G1351gat));
  NAND3_X1  g667(.A1(new_n629), .A2(new_n423), .A3(new_n429), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT126), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n869), .A2(KEYINPUT126), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n850), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(G197gat), .B1(new_n872), .B2(new_n614), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n837), .A2(new_n838), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n465), .A2(new_n485), .A3(new_n620), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n614), .A2(G197gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n873), .B1(new_n877), .B2(new_n878), .ZN(G1352gat));
  XOR2_X1   g678(.A(KEYINPUT127), .B(G204gat), .Z(new_n880));
  NAND3_X1  g679(.A1(new_n872), .A2(new_n545), .A3(new_n880), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT62), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(KEYINPUT62), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n874), .A2(new_n638), .A3(new_n876), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n880), .ZN(G1353gat));
  NAND3_X1  g684(.A1(new_n872), .A2(new_n205), .A3(new_n761), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n761), .B(new_n875), .C1(new_n837), .C2(new_n838), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n887), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT63), .B1(new_n887), .B2(G211gat), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(G1354gat));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n206), .A3(new_n668), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n874), .A2(new_n635), .A3(new_n876), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n206), .ZN(G1355gat));
endmodule


