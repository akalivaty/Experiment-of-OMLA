

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XOR2_X1 U324 ( .A(G99GAT), .B(G85GAT), .Z(n399) );
  INV_X1 U325 ( .A(KEYINPUT33), .ZN(n408) );
  XNOR2_X1 U326 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U327 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U328 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U329 ( .A(n364), .B(n363), .ZN(n370) );
  NOR2_X1 U330 ( .A1(n538), .A2(n454), .ZN(n573) );
  XNOR2_X1 U331 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U332 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G120GAT), .B(G71GAT), .Z(n393) );
  XOR2_X1 U335 ( .A(G15GAT), .B(G127GAT), .Z(n377) );
  XNOR2_X1 U336 ( .A(n393), .B(n377), .ZN(n294) );
  XOR2_X1 U337 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n293) );
  XNOR2_X1 U338 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n292) );
  XNOR2_X1 U339 ( .A(n293), .B(n292), .ZN(n449) );
  XNOR2_X1 U340 ( .A(n294), .B(n449), .ZN(n300) );
  XOR2_X1 U341 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n296) );
  XNOR2_X1 U342 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n325) );
  XOR2_X1 U344 ( .A(n325), .B(G176GAT), .Z(n298) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U347 ( .A(n300), .B(n299), .Z(n308) );
  XOR2_X1 U348 ( .A(G99GAT), .B(G190GAT), .Z(n302) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G134GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U351 ( .A(G183GAT), .B(KEYINPUT85), .Z(n304) );
  XNOR2_X1 U352 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n538) );
  XOR2_X1 U356 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n310) );
  NAND2_X1 U357 ( .A1(G228GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U359 ( .A(n311), .B(KEYINPUT22), .Z(n313) );
  XOR2_X1 U360 ( .A(G141GAT), .B(G22GAT), .Z(n335) );
  XOR2_X1 U361 ( .A(G50GAT), .B(G162GAT), .Z(n368) );
  XNOR2_X1 U362 ( .A(n335), .B(n368), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n315) );
  XNOR2_X1 U364 ( .A(G106GAT), .B(G78GAT), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n314), .B(G148GAT), .ZN(n407) );
  XOR2_X1 U366 ( .A(n315), .B(n407), .Z(n323) );
  XOR2_X1 U367 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n317) );
  XNOR2_X1 U368 ( .A(G218GAT), .B(KEYINPUT88), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U370 ( .A(n318), .B(G211GAT), .Z(n320) );
  XNOR2_X1 U371 ( .A(G197GAT), .B(G204GAT), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n329) );
  XNOR2_X1 U373 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n321) );
  XOR2_X1 U374 ( .A(n321), .B(KEYINPUT3), .Z(n450) );
  XOR2_X1 U375 ( .A(n329), .B(n450), .Z(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n479) );
  XOR2_X1 U377 ( .A(G176GAT), .B(G92GAT), .Z(n324) );
  XOR2_X1 U378 ( .A(G64GAT), .B(n324), .Z(n392) );
  XOR2_X1 U379 ( .A(KEYINPUT92), .B(n325), .Z(n327) );
  NAND2_X1 U380 ( .A1(G226GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U382 ( .A(G8GAT), .B(G183GAT), .Z(n376) );
  XOR2_X1 U383 ( .A(n328), .B(n376), .Z(n331) );
  XOR2_X1 U384 ( .A(G36GAT), .B(G190GAT), .Z(n357) );
  XNOR2_X1 U385 ( .A(n329), .B(n357), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U387 ( .A(n392), .B(n332), .Z(n536) );
  INV_X1 U388 ( .A(KEYINPUT111), .ZN(n418) );
  XOR2_X1 U389 ( .A(G197GAT), .B(G113GAT), .Z(n334) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(G15GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n350) );
  XOR2_X1 U392 ( .A(n335), .B(G36GAT), .Z(n339) );
  XOR2_X1 U393 ( .A(G29GAT), .B(G43GAT), .Z(n337) );
  XNOR2_X1 U394 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n360) );
  XNOR2_X1 U396 ( .A(n360), .B(G50GAT), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U398 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n341) );
  NAND2_X1 U399 ( .A1(G229GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U401 ( .A(n343), .B(n342), .Z(n348) );
  XOR2_X1 U402 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n345) );
  XNOR2_X1 U403 ( .A(G1GAT), .B(G8GAT), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n346), .B(KEYINPUT29), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U407 ( .A(n350), .B(n349), .Z(n517) );
  XOR2_X1 U408 ( .A(KEYINPUT80), .B(KEYINPUT10), .Z(n352) );
  XNOR2_X1 U409 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n353), .B(KEYINPUT75), .ZN(n355) );
  XOR2_X1 U412 ( .A(G218GAT), .B(n399), .Z(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n356), .B(KEYINPUT76), .ZN(n364) );
  XOR2_X1 U415 ( .A(G134GAT), .B(KEYINPUT79), .Z(n441) );
  XOR2_X1 U416 ( .A(n357), .B(n441), .Z(n359) );
  NAND2_X1 U417 ( .A1(G232GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n360), .B(KEYINPUT78), .ZN(n361) );
  XOR2_X1 U420 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n366) );
  XNOR2_X1 U421 ( .A(G92GAT), .B(KEYINPUT77), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n562) );
  INV_X1 U425 ( .A(KEYINPUT36), .ZN(n371) );
  XNOR2_X1 U426 ( .A(n562), .B(n371), .ZN(n588) );
  XOR2_X1 U427 ( .A(KEYINPUT15), .B(G64GAT), .Z(n373) );
  XNOR2_X1 U428 ( .A(G1GAT), .B(G78GAT), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n375) );
  XNOR2_X1 U430 ( .A(G57GAT), .B(KEYINPUT68), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n374), .B(KEYINPUT13), .ZN(n391) );
  XOR2_X1 U432 ( .A(n375), .B(n391), .Z(n379) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U435 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n381) );
  NAND2_X1 U436 ( .A1(G231GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U438 ( .A(n383), .B(n382), .Z(n388) );
  XOR2_X1 U439 ( .A(G155GAT), .B(G211GAT), .Z(n385) );
  XNOR2_X1 U440 ( .A(G22GAT), .B(G71GAT), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n386), .B(KEYINPUT81), .ZN(n387) );
  XOR2_X1 U443 ( .A(n388), .B(n387), .Z(n585) );
  INV_X1 U444 ( .A(n585), .ZN(n502) );
  NOR2_X1 U445 ( .A1(n588), .A2(n502), .ZN(n390) );
  INV_X1 U446 ( .A(KEYINPUT45), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n414) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n413) );
  XNOR2_X1 U449 ( .A(n393), .B(G204GAT), .ZN(n397) );
  XOR2_X1 U450 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n395) );
  XNOR2_X1 U451 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n404) );
  INV_X1 U454 ( .A(n399), .ZN(n398) );
  NAND2_X1 U455 ( .A1(KEYINPUT32), .A2(n398), .ZN(n402) );
  INV_X1 U456 ( .A(KEYINPUT32), .ZN(n400) );
  NAND2_X1 U457 ( .A1(n400), .A2(n399), .ZN(n401) );
  NAND2_X1 U458 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n406) );
  AND2_X1 U460 ( .A1(G230GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n411) );
  XNOR2_X1 U462 ( .A(n407), .B(KEYINPUT31), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n413), .B(n412), .ZN(n582) );
  NOR2_X1 U464 ( .A1(n414), .A2(n582), .ZN(n415) );
  XNOR2_X1 U465 ( .A(n415), .B(KEYINPUT110), .ZN(n416) );
  AND2_X1 U466 ( .A1(n517), .A2(n416), .ZN(n417) );
  XOR2_X1 U467 ( .A(n418), .B(n417), .Z(n425) );
  XOR2_X1 U468 ( .A(KEYINPUT41), .B(n582), .Z(n570) );
  INV_X1 U469 ( .A(n570), .ZN(n518) );
  NOR2_X1 U470 ( .A1(n518), .A2(n517), .ZN(n420) );
  XNOR2_X1 U471 ( .A(KEYINPUT109), .B(KEYINPUT46), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n421) );
  NAND2_X1 U473 ( .A1(n421), .A2(n502), .ZN(n422) );
  NOR2_X1 U474 ( .A1(n562), .A2(n422), .ZN(n423) );
  XNOR2_X1 U475 ( .A(KEYINPUT47), .B(n423), .ZN(n424) );
  AND2_X1 U476 ( .A1(n425), .A2(n424), .ZN(n428) );
  XNOR2_X1 U477 ( .A(KEYINPUT64), .B(KEYINPUT112), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n426), .B(KEYINPUT48), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n428), .B(n427), .ZN(n460) );
  NOR2_X1 U480 ( .A1(n536), .A2(n460), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n429), .B(KEYINPUT54), .ZN(n452) );
  XOR2_X1 U482 ( .A(G148GAT), .B(G127GAT), .Z(n431) );
  XNOR2_X1 U483 ( .A(G1GAT), .B(G141GAT), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U485 ( .A(G57GAT), .B(KEYINPUT89), .Z(n433) );
  XNOR2_X1 U486 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U488 ( .A(n435), .B(n434), .Z(n447) );
  XOR2_X1 U489 ( .A(KEYINPUT91), .B(KEYINPUT4), .Z(n437) );
  XNOR2_X1 U490 ( .A(KEYINPUT90), .B(KEYINPUT5), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n445) );
  XOR2_X1 U492 ( .A(G85GAT), .B(G162GAT), .Z(n439) );
  XNOR2_X1 U493 ( .A(G29GAT), .B(G120GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U495 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U496 ( .A1(G225GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n451) );
  XOR2_X1 U501 ( .A(n451), .B(n450), .Z(n459) );
  INV_X1 U502 ( .A(n459), .ZN(n532) );
  NAND2_X1 U503 ( .A1(n452), .A2(n532), .ZN(n576) );
  NOR2_X1 U504 ( .A1(n479), .A2(n576), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n453), .B(KEYINPUT55), .ZN(n454) );
  NAND2_X1 U506 ( .A1(n573), .A2(n562), .ZN(n458) );
  XOR2_X1 U507 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n456) );
  XNOR2_X1 U508 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n455) );
  XOR2_X1 U509 ( .A(n479), .B(KEYINPUT28), .Z(n541) );
  INV_X1 U510 ( .A(n541), .ZN(n473) );
  XOR2_X1 U511 ( .A(n536), .B(KEYINPUT27), .Z(n481) );
  NAND2_X1 U512 ( .A1(n459), .A2(n481), .ZN(n472) );
  NOR2_X1 U513 ( .A1(n472), .A2(n460), .ZN(n461) );
  XNOR2_X1 U514 ( .A(n461), .B(KEYINPUT113), .ZN(n553) );
  NOR2_X1 U515 ( .A1(n553), .A2(n538), .ZN(n463) );
  INV_X1 U516 ( .A(KEYINPUT114), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n463), .B(n462), .ZN(n464) );
  NOR2_X2 U518 ( .A1(n473), .A2(n464), .ZN(n548) );
  NAND2_X1 U519 ( .A1(n548), .A2(n562), .ZN(n468) );
  XOR2_X1 U520 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n466) );
  INV_X1 U521 ( .A(G134GAT), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n468), .B(n467), .ZN(G1343GAT) );
  XOR2_X1 U523 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n470) );
  XNOR2_X1 U524 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n470), .B(n469), .ZN(n492) );
  NOR2_X1 U526 ( .A1(n517), .A2(n582), .ZN(n471) );
  XOR2_X1 U527 ( .A(KEYINPUT73), .B(n471), .Z(n504) );
  NOR2_X1 U528 ( .A1(n473), .A2(n472), .ZN(n474) );
  NAND2_X1 U529 ( .A1(n538), .A2(n474), .ZN(n475) );
  XOR2_X1 U530 ( .A(KEYINPUT93), .B(n475), .Z(n486) );
  XNOR2_X1 U531 ( .A(KEYINPUT94), .B(KEYINPUT25), .ZN(n478) );
  NOR2_X1 U532 ( .A1(n538), .A2(n536), .ZN(n476) );
  NOR2_X1 U533 ( .A1(n479), .A2(n476), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n478), .B(n477), .ZN(n483) );
  NAND2_X1 U535 ( .A1(n479), .A2(n538), .ZN(n480) );
  XOR2_X1 U536 ( .A(n480), .B(KEYINPUT26), .Z(n552) );
  NAND2_X1 U537 ( .A1(n481), .A2(n552), .ZN(n482) );
  NAND2_X1 U538 ( .A1(n483), .A2(n482), .ZN(n484) );
  NAND2_X1 U539 ( .A1(n532), .A2(n484), .ZN(n485) );
  NAND2_X1 U540 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U541 ( .A(KEYINPUT95), .B(n487), .ZN(n500) );
  NOR2_X1 U542 ( .A1(n562), .A2(n502), .ZN(n488) );
  XOR2_X1 U543 ( .A(KEYINPUT16), .B(n488), .Z(n489) );
  XNOR2_X1 U544 ( .A(n489), .B(KEYINPUT82), .ZN(n490) );
  NOR2_X1 U545 ( .A1(n500), .A2(n490), .ZN(n519) );
  NAND2_X1 U546 ( .A1(n504), .A2(n519), .ZN(n496) );
  NOR2_X1 U547 ( .A1(n532), .A2(n496), .ZN(n491) );
  XOR2_X1 U548 ( .A(n492), .B(n491), .Z(G1324GAT) );
  NOR2_X1 U549 ( .A1(n536), .A2(n496), .ZN(n493) );
  XOR2_X1 U550 ( .A(G8GAT), .B(n493), .Z(G1325GAT) );
  NOR2_X1 U551 ( .A1(n538), .A2(n496), .ZN(n495) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NOR2_X1 U554 ( .A1(n541), .A2(n496), .ZN(n498) );
  XNOR2_X1 U555 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(n499), .ZN(G1327GAT) );
  NOR2_X1 U558 ( .A1(n588), .A2(n500), .ZN(n501) );
  NAND2_X1 U559 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U560 ( .A(KEYINPUT37), .B(n503), .ZN(n531) );
  NAND2_X1 U561 ( .A1(n504), .A2(n531), .ZN(n505) );
  XNOR2_X1 U562 ( .A(n505), .B(KEYINPUT38), .ZN(n515) );
  NOR2_X1 U563 ( .A1(n515), .A2(n532), .ZN(n508) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n506) );
  XNOR2_X1 U565 ( .A(n506), .B(KEYINPUT100), .ZN(n507) );
  XNOR2_X1 U566 ( .A(n508), .B(n507), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n536), .A2(n515), .ZN(n509) );
  XOR2_X1 U568 ( .A(G36GAT), .B(n509), .Z(G1329GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n511) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U572 ( .A(KEYINPUT101), .B(n512), .ZN(n514) );
  NOR2_X1 U573 ( .A1(n538), .A2(n515), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n514), .B(n513), .ZN(G1330GAT) );
  NOR2_X1 U575 ( .A1(n541), .A2(n515), .ZN(n516) );
  XOR2_X1 U576 ( .A(G50GAT), .B(n516), .Z(G1331GAT) );
  INV_X1 U577 ( .A(n517), .ZN(n578) );
  NOR2_X1 U578 ( .A1(n578), .A2(n518), .ZN(n530) );
  NAND2_X1 U579 ( .A1(n530), .A2(n519), .ZN(n524) );
  NOR2_X1 U580 ( .A1(n532), .A2(n524), .ZN(n520) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n520), .Z(n521) );
  XNOR2_X1 U582 ( .A(KEYINPUT42), .B(n521), .ZN(G1332GAT) );
  NOR2_X1 U583 ( .A1(n536), .A2(n524), .ZN(n522) );
  XOR2_X1 U584 ( .A(G64GAT), .B(n522), .Z(G1333GAT) );
  NOR2_X1 U585 ( .A1(n538), .A2(n524), .ZN(n523) );
  XOR2_X1 U586 ( .A(G71GAT), .B(n523), .Z(G1334GAT) );
  NOR2_X1 U587 ( .A1(n541), .A2(n524), .ZN(n529) );
  XOR2_X1 U588 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n526) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(KEYINPUT104), .B(n527), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(G1335GAT) );
  NAND2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n540) );
  NOR2_X1 U594 ( .A1(n532), .A2(n540), .ZN(n534) );
  XNOR2_X1 U595 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U597 ( .A(G85GAT), .B(n535), .ZN(G1336GAT) );
  NOR2_X1 U598 ( .A1(n536), .A2(n540), .ZN(n537) );
  XOR2_X1 U599 ( .A(G92GAT), .B(n537), .Z(G1337GAT) );
  NOR2_X1 U600 ( .A1(n538), .A2(n540), .ZN(n539) );
  XOR2_X1 U601 ( .A(G99GAT), .B(n539), .Z(G1338GAT) );
  NOR2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U603 ( .A(KEYINPUT44), .B(n542), .Z(n543) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(n543), .ZN(G1339GAT) );
  NAND2_X1 U605 ( .A1(n578), .A2(n548), .ZN(n544) );
  XNOR2_X1 U606 ( .A(n544), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n546) );
  NAND2_X1 U608 ( .A1(n548), .A2(n570), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U610 ( .A(G120GAT), .B(n547), .Z(G1341GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n550) );
  NAND2_X1 U612 ( .A1(n548), .A2(n585), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U614 ( .A(G127GAT), .B(n551), .Z(G1342GAT) );
  INV_X1 U615 ( .A(n552), .ZN(n577) );
  NOR2_X1 U616 ( .A1(n577), .A2(n553), .ZN(n563) );
  NAND2_X1 U617 ( .A1(n563), .A2(n578), .ZN(n554) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U621 ( .A1(n563), .A2(n570), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n560) );
  NAND2_X1 U625 ( .A1(n563), .A2(n585), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U630 ( .A(G169GAT), .B(KEYINPUT121), .Z(n566) );
  NAND2_X1 U631 ( .A1(n573), .A2(n578), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n568) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT56), .B(n569), .Z(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1349GAT) );
  NAND2_X1 U639 ( .A1(n585), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT124), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G183GAT), .B(n575), .ZN(G1350GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n587) );
  NAND2_X1 U644 ( .A1(n587), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U648 ( .A1(n587), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n587), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U652 ( .A(KEYINPUT62), .ZN(n591) );
  INV_X1 U653 ( .A(n587), .ZN(n589) );
  NOR2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

