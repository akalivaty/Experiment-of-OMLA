//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(G137), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G131), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n198), .A2(new_n193), .A3(new_n192), .A4(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n203));
  OAI21_X1  g017(.A(G128), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n205), .B1(G143), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT64), .A2(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT64), .A2(G143), .ZN(new_n210));
  AOI21_X1  g024(.A(G146), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(G143), .ZN(new_n212));
  OAI22_X1  g026(.A1(new_n204), .A2(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(G146), .A3(new_n210), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n201), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n214), .A2(new_n205), .A3(G128), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT79), .ZN(new_n219));
  INV_X1    g033(.A(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n219), .A2(new_n224), .A3(new_n220), .A4(G104), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n220), .A2(G104), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n222), .A2(new_n223), .A3(new_n225), .A4(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G107), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n230), .B2(new_n226), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n218), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(G128), .B1(new_n211), .B2(new_n205), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n214), .A2(new_n216), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n232), .B1(new_n237), .B2(new_n217), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n200), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT12), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(new_n207), .B2(KEYINPUT66), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n202), .A2(new_n203), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT64), .A2(G143), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT64), .A2(G143), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n206), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n212), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n243), .A2(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n217), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n241), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n213), .A2(KEYINPUT69), .A3(new_n217), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT10), .A4(new_n233), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n242), .B1(new_n247), .B2(KEYINPUT1), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n245), .A2(new_n246), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n215), .B1(new_n255), .B2(G146), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n217), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n233), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT10), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n226), .B1(new_n221), .B2(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n225), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G101), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT4), .A3(new_n228), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n236), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT0), .B(G128), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(new_n247), .B2(new_n248), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n262), .A2(new_n270), .A3(G101), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n264), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n200), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n253), .A2(new_n260), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  INV_X1    g089(.A(G953), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n276), .A2(G227), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n275), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT12), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n280), .B(new_n200), .C1(new_n234), .C2(new_n238), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n240), .A2(new_n274), .A3(new_n279), .A4(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n253), .A2(new_n260), .A3(new_n272), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n200), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n279), .B1(new_n284), .B2(new_n274), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n282), .B1(new_n285), .B2(KEYINPUT80), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n282), .A2(KEYINPUT80), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G469), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT74), .B(G902), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n240), .A2(new_n274), .A3(new_n281), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n278), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n284), .A2(new_n279), .A3(new_n274), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G469), .B1(new_n295), .B2(G902), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n189), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G214), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G116), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n302));
  INV_X1    g116(.A(G116), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n303), .B2(G119), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n300), .A2(KEYINPUT67), .A3(G116), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT2), .B(G113), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT67), .B1(new_n300), .B2(G116), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n302), .A2(new_n303), .A3(G119), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n313), .A2(new_n314), .B1(G116), .B2(new_n300), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT68), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n310), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G113), .B1(new_n301), .B2(KEYINPUT5), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n309), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n232), .A2(new_n308), .ZN(new_n320));
  INV_X1    g134(.A(new_n318), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n306), .B2(new_n310), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n319), .A2(new_n232), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(G110), .B(G122), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT81), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n325), .B(KEYINPUT8), .Z(new_n326));
  OAI21_X1  g140(.A(KEYINPUT82), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT82), .ZN(new_n328));
  INV_X1    g142(.A(new_n326), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n306), .A2(new_n311), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n315), .A2(KEYINPUT68), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT5), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n321), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n233), .B1(new_n333), .B2(new_n309), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n320), .A2(new_n322), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n328), .B(new_n329), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n327), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n320), .B1(new_n317), .B2(new_n318), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n312), .A2(new_n316), .ZN(new_n339));
  INV_X1    g153(.A(new_n307), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n309), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n264), .A2(new_n271), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n325), .B(new_n338), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G125), .B1(new_n266), .B2(new_n268), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n218), .B2(G125), .ZN(new_n346));
  INV_X1    g160(.A(G224), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT7), .B1(new_n347), .B2(G953), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n346), .A2(new_n348), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n344), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(G902), .B1(new_n337), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n338), .B1(new_n342), .B2(new_n343), .ZN(new_n353));
  INV_X1    g167(.A(new_n325), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT6), .A3(new_n344), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n357), .A3(new_n354), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n347), .A2(G953), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n346), .B(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n352), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G210), .B1(G237), .B2(G902), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n352), .A2(new_n363), .A3(new_n361), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n299), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(G234), .A2(G237), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(G952), .A3(new_n276), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n369), .B(KEYINPUT92), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n290), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n372), .A2(G953), .A3(new_n368), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT21), .B(G898), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n375), .B(KEYINPUT93), .Z(new_n376));
  NAND3_X1  g190(.A1(new_n297), .A2(new_n367), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT17), .ZN(new_n379));
  INV_X1    g193(.A(new_n198), .ZN(new_n380));
  INV_X1    g194(.A(G237), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n276), .A3(G214), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT83), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n209), .A3(new_n383), .A4(new_n210), .ZN(new_n384));
  INV_X1    g198(.A(G214), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n385), .A2(G237), .A3(G953), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G143), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n383), .B1(new_n255), .B2(new_n382), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n380), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(KEYINPUT84), .B(new_n380), .C1(new_n388), .C2(new_n389), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n379), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G125), .ZN(new_n396));
  INV_X1    g210(.A(G125), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G140), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n398), .A3(KEYINPUT16), .ZN(new_n399));
  OR3_X1    g213(.A1(new_n397), .A2(KEYINPUT16), .A3(G140), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(new_n206), .ZN(new_n402));
  AOI21_X1  g216(.A(G146), .B1(new_n399), .B2(new_n400), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n378), .B1(new_n394), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n393), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT64), .B(G143), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT83), .B1(new_n408), .B2(new_n386), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n387), .A3(new_n384), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT84), .B1(new_n410), .B2(new_n380), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT17), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT87), .A3(new_n404), .ZN(new_n413));
  INV_X1    g227(.A(new_n410), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n198), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n415), .A2(new_n392), .A3(new_n379), .A4(new_n393), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n406), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(KEYINPUT18), .A2(G131), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n410), .A2(KEYINPUT18), .A3(G131), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n396), .A2(new_n398), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(new_n206), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G113), .B(G122), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT86), .B(G104), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n424), .B(new_n425), .Z(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT85), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT19), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n206), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n415), .A2(new_n392), .A3(new_n393), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT77), .B1(new_n401), .B2(new_n206), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT77), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n399), .A2(new_n400), .A3(new_n435), .A4(G146), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n432), .A2(new_n433), .A3(new_n434), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n423), .ZN(new_n438));
  INV_X1    g252(.A(new_n426), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n427), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(G475), .A2(G902), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT20), .ZN(new_n445));
  INV_X1    g259(.A(new_n442), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n427), .B2(new_n440), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT88), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n445), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n427), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n426), .B1(new_n417), .B2(new_n423), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G475), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n303), .A2(KEYINPUT14), .A3(G122), .ZN(new_n457));
  XOR2_X1   g271(.A(G116), .B(G122), .Z(new_n458));
  OAI211_X1 g272(.A(G107), .B(new_n457), .C1(new_n458), .C2(KEYINPUT14), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT91), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n458), .A2(G107), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT90), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n255), .A2(G128), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n242), .A2(G143), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(G134), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n460), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n466), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n458), .A2(G107), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n469), .A2(new_n191), .B1(new_n461), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n255), .A2(KEYINPUT13), .A3(G128), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT89), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n465), .A2(KEYINPUT13), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n474), .B1(new_n464), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G134), .B1(new_n472), .B2(new_n473), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G217), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n187), .A2(new_n479), .A3(G953), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n468), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n480), .B1(new_n468), .B2(new_n478), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n290), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G478), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI221_X1 g301(.A(new_n290), .B1(KEYINPUT15), .B2(new_n485), .C1(new_n482), .C2(new_n483), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n451), .A2(new_n456), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n377), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n479), .B1(new_n290), .B2(G234), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n300), .A2(G128), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n242), .A2(KEYINPUT23), .A3(G119), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n300), .A2(G128), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(KEYINPUT23), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G110), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n242), .A2(G119), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT24), .B(G110), .ZN(new_n502));
  OAI221_X1 g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .C1(new_n402), .C2(new_n403), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n276), .A2(G221), .A3(G234), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT78), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT22), .B(G137), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(KEYINPUT75), .A2(G110), .ZN(new_n508));
  NOR2_X1   g322(.A1(KEYINPUT75), .A2(G110), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT23), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n500), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n510), .A2(new_n512), .A3(new_n495), .A4(new_n496), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n501), .A2(new_n502), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(KEYINPUT76), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT76), .B1(new_n513), .B2(new_n514), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n421), .A2(new_n206), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n434), .A2(new_n436), .A3(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n503), .B(new_n507), .C1(new_n518), .C2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n434), .A2(new_n436), .A3(new_n519), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n508), .A2(new_n509), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n514), .B1(new_n498), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT76), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n515), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n507), .B1(new_n529), .B2(new_n503), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n290), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT25), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n503), .B1(new_n518), .B2(new_n520), .ZN(new_n534));
  INV_X1    g348(.A(new_n507), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n521), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT25), .A3(new_n290), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n494), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n494), .A2(new_n452), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n536), .B2(new_n521), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n194), .A2(G134), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n193), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G131), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n199), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n251), .A2(new_n548), .A3(new_n252), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n269), .A2(new_n200), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(KEYINPUT30), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n273), .A2(new_n268), .A3(new_n266), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n547), .B1(new_n213), .B2(new_n217), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n551), .A2(new_n555), .A3(new_n341), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n342), .A2(new_n549), .A3(new_n550), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n381), .A2(new_n276), .A3(G210), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT27), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT26), .B(G101), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT31), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n556), .A2(new_n557), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT28), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n341), .B1(new_n553), .B2(new_n554), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n566), .B1(new_n557), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n549), .A2(new_n550), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT71), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT71), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n549), .A2(new_n571), .A3(new_n550), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n342), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n568), .B1(new_n573), .B2(new_n566), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n563), .B(new_n565), .C1(new_n574), .C2(new_n561), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n575), .B2(new_n576), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n341), .B1(new_n569), .B2(KEYINPUT71), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT28), .B1(new_n581), .B2(new_n572), .ZN(new_n582));
  INV_X1    g396(.A(new_n561), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n582), .A2(new_n568), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n556), .A2(new_n557), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n583), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT29), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT73), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n573), .A2(new_n566), .ZN(new_n590));
  INV_X1    g404(.A(new_n557), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n342), .B1(new_n549), .B2(new_n550), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT28), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n583), .A2(new_n587), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n595), .A2(new_n290), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n574), .A2(new_n561), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT73), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT29), .B1(new_n585), .B2(new_n583), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n589), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G472), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n543), .B1(new_n580), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n492), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  NAND2_X1  g419(.A1(new_n575), .A2(new_n576), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n575), .A2(new_n290), .ZN(new_n607));
  OAI21_X1  g421(.A(G472), .B1(new_n607), .B2(KEYINPUT94), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n575), .B2(new_n290), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n606), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n297), .A2(new_n542), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n482), .A2(new_n483), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n372), .A2(new_n485), .ZN(new_n617));
  NAND2_X1  g431(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n616), .B(new_n617), .C1(new_n614), .C2(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n485), .A2(KEYINPUT96), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n485), .A2(KEYINPUT96), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n484), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n451), .B2(new_n456), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n352), .A2(new_n363), .A3(new_n361), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n363), .B1(new_n352), .B2(new_n361), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n298), .B(new_n376), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n613), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  AOI21_X1  g447(.A(new_n444), .B1(new_n443), .B2(KEYINPUT20), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n447), .A2(KEYINPUT88), .A3(new_n448), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT97), .B1(new_n445), .B2(new_n449), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n450), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n456), .A2(new_n489), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n630), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n636), .B1(new_n634), .B2(new_n635), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n445), .A2(KEYINPUT97), .A3(new_n449), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n640), .B1(new_n647), .B2(new_n450), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(KEYINPUT98), .A3(new_n630), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n613), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n507), .A2(KEYINPUT36), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n534), .B(new_n654), .Z(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n540), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT99), .B1(new_n539), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT25), .B1(new_n537), .B2(new_n290), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n532), .B(new_n372), .C1(new_n536), .C2(new_n521), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n493), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n655), .A2(new_n540), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT99), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n606), .B(new_n664), .C1(new_n608), .C2(new_n610), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n492), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  NAND2_X1  g483(.A1(new_n580), .A2(new_n602), .ZN(new_n670));
  AND4_X1   g484(.A1(new_n670), .A2(new_n367), .A3(new_n297), .A4(new_n664), .ZN(new_n671));
  INV_X1    g485(.A(new_n450), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n645), .B2(new_n646), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n373), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n675), .A2(new_n370), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n673), .A2(new_n640), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  NOR2_X1   g493(.A1(new_n627), .A2(new_n628), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(G472), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n583), .B1(new_n591), .B2(new_n592), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n562), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n685), .B1(new_n687), .B2(new_n452), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n577), .A2(new_n579), .A3(new_n688), .ZN(new_n689));
  NOR4_X1   g503(.A1(new_n684), .A2(new_n689), .A3(new_n299), .A4(new_n664), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n291), .A2(new_n296), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n188), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n676), .B(KEYINPUT39), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n490), .B1(new_n451), .B2(new_n456), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n690), .A2(new_n695), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n408), .ZN(G45));
  AOI211_X1 g513(.A(new_n676), .B(new_n625), .C1(new_n451), .C2(new_n456), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n671), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  AND2_X1   g516(.A1(new_n286), .A2(new_n287), .ZN(new_n703));
  OAI21_X1  g517(.A(G469), .B1(new_n703), .B2(new_n372), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n188), .A3(new_n291), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n603), .A2(new_n626), .A3(new_n630), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND2_X1  g523(.A1(new_n603), .A2(new_n706), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT98), .B1(new_n648), .B2(new_n630), .ZN(new_n712));
  NOR4_X1   g526(.A1(new_n673), .A2(new_n643), .A3(new_n629), .A4(new_n640), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  NOR2_X1   g529(.A1(new_n705), .A2(new_n629), .ZN(new_n716));
  INV_X1    g530(.A(new_n491), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n670), .A4(new_n664), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  OR3_X1    g533(.A1(new_n539), .A2(KEYINPUT102), .A3(new_n541), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT102), .B1(new_n539), .B2(new_n541), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n563), .A2(new_n565), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n561), .B1(new_n590), .B2(new_n593), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n576), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT101), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n607), .A2(G472), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT101), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n728), .B(new_n576), .C1(new_n723), .C2(new_n724), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n722), .A2(new_n726), .A3(new_n727), .A4(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n716), .A2(new_n730), .A3(new_n696), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND4_X1  g546(.A1(new_n727), .A2(new_n726), .A3(new_n664), .A4(new_n729), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n705), .A2(new_n299), .A3(new_n680), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n700), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  NAND2_X1  g552(.A1(new_n595), .A2(new_n290), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n597), .A2(new_n599), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n739), .B1(new_n740), .B2(KEYINPUT73), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n685), .B1(new_n741), .B2(new_n600), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT32), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n606), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n576), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n722), .B1(new_n742), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n365), .A2(new_n298), .A3(new_n366), .A4(new_n188), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  AOI211_X1 g564(.A(G469), .B(new_n372), .C1(new_n286), .C2(new_n287), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n294), .A2(KEYINPUT104), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n284), .A2(new_n753), .A3(new_n279), .A4(new_n274), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n752), .A2(G469), .A3(new_n293), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(G469), .A2(G902), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n750), .B1(new_n751), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n755), .A2(new_n756), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n291), .A3(KEYINPUT105), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n749), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n748), .A2(KEYINPUT42), .A3(new_n700), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n761), .A2(new_n670), .A3(new_n542), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n763), .B1(new_n764), .B2(new_n700), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n700), .A2(new_n603), .A3(new_n763), .A4(new_n761), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n762), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  NAND2_X1  g584(.A1(new_n764), .A2(new_n677), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  AND2_X1   g586(.A1(new_n451), .A2(new_n456), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n624), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT43), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n611), .A2(new_n664), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n451), .A2(new_n456), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n777), .A2(KEYINPUT43), .A3(new_n625), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(KEYINPUT44), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n680), .A2(new_n298), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n752), .A2(KEYINPUT45), .A3(new_n293), .A4(new_n754), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT107), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(KEYINPUT107), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n295), .A2(KEYINPUT45), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n784), .A2(G469), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT46), .B1(new_n787), .B2(new_n756), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n751), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n756), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n189), .A3(new_n693), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n775), .A2(new_n778), .A3(new_n776), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n782), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(KEYINPUT108), .B(G137), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(G39));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n189), .B1(new_n789), .B2(new_n790), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n676), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n626), .A2(new_n803), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n804), .A2(new_n670), .A3(new_n542), .A4(new_n780), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT109), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n799), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n801), .B1(new_n791), .B2(new_n189), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n800), .A2(KEYINPUT47), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n805), .B(KEYINPUT109), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(KEYINPUT110), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G140), .ZN(G42));
  NAND2_X1  g629(.A1(new_n704), .A2(new_n291), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT111), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT49), .ZN(new_n818));
  INV_X1    g632(.A(new_n774), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n298), .A2(new_n684), .A3(new_n188), .A4(new_n722), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n818), .A2(new_n689), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n671), .B1(new_n677), .B2(new_n700), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n660), .A2(new_n661), .A3(new_n188), .A4(new_n803), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n689), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n758), .A2(new_n760), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n367), .A3(new_n696), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n822), .A2(new_n737), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n822), .A2(new_n737), .A3(KEYINPUT52), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND4_X1   g645(.A1(KEYINPUT42), .A2(new_n748), .A3(new_n700), .A4(new_n761), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n766), .A2(new_n767), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n603), .A2(new_n761), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT106), .B1(new_n834), .B2(new_n804), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n832), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n707), .A2(new_n718), .A3(new_n731), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n714), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n487), .A2(new_n488), .A3(new_n803), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n455), .B2(G475), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n680), .A2(new_n664), .A3(new_n841), .A4(new_n298), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n692), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n639), .A3(new_n670), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n639), .A3(KEYINPUT112), .A4(new_n670), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n846), .A2(new_n847), .B1(new_n677), .B2(new_n764), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n777), .A2(new_n624), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n777), .B2(new_n490), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n630), .A3(new_n613), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n492), .B1(new_n666), .B2(new_n603), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n735), .A2(new_n700), .A3(new_n761), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n848), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n831), .A2(new_n839), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n707), .A2(new_n718), .A3(new_n731), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n650), .B2(new_n711), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n769), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n855), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(KEYINPUT53), .A3(new_n831), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n859), .A2(KEYINPUT113), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n857), .A2(new_n866), .A3(new_n858), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(KEYINPUT54), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n705), .A2(new_n780), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n689), .A3(new_n542), .A4(new_n371), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n777), .A3(new_n624), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n371), .A2(new_n775), .A3(new_n778), .A4(new_n869), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n871), .B1(new_n872), .B2(new_n735), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n298), .B1(new_n682), .B2(new_n683), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n706), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT115), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n877), .A3(new_n706), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n775), .A2(new_n371), .A3(new_n730), .A4(new_n778), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT50), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n876), .A2(new_n878), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT50), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(new_n884), .A3(new_n880), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n873), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n879), .A2(KEYINPUT50), .A3(new_n881), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n884), .B1(new_n883), .B2(new_n880), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(KEYINPUT116), .A3(new_n873), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n817), .A2(new_n189), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n809), .A2(new_n810), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n880), .A2(new_n780), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n888), .A2(new_n892), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g712(.A(G952), .B(new_n276), .C1(new_n870), .C2(new_n849), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n881), .B2(new_n736), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT48), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n872), .A2(new_n901), .A3(new_n748), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n872), .B2(new_n748), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n895), .A2(new_n896), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n891), .A3(new_n873), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n904), .B1(new_n906), .B2(new_n893), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n898), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT114), .B1(new_n836), .B2(new_n838), .ZN(new_n910));
  AND4_X1   g724(.A1(KEYINPUT53), .A2(new_n848), .A3(new_n853), .A4(new_n854), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT114), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n861), .A2(new_n769), .A3(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n910), .A2(new_n831), .A3(new_n911), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n859), .A2(new_n909), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n868), .A2(new_n908), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(G952), .A2(G953), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT118), .Z(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n916), .B2(new_n917), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n821), .B1(new_n918), .B2(new_n921), .ZN(G75));
  NOR2_X1   g736(.A1(new_n276), .A2(G952), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT56), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n859), .A2(new_n914), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n372), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n925), .B1(new_n927), .B2(new_n363), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n356), .A2(new_n358), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(new_n360), .Z(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n924), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n931), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT119), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n928), .A2(KEYINPUT119), .A3(new_n931), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G51));
  NOR2_X1   g751(.A1(new_n927), .A2(new_n787), .ZN(new_n938));
  AND4_X1   g752(.A1(new_n831), .A2(new_n910), .A3(new_n911), .A4(new_n913), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT53), .B1(new_n863), .B2(new_n831), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT54), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n915), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n756), .B(KEYINPUT57), .Z(new_n943));
  AOI21_X1  g757(.A(new_n703), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n938), .B1(new_n944), .B2(KEYINPUT120), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT120), .ZN(new_n946));
  INV_X1    g760(.A(new_n943), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n941), .B2(new_n915), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n948), .B2(new_n703), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n923), .B1(new_n945), .B2(new_n949), .ZN(G54));
  AND4_X1   g764(.A1(KEYINPUT58), .A2(new_n926), .A3(G475), .A4(new_n372), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n924), .B1(new_n951), .B2(new_n441), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n441), .B2(new_n951), .ZN(G60));
  INV_X1    g767(.A(new_n942), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n616), .B1(new_n614), .B2(new_n619), .ZN(new_n955));
  NAND2_X1  g769(.A1(G478), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT59), .Z(new_n957));
  OR2_X1    g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n924), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n868), .A2(new_n915), .ZN(new_n960));
  INV_X1    g774(.A(new_n957), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n959), .B1(new_n955), .B2(new_n962), .ZN(G63));
  NAND2_X1  g777(.A1(G217), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT60), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n859), .B2(new_n914), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n924), .B1(new_n966), .B2(new_n537), .ZN(new_n967));
  AOI211_X1 g781(.A(new_n655), .B(new_n965), .C1(new_n859), .C2(new_n914), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n969));
  OAI22_X1  g783(.A1(new_n967), .A2(new_n968), .B1(KEYINPUT121), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(KEYINPUT121), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT122), .Z(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  OAI221_X1 g788(.A(new_n972), .B1(KEYINPUT121), .B2(new_n969), .C1(new_n967), .C2(new_n968), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(G66));
  OAI21_X1  g790(.A(G953), .B1(new_n374), .B2(new_n347), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT123), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n861), .A2(new_n853), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n978), .B1(new_n980), .B2(G953), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n929), .B1(G898), .B2(new_n276), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G69));
  NAND4_X1  g797(.A1(new_n792), .A2(new_n367), .A3(new_n696), .A4(new_n748), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n822), .A2(new_n737), .A3(new_n771), .ZN(new_n985));
  AND4_X1   g799(.A1(new_n769), .A2(new_n984), .A3(new_n796), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n814), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n276), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n276), .A2(G900), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n988), .A2(KEYINPUT125), .A3(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT125), .ZN(new_n992));
  AOI21_X1  g806(.A(G953), .B1(new_n986), .B2(new_n814), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(new_n989), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n551), .A2(new_n555), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(new_n431), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n276), .B1(G227), .B2(G900), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n694), .A2(new_n780), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1002), .A2(new_n603), .A3(new_n850), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n796), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT124), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n796), .A2(KEYINPUT124), .A3(new_n1003), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n698), .A2(new_n737), .A3(new_n822), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT62), .Z(new_n1010));
  NAND3_X1  g824(.A1(new_n1008), .A2(new_n814), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n998), .B1(new_n1011), .B2(new_n276), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n999), .A2(new_n1001), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n997), .B1(new_n991), .B2(new_n994), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1000), .B1(new_n1015), .B2(new_n1012), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1014), .A2(new_n1016), .ZN(G72));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  OAI21_X1  g833(.A(new_n1019), .B1(new_n987), .B2(new_n979), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n585), .B(KEYINPUT126), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1020), .A2(new_n583), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n586), .A2(new_n562), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n865), .A2(new_n867), .A3(new_n1019), .A4(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1023), .A2(new_n924), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1021), .A2(new_n561), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1008), .A2(new_n814), .A3(new_n980), .A4(new_n1010), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(new_n1019), .ZN(new_n1029));
  OR2_X1    g843(.A1(new_n1029), .A2(KEYINPUT127), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(KEYINPUT127), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1026), .B1(new_n1030), .B2(new_n1031), .ZN(G57));
endmodule


