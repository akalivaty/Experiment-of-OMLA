//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  OAI21_X1  g005(.A(G214), .B1(G237), .B2(G902), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT79), .B1(new_n193), .B2(G104), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G107), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(G104), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G101), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n196), .B2(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n193), .A2(KEYINPUT3), .A3(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n196), .A2(G107), .ZN(new_n207));
  AND4_X1   g021(.A1(new_n201), .A2(new_n205), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n193), .A2(G104), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(new_n203), .B2(new_n204), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n201), .B1(new_n210), .B2(new_n206), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n200), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT85), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT5), .ZN(new_n214));
  INV_X1    g028(.A(G116), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G119), .ZN(new_n216));
  INV_X1    g030(.A(G119), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G116), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT70), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(G116), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(G119), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n214), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G113), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(new_n216), .B2(new_n214), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n213), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n222), .B1(new_n220), .B2(new_n221), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(KEYINPUT85), .B(new_n226), .C1(new_n231), .C2(new_n214), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT2), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n225), .A3(KEYINPUT69), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(KEYINPUT2), .B2(G113), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n234), .A2(new_n236), .B1(KEYINPUT2), .B2(G113), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n220), .A3(new_n221), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n212), .A2(new_n228), .A3(new_n232), .A4(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(G110), .B(G122), .Z(new_n240));
  XOR2_X1   g054(.A(new_n240), .B(KEYINPUT8), .Z(new_n241));
  NAND3_X1  g055(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT5), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n226), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n239), .B(new_n241), .C1(new_n212), .C2(new_n244), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n193), .A2(KEYINPUT3), .A3(G104), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT3), .B1(new_n193), .B2(G104), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n207), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G101), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT78), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT78), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n248), .A2(new_n252), .A3(new_n249), .A4(G101), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n237), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n231), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n238), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n249), .B1(new_n248), .B2(G101), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(new_n208), .B2(new_n211), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n254), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n199), .A2(G101), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n206), .B(new_n207), .C1(new_n246), .C2(new_n247), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT77), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n210), .A2(new_n201), .A3(new_n206), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n265), .A2(new_n228), .A3(new_n232), .A4(new_n238), .ZN(new_n266));
  INV_X1    g080(.A(new_n240), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n260), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n245), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G224), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT7), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G146), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT65), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G146), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n277), .A3(G143), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n274), .A2(G143), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n278), .A2(G128), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n274), .A2(G143), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT65), .B(G146), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(G143), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n281), .B1(G143), .B2(new_n285), .ZN(new_n287));
  INV_X1    g101(.A(G128), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT68), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT1), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT67), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT67), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT1), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n288), .B1(new_n278), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n284), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n275), .A2(new_n277), .ZN(new_n298));
  INV_X1    g112(.A(G143), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n290), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n283), .B1(new_n289), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G125), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(KEYINPUT0), .A2(G128), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n278), .A2(new_n280), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(KEYINPUT0), .A2(G128), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n306), .B1(new_n300), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n273), .B1(new_n304), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n269), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n304), .A2(new_n311), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT89), .B1(new_n314), .B2(new_n272), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n304), .A2(new_n316), .A3(new_n311), .A4(new_n273), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(G902), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n260), .A2(new_n266), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT86), .A3(new_n240), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT6), .A3(new_n268), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n267), .B1(new_n260), .B2(new_n266), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(KEYINPUT86), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT87), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT6), .ZN(new_n326));
  AND4_X1   g140(.A1(new_n325), .A2(new_n320), .A3(new_n326), .A4(new_n240), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n325), .B1(new_n323), .B2(new_n326), .ZN(new_n328));
  OAI22_X1  g142(.A1(new_n322), .A2(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n271), .B(KEYINPUT88), .Z(new_n330));
  XNOR2_X1  g144(.A(new_n314), .B(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n319), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(G210), .B1(G237), .B2(G902), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n327), .A2(new_n328), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n323), .A2(KEYINPUT86), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n337), .A2(KEYINPUT6), .A3(new_n321), .A4(new_n268), .ZN(new_n338));
  INV_X1    g152(.A(new_n331), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n333), .B1(new_n340), .B2(new_n319), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n192), .B1(new_n335), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT12), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n279), .B1(new_n285), .B2(G143), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n288), .B1(new_n284), .B2(KEYINPUT1), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n282), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n344), .B1(new_n212), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n265), .A2(KEYINPUT80), .A3(new_n347), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n349), .A2(new_n350), .B1(new_n302), .B2(new_n212), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT11), .ZN(new_n352));
  INV_X1    g166(.A(G134), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n352), .B1(new_n353), .B2(G137), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(G137), .ZN(new_n355));
  INV_X1    g169(.A(G137), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT11), .A3(G134), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G131), .ZN(new_n359));
  INV_X1    g173(.A(G131), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n354), .A2(new_n357), .A3(new_n360), .A4(new_n355), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n343), .B1(new_n351), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n302), .A2(new_n212), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n263), .A2(new_n264), .ZN(new_n365));
  AND4_X1   g179(.A1(KEYINPUT80), .A2(new_n365), .A3(new_n200), .A4(new_n347), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT80), .B1(new_n265), .B2(new_n347), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n359), .A2(new_n361), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(KEYINPUT12), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n363), .A2(new_n370), .A3(KEYINPUT83), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT83), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n372), .B(new_n343), .C1(new_n351), .C2(new_n362), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G110), .B(G140), .ZN(new_n375));
  INV_X1    g189(.A(G227), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(G953), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n375), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n310), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n251), .A2(new_n253), .B1(new_n365), .B2(new_n258), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n278), .A2(new_n295), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G128), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT68), .B1(new_n383), .B2(new_n286), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n296), .A2(new_n300), .A3(new_n290), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n282), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT10), .ZN(new_n387));
  AOI211_X1 g201(.A(new_n387), .B(new_n261), .C1(new_n263), .C2(new_n264), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n380), .A2(new_n381), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n366), .B2(new_n367), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n391), .A3(new_n362), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT82), .A4(new_n362), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n374), .A2(KEYINPUT84), .A3(new_n379), .A4(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n398));
  INV_X1    g212(.A(new_n390), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(new_n349), .B2(new_n350), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n254), .A2(new_n259), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n365), .A2(KEYINPUT10), .A3(new_n200), .ZN(new_n402));
  OAI22_X1  g216(.A1(new_n401), .A2(new_n310), .B1(new_n302), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT82), .B1(new_n404), .B2(new_n362), .ZN(new_n405));
  INV_X1    g219(.A(new_n395), .ZN(new_n406));
  OAI22_X1  g220(.A1(new_n405), .A2(new_n406), .B1(new_n362), .B2(new_n404), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n398), .B1(new_n407), .B2(new_n378), .ZN(new_n408));
  AND4_X1   g222(.A1(new_n379), .A2(new_n396), .A3(new_n373), .A4(new_n371), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n397), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G469), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n190), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n373), .B(new_n371), .C1(new_n405), .C2(new_n406), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n378), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n362), .B1(new_n389), .B2(new_n391), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n394), .B2(new_n395), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n379), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(G469), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(G469), .A2(G902), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n191), .B(new_n342), .C1(new_n412), .C2(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(G119), .B(G128), .Z(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT24), .B(G110), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT23), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n217), .B2(G128), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n288), .A2(KEYINPUT23), .A3(G119), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n426), .B(new_n427), .C1(G119), .C2(new_n288), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n424), .B1(new_n428), .B2(G110), .ZN(new_n429));
  INV_X1    g243(.A(G140), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G125), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n303), .A2(G140), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n275), .A2(new_n277), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT16), .ZN(new_n434));
  OR3_X1    g248(.A1(new_n303), .A2(KEYINPUT16), .A3(G140), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(G146), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n429), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT76), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n422), .A2(new_n423), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(G110), .B2(new_n428), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n435), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT75), .A3(G146), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT75), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n274), .ZN(new_n444));
  NAND2_X1  g258(.A1(KEYINPUT75), .A2(G146), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n434), .A2(new_n435), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n440), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n438), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT22), .B(G137), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n270), .A2(G221), .A3(G234), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n449), .B(new_n450), .Z(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n438), .A2(new_n447), .A3(new_n451), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G217), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(G234), .B2(new_n190), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G902), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT25), .B1(new_n455), .B2(new_n190), .ZN(new_n460));
  AND4_X1   g274(.A1(KEYINPUT25), .A2(new_n453), .A3(new_n190), .A4(new_n454), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n457), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT32), .ZN(new_n465));
  INV_X1    g279(.A(new_n355), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n353), .A2(G137), .ZN(new_n467));
  OAI21_X1  g281(.A(G131), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n361), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n386), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT28), .ZN(new_n472));
  INV_X1    g286(.A(new_n257), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n380), .A2(new_n369), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n471), .A2(new_n472), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n473), .B(new_n474), .C1(new_n302), .C2(new_n469), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT28), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT66), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n362), .B2(new_n310), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n286), .A2(new_n308), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n369), .A2(new_n480), .A3(KEYINPUT66), .A4(new_n306), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n302), .B2(new_n469), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n475), .A2(new_n477), .B1(new_n257), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(G237), .A2(G953), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G210), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT27), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT26), .B(G101), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT31), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n386), .A2(new_n470), .B1(new_n479), .B2(new_n481), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n257), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(KEYINPUT30), .B(new_n474), .C1(new_n302), .C2(new_n469), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT71), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n471), .A2(KEYINPUT71), .A3(KEYINPUT30), .A4(new_n474), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT72), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n476), .A2(new_n500), .A3(new_n489), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n476), .B2(new_n489), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n491), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n498), .A2(new_n497), .ZN(new_n505));
  INV_X1    g319(.A(new_n493), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n473), .B1(new_n483), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n476), .A2(new_n489), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n476), .A2(new_n500), .A3(new_n489), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n512), .A3(KEYINPUT31), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n490), .B1(new_n504), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(G472), .A2(G902), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n465), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(KEYINPUT32), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT74), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n490), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n508), .A2(new_n512), .A3(KEYINPUT31), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT31), .B1(new_n508), .B2(new_n512), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT32), .A4(new_n515), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n517), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT73), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n489), .B1(new_n508), .B2(new_n476), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n475), .A2(new_n477), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n483), .A2(new_n257), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n489), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT29), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n527), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT29), .B1(new_n484), .B2(new_n489), .ZN(new_n535));
  INV_X1    g349(.A(new_n476), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n505), .B2(new_n507), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n535), .B(KEYINPUT73), .C1(new_n489), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n471), .A2(new_n474), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n257), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n529), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n489), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n532), .ZN(new_n543));
  AOI21_X1  g357(.A(G902), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n534), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G472), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n464), .B1(new_n526), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT97), .ZN(new_n548));
  XOR2_X1   g362(.A(G113), .B(G122), .Z(new_n549));
  XOR2_X1   g363(.A(KEYINPUT93), .B(G104), .Z(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G113), .B(G122), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT93), .B(G104), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n431), .A2(new_n432), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G146), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n433), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT18), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(new_n360), .ZN(new_n560));
  INV_X1    g374(.A(G237), .ZN(new_n561));
  AND4_X1   g375(.A1(G143), .A2(new_n561), .A3(new_n270), .A4(G214), .ZN(new_n562));
  AOI21_X1  g376(.A(G143), .B1(new_n485), .B2(G214), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n270), .A3(G214), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n299), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n485), .A2(G143), .A3(G214), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT90), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(new_n559), .B2(new_n360), .ZN(new_n569));
  NAND3_X1  g383(.A1(KEYINPUT90), .A2(KEYINPUT18), .A3(G131), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n566), .A2(new_n567), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n558), .A2(new_n564), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT91), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT91), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n558), .A2(new_n564), .A3(new_n571), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G131), .B1(new_n562), .B2(new_n563), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n566), .A2(new_n360), .A3(new_n567), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(G125), .B(G140), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n580), .A2(KEYINPUT92), .A3(KEYINPUT19), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT19), .B1(new_n580), .B2(KEYINPUT92), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n436), .B(new_n579), .C1(new_n583), .C2(new_n298), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n555), .B1(new_n576), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n360), .B1(new_n566), .B2(new_n567), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n442), .A2(new_n446), .B1(KEYINPUT17), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n577), .A2(new_n590), .A3(new_n578), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n573), .A2(new_n575), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n551), .A2(new_n593), .A3(new_n554), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n551), .B2(new_n554), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n587), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n588), .A2(KEYINPUT17), .ZN(new_n598));
  INV_X1    g412(.A(new_n446), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n443), .B(new_n274), .C1(new_n434), .C2(new_n435), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n591), .B(new_n598), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n576), .A2(new_n587), .A3(new_n601), .A4(new_n596), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n586), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT20), .ZN(new_n605));
  NOR2_X1   g419(.A1(G475), .A2(G902), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n604), .A2(KEYINPUT96), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n566), .A2(new_n567), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n609), .A2(new_n560), .B1(new_n557), .B2(new_n433), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n574), .B1(new_n610), .B2(new_n571), .ZN(new_n611));
  INV_X1    g425(.A(new_n575), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n601), .B(new_n596), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT95), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n602), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n586), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n608), .A2(new_n606), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n607), .B1(new_n618), .B2(KEYINPUT20), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n615), .B1(new_n592), .B2(new_n555), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n190), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G475), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n548), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n616), .B1(new_n615), .B2(new_n586), .ZN(new_n625));
  AOI211_X1 g439(.A(KEYINPUT96), .B(new_n585), .C1(new_n614), .C2(new_n602), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n605), .B1(new_n627), .B2(new_n606), .ZN(new_n628));
  OAI211_X1 g442(.A(KEYINPUT97), .B(new_n622), .C1(new_n628), .C2(new_n607), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n270), .A2(G952), .ZN(new_n631));
  NAND2_X1  g445(.A1(G234), .A2(G237), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT21), .B(G898), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n632), .A2(G902), .A3(G953), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT100), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(G116), .B(G122), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n193), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n288), .A2(G143), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n642), .A2(KEYINPUT13), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n288), .A2(G143), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n642), .B2(KEYINPUT13), .ZN(new_n645));
  OAI21_X1  g459(.A(G134), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(G128), .B(G143), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n353), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n641), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n647), .B(new_n353), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n215), .A2(KEYINPUT14), .A3(G122), .ZN(new_n652));
  INV_X1    g466(.A(new_n640), .ZN(new_n653));
  OAI211_X1 g467(.A(G107), .B(new_n652), .C1(new_n653), .C2(KEYINPUT14), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n651), .B(new_n654), .C1(G107), .C2(new_n653), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n650), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n188), .A2(new_n456), .A3(G953), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n657), .A2(new_n659), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n190), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(G478), .ZN(new_n663));
  NOR2_X1   g477(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n662), .B(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n630), .A2(new_n639), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n421), .A2(new_n547), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G101), .ZN(G3));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n514), .B2(G902), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n523), .A2(new_n515), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n523), .A2(new_n190), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT101), .B1(new_n676), .B2(G472), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n675), .A2(new_n464), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n191), .B1(new_n412), .B2(new_n420), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n342), .A2(new_n639), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n662), .A2(new_n663), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n658), .B(KEYINPUT102), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n657), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT103), .Z(new_n685));
  INV_X1    g499(.A(KEYINPUT33), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n661), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n660), .A2(new_n661), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n686), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n663), .A2(G902), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n624), .A2(new_n629), .B1(new_n682), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n681), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n680), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT34), .B(G104), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G6));
  AND4_X1   g511(.A1(new_n605), .A2(new_n608), .A3(new_n606), .A4(new_n617), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n622), .B(new_n668), .C1(new_n628), .C2(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT104), .B1(new_n699), .B2(new_n639), .ZN(new_n700));
  INV_X1    g514(.A(new_n342), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n618), .A2(KEYINPUT20), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n627), .A2(new_n605), .A3(new_n606), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n623), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n705), .A3(new_n638), .A4(new_n668), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n700), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n680), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT35), .B(G107), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G9));
  NOR2_X1   g524(.A1(new_n462), .A2(new_n463), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n452), .A2(KEYINPUT36), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n448), .B(new_n712), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n713), .A2(new_n458), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n675), .A2(new_n677), .A3(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n679), .A3(new_n701), .A4(new_n669), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT37), .B(G110), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G12));
  NAND4_X1  g533(.A1(new_n546), .A2(new_n525), .A3(new_n517), .A4(new_n519), .ZN(new_n720));
  INV_X1    g534(.A(new_n715), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n421), .A2(new_n723), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n636), .A2(G900), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n633), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n699), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n288), .ZN(G30));
  XNOR2_X1  g544(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n726), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n679), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n733), .A2(KEYINPUT40), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(KEYINPUT40), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n489), .B1(new_n540), .B2(new_n476), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n508), .B2(new_n512), .ZN(new_n737));
  OAI21_X1  g551(.A(G472), .B1(new_n737), .B2(G902), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n517), .A2(new_n519), .A3(new_n525), .A4(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n335), .A2(new_n341), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT38), .ZN(new_n741));
  INV_X1    g555(.A(new_n192), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n630), .A2(new_n668), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .A4(new_n721), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n734), .A2(new_n735), .A3(new_n739), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT106), .B(G143), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G45));
  NAND2_X1  g561(.A1(new_n692), .A2(new_n682), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n630), .A2(new_n748), .A3(new_n726), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n724), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n274), .ZN(G48));
  OAI21_X1  g566(.A(KEYINPUT84), .B1(new_n416), .B2(new_n379), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n396), .A2(new_n379), .A3(new_n373), .A4(new_n371), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(G902), .B1(new_n755), .B2(new_n397), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n411), .ZN(new_n757));
  AOI211_X1 g571(.A(G469), .B(G902), .C1(new_n755), .C2(new_n397), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n757), .A2(new_n758), .A3(new_n191), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n547), .A2(new_n759), .A3(new_n694), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT41), .B(G113), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G15));
  NAND3_X1  g576(.A1(new_n547), .A2(new_n759), .A3(new_n707), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G116), .ZN(G18));
  NAND4_X1  g578(.A1(new_n723), .A2(new_n759), .A3(new_n701), .A4(new_n669), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G119), .ZN(G21));
  NOR2_X1   g580(.A1(new_n743), .A2(new_n342), .ZN(new_n767));
  INV_X1    g581(.A(new_n673), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n504), .A2(new_n513), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n541), .A2(new_n489), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n516), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n768), .A2(new_n464), .A3(new_n771), .A4(new_n639), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n759), .A2(new_n767), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  NOR4_X1   g588(.A1(new_n757), .A2(new_n758), .A3(new_n191), .A4(new_n342), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n749), .A2(KEYINPUT107), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n693), .A2(new_n777), .A3(new_n726), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n768), .A2(new_n715), .A3(new_n771), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n775), .A2(new_n776), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G125), .ZN(G27));
  NAND2_X1  g595(.A1(new_n776), .A2(new_n778), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n332), .A2(new_n334), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n340), .A2(new_n319), .A3(new_n333), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n192), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT108), .ZN(new_n787));
  INV_X1    g601(.A(new_n191), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n784), .A2(new_n785), .A3(new_n789), .A4(new_n192), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n418), .A2(new_n419), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n756), .B2(new_n411), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n514), .A2(new_n518), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n465), .B2(new_n674), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n464), .B1(new_n796), .B2(new_n546), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n783), .A2(KEYINPUT42), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT42), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n794), .A2(new_n547), .A3(new_n776), .A4(new_n778), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n799), .B1(new_n800), .B2(KEYINPUT109), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT109), .ZN(new_n802));
  INV_X1    g616(.A(new_n464), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n720), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n804), .A2(new_n793), .A3(new_n791), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n802), .B1(new_n783), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n798), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G131), .ZN(G33));
  OAI21_X1  g622(.A(KEYINPUT110), .B1(new_n699), .B2(new_n727), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n704), .A2(new_n810), .A3(new_n668), .A4(new_n726), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n794), .A2(new_n547), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G134), .ZN(G36));
  NAND2_X1  g628(.A1(new_n414), .A2(new_n417), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT45), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n414), .A2(KEYINPUT45), .A3(new_n417), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(G469), .A3(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(new_n419), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(KEYINPUT111), .A3(KEYINPUT46), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT111), .B1(new_n820), .B2(KEYINPUT46), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n758), .B1(new_n820), .B2(KEYINPUT46), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n788), .A3(new_n732), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n624), .A2(new_n629), .A3(new_n748), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT43), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT44), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n721), .B1(new_n675), .B2(new_n677), .ZN(new_n830));
  OR3_X1    g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n787), .A2(new_n790), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n829), .B1(new_n828), .B2(new_n830), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n826), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(new_n356), .ZN(G39));
  NAND2_X1  g651(.A1(new_n825), .A2(new_n788), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT47), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n838), .B1(new_n843), .B2(new_n841), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n749), .A2(new_n832), .A3(new_n720), .A4(new_n803), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n842), .A2(new_n848), .A3(new_n844), .A4(new_n845), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(G140), .ZN(G42));
  INV_X1    g665(.A(new_n759), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n832), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n828), .A2(new_n633), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n779), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n856), .A2(KEYINPUT117), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(KEYINPUT117), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n739), .A2(new_n464), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n632), .A2(new_n853), .A3(new_n631), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n630), .A2(new_n748), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n857), .A2(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n741), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n852), .A2(new_n863), .A3(new_n192), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n768), .A2(new_n464), .A3(new_n771), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n854), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT50), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n757), .A2(new_n758), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n842), .A2(new_n844), .B1(new_n191), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n867), .A2(new_n832), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n870), .A2(new_n875), .A3(KEYINPUT51), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n855), .A2(new_n797), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT48), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n854), .A2(new_n775), .A3(new_n866), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n860), .A2(new_n693), .ZN(new_n883));
  AND4_X1   g697(.A1(new_n631), .A2(new_n881), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n878), .A2(new_n879), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n765), .A2(new_n760), .A3(new_n763), .A4(new_n773), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n794), .A2(new_n776), .A3(new_n778), .A4(new_n779), .ZN(new_n887));
  INV_X1    g701(.A(new_n668), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n704), .A2(new_n888), .A3(new_n726), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n720), .A2(new_n721), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n794), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n813), .A3(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n624), .A2(new_n629), .A3(new_n888), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n748), .B1(new_n624), .B2(new_n629), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n678), .A2(new_n895), .A3(new_n679), .A4(new_n681), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n670), .A2(new_n717), .A3(new_n896), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n886), .A2(new_n892), .A3(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n711), .A2(new_n714), .A3(new_n727), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n788), .B(new_n899), .C1(new_n758), .C2(new_n792), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT114), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT114), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n679), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n701), .A2(new_n739), .A3(new_n630), .A4(new_n668), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n723), .B(new_n421), .C1(new_n728), .C2(new_n750), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT52), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n780), .A2(new_n905), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n780), .A2(new_n905), .A3(new_n906), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT52), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n898), .A2(new_n807), .A3(new_n908), .A4(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n898), .A2(new_n807), .A3(new_n908), .A4(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n912), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n916), .A2(new_n912), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n912), .B2(new_n911), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  OAI22_X1  g738(.A1(new_n885), .A2(new_n924), .B1(G952), .B2(G953), .ZN(new_n925));
  NOR4_X1   g739(.A1(new_n863), .A2(new_n827), .A3(new_n191), .A4(new_n742), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n871), .B(KEYINPUT49), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n927), .A3(new_n859), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n925), .A2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n270), .A2(G952), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(G210), .B(G902), .C1(new_n913), .C2(new_n917), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT56), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n329), .B(KEYINPUT118), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n331), .B(KEYINPUT55), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n935), .B(new_n936), .Z(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT119), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n940), .B(new_n937), .C1(new_n932), .C2(new_n933), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n931), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(G902), .B1(new_n913), .B2(new_n917), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT120), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT120), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n945), .B(G902), .C1(new_n913), .C2(new_n917), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n334), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n938), .A2(KEYINPUT56), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT121), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n947), .A2(KEYINPUT121), .A3(new_n948), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n942), .B1(new_n951), .B2(new_n952), .ZN(G51));
  XOR2_X1   g767(.A(new_n419), .B(KEYINPUT57), .Z(new_n954));
  OR2_X1    g768(.A1(new_n916), .A2(new_n912), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n911), .A2(new_n912), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n919), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n920), .B1(KEYINPUT122), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n957), .A2(KEYINPUT122), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n410), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n944), .A2(new_n946), .ZN(new_n962));
  INV_X1    g776(.A(new_n819), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n930), .B1(new_n961), .B2(new_n964), .ZN(G54));
  AND2_X1   g779(.A1(KEYINPUT58), .A2(G475), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n962), .A2(KEYINPUT123), .A3(new_n627), .A4(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT123), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n944), .A2(new_n946), .A3(new_n966), .ZN(new_n969));
  INV_X1    g783(.A(new_n627), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n930), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n967), .A2(new_n971), .A3(new_n972), .ZN(G60));
  NAND2_X1  g787(.A1(G478), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT59), .Z(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n920), .B2(new_n923), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n688), .A2(new_n690), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n931), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n958), .A2(new_n959), .ZN(new_n979));
  INV_X1    g793(.A(new_n975), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n978), .B1(new_n979), .B2(new_n981), .ZN(G63));
  NAND2_X1  g796(.A1(G217), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT60), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n918), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n930), .B1(new_n985), .B2(new_n713), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n455), .B2(new_n985), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n985), .B2(new_n713), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(KEYINPUT61), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  OAI221_X1 g805(.A(new_n986), .B1(new_n455), .B2(new_n985), .C1(new_n989), .C2(KEYINPUT61), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(G66));
  INV_X1    g807(.A(G224), .ZN(new_n994));
  OAI21_X1  g808(.A(G953), .B1(new_n634), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n886), .A2(new_n897), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(G953), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n935), .B1(G898), .B2(new_n270), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(G69));
  OAI21_X1  g813(.A(new_n505), .B1(new_n492), .B2(new_n493), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(new_n583), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI211_X1 g816(.A(G900), .B(G953), .C1(new_n1002), .C2(G227), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(G227), .B2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n767), .A2(new_n797), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n826), .B1(new_n835), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n807), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n780), .A2(new_n906), .A3(new_n813), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n850), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(G953), .B1(new_n1010), .B2(new_n1002), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n547), .A2(new_n833), .A3(new_n895), .ZN(new_n1012));
  OAI22_X1  g826(.A1(new_n826), .A2(new_n835), .B1(new_n733), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT125), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n745), .A2(new_n780), .A3(new_n906), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT62), .Z(new_n1016));
  NAND3_X1  g830(.A1(new_n850), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n1001), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1004), .B1(new_n1011), .B2(new_n1018), .ZN(G72));
  NAND3_X1  g833(.A1(new_n850), .A2(new_n1009), .A3(new_n996), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1021));
  XNOR2_X1  g835(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1022));
  AND2_X1   g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1022), .B(new_n1023), .Z(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  AND3_X1   g839(.A1(new_n1020), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1021), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n537), .A2(new_n542), .ZN(new_n1028));
  NOR3_X1   g842(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  OR2_X1    g843(.A1(new_n886), .A2(new_n897), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1025), .B1(new_n1017), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n537), .A2(new_n542), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n528), .B1(new_n508), .B2(new_n512), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1034), .A2(new_n1024), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n930), .B1(new_n922), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1029), .A2(new_n1037), .ZN(G57));
endmodule


