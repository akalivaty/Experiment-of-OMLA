

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XOR2_X1 U322 ( .A(n358), .B(n357), .Z(n508) );
  AND2_X1 U323 ( .A1(G230GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U324 ( .A(n454), .B(KEYINPUT46), .ZN(n455) );
  XNOR2_X1 U325 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n329) );
  XNOR2_X1 U326 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U327 ( .A(n429), .B(n290), .ZN(n430) );
  XNOR2_X1 U328 ( .A(n373), .B(KEYINPUT96), .ZN(n482) );
  XNOR2_X1 U329 ( .A(n431), .B(n430), .ZN(n435) );
  INV_X1 U330 ( .A(n482), .ZN(n483) );
  XNOR2_X1 U331 ( .A(n441), .B(n440), .ZN(n442) );
  NOR2_X1 U332 ( .A1(n507), .A2(n485), .ZN(n445) );
  XNOR2_X1 U333 ( .A(n443), .B(n442), .ZN(n576) );
  INV_X1 U334 ( .A(G43GAT), .ZN(n450) );
  XNOR2_X1 U335 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U336 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U337 ( .A(n479), .B(n478), .ZN(G1351GAT) );
  XNOR2_X1 U338 ( .A(n453), .B(n452), .ZN(G1330GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT83), .B(G183GAT), .Z(n292) );
  XNOR2_X1 U340 ( .A(G15GAT), .B(G190GAT), .ZN(n291) );
  XNOR2_X1 U341 ( .A(n292), .B(n291), .ZN(n294) );
  XOR2_X1 U342 ( .A(G43GAT), .B(G99GAT), .Z(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n307) );
  XOR2_X1 U344 ( .A(G127GAT), .B(G134GAT), .Z(n296) );
  XNOR2_X1 U345 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(n297), .ZN(n356) );
  XNOR2_X1 U348 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n298), .B(KEYINPUT17), .ZN(n299) );
  XOR2_X1 U350 ( .A(n299), .B(KEYINPUT84), .Z(n301) );
  XNOR2_X1 U351 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n339) );
  XOR2_X1 U353 ( .A(n356), .B(n339), .Z(n305) );
  XOR2_X1 U354 ( .A(G71GAT), .B(G176GAT), .Z(n303) );
  XNOR2_X1 U355 ( .A(KEYINPUT20), .B(KEYINPUT82), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n309) );
  NAND2_X1 U359 ( .A1(G227GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n475) );
  INV_X1 U361 ( .A(n475), .ZN(n519) );
  XOR2_X1 U362 ( .A(KEYINPUT87), .B(KEYINPUT23), .Z(n311) );
  XOR2_X1 U363 ( .A(G50GAT), .B(G162GAT), .Z(n378) );
  XOR2_X1 U364 ( .A(G22GAT), .B(G155GAT), .Z(n393) );
  XNOR2_X1 U365 ( .A(n378), .B(n393), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U367 ( .A(n312), .B(KEYINPUT89), .Z(n318) );
  XNOR2_X1 U368 ( .A(G106GAT), .B(G78GAT), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n313), .B(G148GAT), .ZN(n437) );
  XOR2_X1 U370 ( .A(n437), .B(KEYINPUT86), .Z(n315) );
  NAND2_X1 U371 ( .A1(G228GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n316), .B(G204GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U375 ( .A(KEYINPUT22), .B(KEYINPUT90), .Z(n320) );
  XNOR2_X1 U376 ( .A(G211GAT), .B(KEYINPUT24), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U378 ( .A(n322), .B(n321), .Z(n327) );
  XNOR2_X1 U379 ( .A(G197GAT), .B(G218GAT), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n323), .B(KEYINPUT21), .ZN(n330) );
  XOR2_X1 U381 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n325) );
  XNOR2_X1 U382 ( .A(G141GAT), .B(KEYINPUT88), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n325), .B(n324), .ZN(n351) );
  XNOR2_X1 U384 ( .A(n330), .B(n351), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n472) );
  XNOR2_X1 U386 ( .A(n472), .B(KEYINPUT66), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n328), .B(KEYINPUT28), .ZN(n518) );
  XOR2_X1 U388 ( .A(G36GAT), .B(G190GAT), .Z(n385) );
  XOR2_X1 U389 ( .A(n385), .B(n331), .Z(n333) );
  NAND2_X1 U390 ( .A1(G226GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n336) );
  XOR2_X1 U392 ( .A(KEYINPUT77), .B(G211GAT), .Z(n335) );
  XNOR2_X1 U393 ( .A(G8GAT), .B(G183GAT), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n398) );
  XOR2_X1 U395 ( .A(n336), .B(n398), .Z(n341) );
  XOR2_X1 U396 ( .A(G64GAT), .B(G92GAT), .Z(n338) );
  XNOR2_X1 U397 ( .A(G176GAT), .B(G204GAT), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n436) );
  XNOR2_X1 U399 ( .A(n339), .B(n436), .ZN(n340) );
  XOR2_X1 U400 ( .A(n341), .B(n340), .Z(n342) );
  XOR2_X1 U401 ( .A(n342), .B(KEYINPUT27), .Z(n367) );
  INV_X1 U402 ( .A(n367), .ZN(n359) );
  XOR2_X1 U403 ( .A(KEYINPUT1), .B(G57GAT), .Z(n344) );
  XNOR2_X1 U404 ( .A(G1GAT), .B(G155GAT), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n344), .B(n343), .ZN(n355) );
  XOR2_X1 U406 ( .A(G85GAT), .B(G162GAT), .Z(n346) );
  XNOR2_X1 U407 ( .A(G29GAT), .B(G148GAT), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U409 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n348) );
  NAND2_X1 U410 ( .A1(G225GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U412 ( .A(n350), .B(n349), .Z(n353) );
  XNOR2_X1 U413 ( .A(n351), .B(KEYINPUT6), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n358) );
  INV_X1 U416 ( .A(n356), .ZN(n357) );
  NAND2_X1 U417 ( .A1(n359), .A2(n508), .ZN(n516) );
  NOR2_X1 U418 ( .A1(n518), .A2(n516), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n360), .B(KEYINPUT93), .ZN(n361) );
  NOR2_X1 U420 ( .A1(n519), .A2(n361), .ZN(n372) );
  XNOR2_X1 U421 ( .A(KEYINPUT25), .B(KEYINPUT95), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n362), .B(KEYINPUT94), .ZN(n365) );
  INV_X1 U423 ( .A(n342), .ZN(n467) );
  NOR2_X1 U424 ( .A1(n475), .A2(n467), .ZN(n363) );
  NOR2_X1 U425 ( .A1(n472), .A2(n363), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n369) );
  NAND2_X1 U427 ( .A1(n472), .A2(n475), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n366), .B(KEYINPUT26), .ZN(n567) );
  NOR2_X1 U429 ( .A1(n367), .A2(n567), .ZN(n368) );
  NOR2_X1 U430 ( .A1(n369), .A2(n368), .ZN(n370) );
  NOR2_X1 U431 ( .A1(n370), .A2(n508), .ZN(n371) );
  NOR2_X1 U432 ( .A1(n372), .A2(n371), .ZN(n373) );
  XOR2_X1 U433 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n375) );
  XNOR2_X1 U434 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n389) );
  XOR2_X1 U436 ( .A(G29GAT), .B(G43GAT), .Z(n377) );
  XNOR2_X1 U437 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n421) );
  XNOR2_X1 U439 ( .A(n378), .B(n421), .ZN(n380) );
  AND2_X1 U440 ( .A1(G232GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U442 ( .A(KEYINPUT9), .B(G92GAT), .Z(n382) );
  XNOR2_X1 U443 ( .A(G134GAT), .B(G106GAT), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n387) );
  XOR2_X1 U446 ( .A(G99GAT), .B(G85GAT), .Z(n429) );
  XOR2_X1 U447 ( .A(n385), .B(n429), .Z(n386) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U449 ( .A(n389), .B(n388), .Z(n532) );
  XNOR2_X1 U450 ( .A(n532), .B(KEYINPUT36), .ZN(n583) );
  NOR2_X1 U451 ( .A1(n482), .A2(n583), .ZN(n410) );
  XOR2_X1 U452 ( .A(KEYINPUT78), .B(G64GAT), .Z(n391) );
  XNOR2_X1 U453 ( .A(G127GAT), .B(G78GAT), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U455 ( .A(n393), .B(n392), .Z(n395) );
  NAND2_X1 U456 ( .A1(G231GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n397) );
  INV_X1 U458 ( .A(KEYINPUT79), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n398), .B(KEYINPUT14), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U462 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n402) );
  XNOR2_X1 U463 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n404), .B(n403), .ZN(n409) );
  XNOR2_X1 U466 ( .A(G15GAT), .B(G1GAT), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n405), .B(KEYINPUT70), .ZN(n419) );
  XOR2_X1 U468 ( .A(G57GAT), .B(KEYINPUT13), .Z(n407) );
  XNOR2_X1 U469 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n431) );
  XOR2_X1 U471 ( .A(n419), .B(n431), .Z(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n480) );
  NAND2_X1 U473 ( .A1(n410), .A2(n480), .ZN(n411) );
  XOR2_X1 U474 ( .A(KEYINPUT37), .B(n411), .Z(n507) );
  XOR2_X1 U475 ( .A(G8GAT), .B(G141GAT), .Z(n413) );
  XNOR2_X1 U476 ( .A(G197GAT), .B(G22GAT), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U478 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n415) );
  XNOR2_X1 U479 ( .A(KEYINPUT69), .B(KEYINPUT67), .ZN(n414) );
  XNOR2_X1 U480 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n428) );
  XNOR2_X1 U482 ( .A(G113GAT), .B(G50GAT), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n418), .B(G36GAT), .ZN(n420) );
  XOR2_X1 U484 ( .A(n420), .B(n419), .Z(n426) );
  XOR2_X1 U485 ( .A(n421), .B(KEYINPUT68), .Z(n423) );
  NAND2_X1 U486 ( .A1(G229GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U488 ( .A(G169GAT), .B(n424), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U490 ( .A(n428), .B(n427), .Z(n521) );
  XOR2_X1 U491 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n433) );
  XNOR2_X1 U492 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n443) );
  XOR2_X1 U495 ( .A(n437), .B(n436), .Z(n441) );
  XOR2_X1 U496 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n439) );
  XNOR2_X1 U497 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  OR2_X1 U499 ( .A1(n521), .A2(n576), .ZN(n485) );
  XNOR2_X1 U500 ( .A(KEYINPUT98), .B(KEYINPUT38), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n495) );
  NAND2_X1 U502 ( .A1(n495), .A2(n508), .ZN(n449) );
  XOR2_X1 U503 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n447) );
  INV_X1 U504 ( .A(G29GAT), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(G1328GAT) );
  NAND2_X1 U507 ( .A1(n495), .A2(n519), .ZN(n453) );
  XOR2_X1 U508 ( .A(KEYINPUT40), .B(KEYINPUT100), .Z(n451) );
  INV_X1 U509 ( .A(n532), .ZN(n549) );
  INV_X1 U510 ( .A(n521), .ZN(n570) );
  XOR2_X1 U511 ( .A(KEYINPUT41), .B(n576), .Z(n556) );
  NAND2_X1 U512 ( .A1(n570), .A2(n556), .ZN(n454) );
  INV_X1 U513 ( .A(n480), .ZN(n579) );
  XNOR2_X1 U514 ( .A(KEYINPUT103), .B(n579), .ZN(n561) );
  NAND2_X1 U515 ( .A1(n455), .A2(n561), .ZN(n456) );
  NOR2_X1 U516 ( .A1(n549), .A2(n456), .ZN(n457) );
  XOR2_X1 U517 ( .A(KEYINPUT47), .B(n457), .Z(n465) );
  NOR2_X1 U518 ( .A1(n480), .A2(n583), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n458), .B(KEYINPUT45), .ZN(n460) );
  INV_X1 U520 ( .A(KEYINPUT65), .ZN(n459) );
  XNOR2_X1 U521 ( .A(n460), .B(n459), .ZN(n462) );
  NOR2_X1 U522 ( .A1(n576), .A2(n570), .ZN(n461) );
  AND2_X1 U523 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT104), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n466), .B(KEYINPUT48), .ZN(n517) );
  NOR2_X1 U527 ( .A1(n517), .A2(n467), .ZN(n469) );
  XNOR2_X1 U528 ( .A(KEYINPUT54), .B(KEYINPUT115), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U530 ( .A1(n470), .A2(n508), .ZN(n471) );
  XOR2_X1 U531 ( .A(KEYINPUT64), .B(n471), .Z(n568) );
  NOR2_X1 U532 ( .A1(n472), .A2(n568), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n473), .B(KEYINPUT55), .ZN(n474) );
  NOR2_X2 U534 ( .A1(n475), .A2(n474), .ZN(n559) );
  NAND2_X1 U535 ( .A1(n559), .A2(n549), .ZN(n479) );
  XOR2_X1 U536 ( .A(KEYINPUT58), .B(KEYINPUT120), .Z(n477) );
  INV_X1 U537 ( .A(G190GAT), .ZN(n476) );
  NOR2_X1 U538 ( .A1(n480), .A2(n549), .ZN(n481) );
  XNOR2_X1 U539 ( .A(KEYINPUT16), .B(n481), .ZN(n484) );
  NAND2_X1 U540 ( .A1(n484), .A2(n483), .ZN(n497) );
  NOR2_X1 U541 ( .A1(n485), .A2(n497), .ZN(n492) );
  NAND2_X1 U542 ( .A1(n508), .A2(n492), .ZN(n488) );
  XOR2_X1 U543 ( .A(G1GAT), .B(KEYINPUT34), .Z(n486) );
  XNOR2_X1 U544 ( .A(KEYINPUT97), .B(n486), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n488), .B(n487), .ZN(G1324GAT) );
  NAND2_X1 U546 ( .A1(n342), .A2(n492), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n489), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .Z(n491) );
  NAND2_X1 U549 ( .A1(n492), .A2(n519), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  NAND2_X1 U551 ( .A1(n492), .A2(n518), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U553 ( .A1(n342), .A2(n495), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U555 ( .A1(n495), .A2(n518), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT101), .B(KEYINPUT42), .Z(n499) );
  NAND2_X1 U558 ( .A1(n521), .A2(n556), .ZN(n506) );
  NOR2_X1 U559 ( .A1(n506), .A2(n497), .ZN(n503) );
  NAND2_X1 U560 ( .A1(n503), .A2(n508), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(n500), .ZN(G1332GAT) );
  NAND2_X1 U563 ( .A1(n342), .A2(n503), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n501), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U565 ( .A1(n519), .A2(n503), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U567 ( .A(G78GAT), .B(KEYINPUT43), .Z(n505) );
  NAND2_X1 U568 ( .A1(n503), .A2(n518), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(G1335GAT) );
  XNOR2_X1 U570 ( .A(G85GAT), .B(KEYINPUT102), .ZN(n510) );
  NOR2_X1 U571 ( .A1(n507), .A2(n506), .ZN(n513) );
  NAND2_X1 U572 ( .A1(n513), .A2(n508), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1336GAT) );
  NAND2_X1 U574 ( .A1(n342), .A2(n513), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U576 ( .A1(n519), .A2(n513), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n518), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(KEYINPUT44), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G106GAT), .B(n515), .ZN(G1339GAT) );
  OR2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n536) );
  NOR2_X1 U582 ( .A1(n518), .A2(n536), .ZN(n520) );
  NAND2_X1 U583 ( .A1(n520), .A2(n519), .ZN(n531) );
  NOR2_X1 U584 ( .A1(n521), .A2(n531), .ZN(n523) );
  XNOR2_X1 U585 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G113GAT), .B(n524), .ZN(G1340GAT) );
  INV_X1 U588 ( .A(n556), .ZN(n525) );
  NOR2_X1 U589 ( .A1(n525), .A2(n531), .ZN(n527) );
  XNOR2_X1 U590 ( .A(KEYINPUT107), .B(KEYINPUT49), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U592 ( .A(G120GAT), .B(n528), .Z(G1341GAT) );
  NOR2_X1 U593 ( .A1(n561), .A2(n531), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT50), .B(n529), .Z(n530) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(n530), .ZN(G1342GAT) );
  NOR2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U597 ( .A(KEYINPUT108), .B(KEYINPUT51), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G134GAT), .B(n535), .ZN(G1343GAT) );
  NOR2_X1 U600 ( .A1(n567), .A2(n536), .ZN(n537) );
  XOR2_X1 U601 ( .A(KEYINPUT109), .B(n537), .Z(n548) );
  NAND2_X1 U602 ( .A1(n548), .A2(n570), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n538), .B(KEYINPUT110), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(n539), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT113), .B(KEYINPUT53), .Z(n541) );
  XNOR2_X1 U606 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n545) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n548), .A2(n556), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(G1345GAT) );
  NAND2_X1 U612 ( .A1(n579), .A2(n548), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT114), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G155GAT), .B(n547), .ZN(G1346GAT) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U617 ( .A1(n559), .A2(n570), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(KEYINPUT116), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G169GAT), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT57), .B(KEYINPUT118), .Z(n554) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U623 ( .A(KEYINPUT117), .B(n555), .Z(n558) );
  NAND2_X1 U624 ( .A1(n559), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  INV_X1 U626 ( .A(n559), .ZN(n560) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT119), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n565) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(KEYINPUT122), .B(n566), .Z(n572) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT121), .B(n569), .ZN(n582) );
  INV_X1 U636 ( .A(n582), .ZN(n580) );
  NAND2_X1 U637 ( .A1(n580), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n574) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT124), .B(n575), .Z(n578) );
  NAND2_X1 U643 ( .A1(n580), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

