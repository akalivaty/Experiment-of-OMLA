//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G125), .B(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n192), .B(G146), .C1(KEYINPUT16), .C2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  OR3_X1    g012(.A1(new_n198), .A2(KEYINPUT75), .A3(G128), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT75), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n203));
  OAI22_X1  g017(.A1(new_n200), .A2(G119), .B1(KEYINPUT74), .B2(KEYINPUT23), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n199), .B(new_n202), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G110), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT76), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n205), .A2(KEYINPUT76), .A3(new_n208), .A4(new_n206), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n198), .A2(G128), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n201), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT24), .B(G110), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n195), .B(new_n197), .C1(new_n209), .C2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G125), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G140), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n194), .A2(new_n218), .A3(KEYINPUT16), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n194), .A2(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n196), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n195), .A2(new_n221), .ZN(new_n222));
  OAI221_X1 g036(.A(new_n222), .B1(new_n212), .B2(new_n213), .C1(new_n207), .C2(new_n208), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT22), .B(G137), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G953), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(G221), .A3(G234), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n228), .B(KEYINPUT77), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT78), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n229), .A2(KEYINPUT78), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n226), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OR2_X1    g047(.A1(new_n229), .A2(KEYINPUT78), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n225), .A3(new_n230), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n224), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n233), .A2(new_n235), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n216), .A2(new_n238), .A3(new_n223), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n188), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n237), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n239), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n190), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n216), .A2(new_n238), .A3(new_n223), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n238), .B1(new_n216), .B2(new_n223), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n189), .A2(G902), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT26), .B(G101), .Z(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n252), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(G137), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT11), .A3(G134), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(G137), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n260), .A2(new_n262), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n260), .A2(new_n262), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G131), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n196), .A2(G143), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT65), .ZN(new_n272));
  INV_X1    g086(.A(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G146), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n196), .A3(G143), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT0), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(new_n200), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n272), .A2(new_n274), .A3(new_n276), .A4(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n276), .A2(new_n274), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n272), .A4(new_n278), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n278), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n271), .A2(new_n274), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n277), .A2(new_n200), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n280), .A2(new_n283), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n270), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(KEYINPUT68), .B(KEYINPUT1), .C1(new_n273), .C2(G146), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G128), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT68), .B1(new_n271), .B2(KEYINPUT1), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n286), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n281), .A2(new_n272), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n261), .A2(G134), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n264), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G131), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n267), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n290), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n198), .A2(G116), .ZN(new_n303));
  INV_X1    g117(.A(G116), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G119), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT2), .B(G113), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n307), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n302), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT69), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n301), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n267), .A2(new_n297), .A3(KEYINPUT69), .A4(new_n300), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n314), .A2(new_n290), .A3(new_n315), .A4(new_n310), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT28), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n302), .B2(new_n311), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n257), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n265), .A2(new_n266), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n265), .A2(new_n266), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n323), .A2(new_n324), .B1(G131), .B2(new_n299), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n270), .A2(new_n289), .B1(new_n325), .B2(new_n297), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n311), .B1(new_n326), .B2(KEYINPUT30), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT70), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT69), .B1(new_n325), .B2(new_n297), .ZN(new_n330));
  INV_X1    g144(.A(new_n315), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n270), .B2(new_n289), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n329), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n314), .A3(new_n329), .A4(new_n315), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n328), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n316), .A2(new_n257), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT31), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n314), .A2(new_n290), .A3(KEYINPUT30), .A4(new_n315), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT70), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n327), .B1(new_n343), .B2(new_n336), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT31), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n344), .A2(new_n345), .A3(new_n339), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n322), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(G472), .A2(G902), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n251), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n338), .A2(KEYINPUT31), .A3(new_n340), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n345), .B1(new_n344), .B2(new_n339), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n321), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n353));
  INV_X1    g167(.A(new_n348), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n314), .A2(new_n315), .A3(new_n290), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n311), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n319), .B1(new_n358), .B2(new_n316), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n320), .A2(KEYINPUT29), .A3(new_n257), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n188), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n257), .ZN(new_n362));
  INV_X1    g176(.A(new_n316), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n362), .B1(new_n344), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT28), .B1(new_n326), .B2(new_n310), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(new_n362), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n318), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n361), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT73), .A3(G472), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT73), .ZN(new_n371));
  INV_X1    g185(.A(G472), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n371), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n250), .B1(new_n356), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT9), .B(G234), .ZN(new_n376));
  OAI21_X1  g190(.A(G221), .B1(new_n376), .B2(G902), .ZN(new_n377));
  XOR2_X1   g191(.A(new_n377), .B(KEYINPUT79), .Z(new_n378));
  NAND2_X1  g192(.A1(new_n227), .A2(G227), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT80), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G140), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G107), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G104), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(G104), .B2(new_n383), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n384), .A2(new_n385), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT82), .B1(new_n383), .B2(G104), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G107), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n390), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n383), .A2(KEYINPUT81), .A3(G104), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n383), .A2(KEYINPUT81), .A3(KEYINPUT3), .A4(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n395), .A2(new_n400), .A3(KEYINPUT84), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT84), .B1(new_n395), .B2(new_n400), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n389), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT86), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT86), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n389), .B(new_n405), .C1(new_n401), .C2(new_n402), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT10), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(new_n294), .B2(new_n296), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT87), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n404), .A2(KEYINPUT87), .A3(new_n406), .A4(new_n408), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n270), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n390), .A2(new_n393), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT83), .B1(new_n400), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n400), .A2(new_n415), .A3(KEYINPUT83), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(G101), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT4), .B1(new_n401), .B2(new_n402), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n417), .A2(KEYINPUT4), .A3(G101), .A4(new_n418), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n281), .A2(new_n272), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n271), .A2(KEYINPUT1), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n424), .B1(new_n200), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n296), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n427), .B(new_n389), .C1(new_n402), .C2(new_n401), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n423), .A2(new_n289), .B1(new_n407), .B2(new_n428), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n413), .A2(new_n414), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n414), .B1(new_n413), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n382), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT88), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n428), .A2(new_n407), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n418), .A2(G101), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n436), .A2(new_n437), .A3(new_n416), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n420), .B2(new_n419), .ZN(new_n439));
  INV_X1    g253(.A(new_n289), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(new_n411), .B2(new_n412), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n382), .B1(new_n442), .B2(new_n414), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n403), .A2(new_n296), .A3(new_n294), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n414), .B1(new_n428), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT12), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g261(.A(KEYINPUT88), .B(new_n382), .C1(new_n430), .C2(new_n431), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n434), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G469), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n188), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n413), .A2(new_n429), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n270), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n413), .A2(new_n414), .A3(new_n429), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n446), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n443), .A2(new_n453), .B1(new_n455), .B2(new_n382), .ZN(new_n456));
  OAI21_X1  g270(.A(G469), .B1(new_n456), .B2(G902), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n378), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G214), .B1(G237), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n294), .A2(new_n296), .A3(new_n217), .ZN(new_n461));
  INV_X1    g275(.A(G224), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(G953), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT89), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT7), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n461), .B(new_n466), .C1(new_n289), .C2(new_n217), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT91), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n440), .A2(G125), .B1(KEYINPUT90), .B2(new_n461), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n461), .A2(KEYINPUT90), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G122), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n472), .B(KEYINPUT8), .Z(new_n473));
  NAND3_X1  g287(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT5), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(G113), .C1(KEYINPUT5), .C2(new_n303), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n308), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n403), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n403), .A2(new_n476), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n468), .A2(new_n471), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n476), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n404), .A2(new_n406), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n482), .B(new_n472), .C1(new_n439), .C2(new_n310), .ZN(new_n483));
  AOI21_X1  g297(.A(G902), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n472), .ZN(new_n485));
  INV_X1    g299(.A(new_n482), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n310), .B1(new_n421), .B2(new_n422), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(KEYINPUT6), .A3(new_n483), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n490), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n461), .B1(new_n289), .B2(new_n217), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(new_n464), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n484), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G210), .B1(G237), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n484), .A2(new_n494), .A3(new_n496), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n460), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G237), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n227), .A3(G214), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(new_n273), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n253), .B(G214), .C1(KEYINPUT92), .C2(G143), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n263), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT17), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n507), .A2(new_n221), .A3(new_n195), .ZN(new_n508));
  INV_X1    g322(.A(new_n506), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n263), .A3(new_n505), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n504), .A2(new_n505), .ZN(new_n513));
  NAND2_X1  g327(.A1(KEYINPUT18), .A2(G131), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n513), .A2(new_n515), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n194), .A2(new_n218), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G146), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n519), .A2(new_n197), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n508), .A2(new_n512), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(G113), .B(G122), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(new_n392), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT93), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n517), .ZN(new_n529));
  INV_X1    g343(.A(new_n520), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n516), .ZN(new_n531));
  INV_X1    g345(.A(new_n511), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n532), .A2(KEYINPUT17), .A3(new_n506), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n507), .A2(new_n221), .A3(new_n195), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n526), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n528), .A2(new_n188), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G475), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n524), .B1(new_n521), .B2(new_n516), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n191), .A2(KEYINPUT19), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n191), .A2(KEYINPUT19), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI221_X1 g356(.A(new_n195), .B1(new_n532), .B2(new_n506), .C1(G146), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(G475), .A2(G902), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n544), .B(new_n545), .C1(new_n522), .C2(new_n525), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(KEYINPUT20), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT20), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n535), .A2(new_n524), .B1(new_n539), .B2(new_n543), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n549), .B2(new_n545), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n538), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n273), .A2(G128), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n200), .A2(G143), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(new_n259), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n304), .A2(KEYINPUT14), .A3(G122), .ZN(new_n558));
  XNOR2_X1  g372(.A(G116), .B(G122), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(G107), .B(new_n558), .C1(new_n560), .C2(KEYINPUT14), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n557), .B(new_n561), .C1(G107), .C2(new_n560), .ZN(new_n562));
  INV_X1    g376(.A(new_n554), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n563), .A2(KEYINPUT13), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n555), .B1(new_n563), .B2(KEYINPUT13), .ZN(new_n565));
  OAI21_X1  g379(.A(G134), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n556), .A2(new_n259), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n559), .B(new_n383), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n376), .A2(new_n187), .A3(G953), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n562), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n562), .B2(new_n569), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n188), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G478), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n562), .A2(new_n569), .ZN(new_n577));
  INV_X1    g391(.A(new_n570), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n562), .A2(new_n569), .A3(new_n570), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n575), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n188), .A3(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n576), .A2(new_n583), .A3(KEYINPUT95), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT95), .B1(new_n576), .B2(new_n583), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n538), .B(KEYINPUT94), .C1(new_n547), .C2(new_n550), .ZN(new_n587));
  NOR2_X1   g401(.A1(KEYINPUT96), .A2(G952), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(KEYINPUT96), .A2(G952), .ZN(new_n590));
  AOI21_X1  g404(.A(G953), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G234), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(new_n501), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n188), .B(new_n227), .C1(G234), .C2(G237), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT21), .B(G898), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AND4_X1   g412(.A1(new_n553), .A2(new_n586), .A3(new_n587), .A4(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n375), .A2(new_n458), .A3(new_n500), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  OAI21_X1  g415(.A(G472), .B1(new_n352), .B2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n347), .A2(new_n348), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n458), .A2(new_n249), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n498), .A2(new_n499), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n459), .A3(new_n598), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT97), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT33), .B1(new_n570), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n581), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n610), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n579), .B2(new_n580), .ZN(new_n613));
  OAI21_X1  g427(.A(G478), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n581), .A2(new_n574), .A3(new_n188), .ZN(new_n615));
  NAND2_X1  g429(.A1(G478), .A2(G902), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n553), .B2(new_n587), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n606), .A2(new_n608), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT99), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT34), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(new_n547), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n546), .A2(KEYINPUT20), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n627), .B2(KEYINPUT100), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n629), .B(KEYINPUT101), .C1(new_n546), .C2(KEYINPUT20), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n625), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT101), .B1(new_n550), .B2(new_n629), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n627), .A2(KEYINPUT100), .A3(new_n626), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n547), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n631), .A2(new_n538), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n576), .A2(new_n583), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT95), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n576), .A2(new_n583), .A3(KEYINPUT95), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n635), .A2(new_n636), .A3(new_n641), .A4(new_n598), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n631), .A2(new_n641), .A3(new_n634), .A4(new_n538), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT102), .B1(new_n643), .B2(new_n597), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n642), .A2(new_n500), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n606), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT103), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n224), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n248), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT104), .B1(new_n244), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(KEYINPUT25), .B1(new_n247), .B2(new_n188), .ZN(new_n656));
  INV_X1    g470(.A(new_n243), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n189), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n659), .A3(new_n653), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n459), .A2(new_n607), .A3(new_n655), .A4(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n458), .A2(new_n661), .A3(new_n599), .A4(new_n605), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  INV_X1    g478(.A(new_n251), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n603), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n347), .A2(KEYINPUT32), .A3(new_n348), .ZN(new_n667));
  INV_X1    g481(.A(new_n373), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n368), .A2(new_n371), .A3(new_n372), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n666), .B(new_n667), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n593), .ZN(new_n671));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n671), .B1(new_n672), .B2(new_n594), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n643), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n458), .A2(new_n661), .A3(new_n670), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT105), .B(G128), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G30));
  NAND2_X1  g491(.A1(new_n338), .A2(new_n316), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n362), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n358), .A2(new_n316), .A3(new_n362), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n188), .ZN(new_n682));
  OAI21_X1  g496(.A(G472), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n356), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n607), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n498), .A2(new_n499), .A3(new_n686), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n553), .A2(new_n587), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n641), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n658), .A2(new_n653), .ZN(new_n693));
  OR3_X1    g507(.A1(new_n692), .A2(new_n693), .A3(new_n460), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n685), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n673), .B(KEYINPUT39), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n458), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT40), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n458), .A2(new_n699), .A3(new_n696), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n695), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  AOI211_X1 g516(.A(new_n673), .B(new_n617), .C1(new_n553), .C2(new_n587), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n458), .A2(new_n661), .A3(new_n670), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  INV_X1    g519(.A(new_n451), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n450), .B1(new_n449), .B2(new_n188), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n620), .A2(new_n608), .ZN(new_n709));
  INV_X1    g523(.A(new_n378), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n375), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT107), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT41), .B(G113), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NAND4_X1  g528(.A1(new_n708), .A2(new_n375), .A3(new_n645), .A4(new_n710), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  NAND3_X1  g530(.A1(new_n599), .A2(new_n660), .A3(new_n655), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n356), .B2(new_n374), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n708), .A2(new_n718), .A3(new_n710), .A4(new_n500), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  OAI21_X1  g534(.A(new_n362), .B1(new_n359), .B2(new_n365), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n341), .B2(new_n346), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n348), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n602), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n724), .A2(new_n249), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n608), .A2(new_n692), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n708), .A2(new_n725), .A3(new_n710), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  NAND2_X1  g542(.A1(new_n449), .A2(new_n188), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G469), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n710), .A3(new_n451), .A4(new_n500), .ZN(new_n731));
  AND4_X1   g545(.A1(new_n602), .A2(new_n703), .A3(new_n723), .A4(new_n693), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n217), .ZN(G27));
  NAND4_X1  g549(.A1(new_n498), .A2(new_n710), .A3(new_n459), .A4(new_n499), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n451), .B2(new_n457), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n375), .A2(new_n703), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n451), .A2(new_n457), .ZN(new_n742));
  INV_X1    g556(.A(new_n736), .ZN(new_n743));
  INV_X1    g557(.A(new_n673), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n618), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n739), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n742), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n668), .A2(new_n669), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n353), .B1(new_n352), .B2(new_n354), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n667), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n249), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n741), .B1(new_n747), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n737), .A2(new_n746), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n754), .A2(new_n751), .A3(KEYINPUT108), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n740), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  NAND4_X1  g571(.A1(new_n737), .A2(new_n670), .A3(new_n249), .A4(new_n674), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n455), .A2(new_n382), .ZN(new_n761));
  INV_X1    g575(.A(new_n382), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n453), .A2(new_n762), .A3(new_n454), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n760), .B1(new_n764), .B2(new_n450), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n456), .A2(KEYINPUT45), .ZN(new_n766));
  OAI211_X1 g580(.A(KEYINPUT109), .B(G469), .C1(new_n456), .C2(KEYINPUT45), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(G469), .A2(G902), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n768), .A2(KEYINPUT46), .A3(new_n769), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n451), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT43), .B1(new_n691), .B2(new_n617), .ZN(new_n775));
  INV_X1    g589(.A(new_n617), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n553), .A4(new_n587), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(KEYINPUT44), .A3(new_n604), .A4(new_n693), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n775), .A2(new_n693), .A3(new_n778), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n605), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n498), .A2(new_n459), .A3(new_n499), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n780), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n774), .A2(new_n786), .A3(new_n710), .A4(new_n696), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  NOR4_X1   g602(.A1(new_n670), .A2(new_n249), .A3(new_n745), .A4(new_n784), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n706), .B1(new_n770), .B2(new_n771), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n790), .B(new_n378), .C1(new_n791), .C2(new_n773), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT47), .B1(new_n774), .B2(new_n710), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT110), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n768), .A2(KEYINPUT46), .A3(new_n769), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT46), .B1(new_n768), .B2(new_n769), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n796), .A2(new_n797), .A3(new_n706), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n790), .B1(new_n798), .B2(new_n378), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n774), .A2(KEYINPUT47), .A3(new_n710), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n789), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  NAND4_X1  g619(.A1(new_n711), .A2(new_n715), .A3(new_n719), .A4(new_n662), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n553), .A2(new_n587), .A3(new_n637), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT112), .B1(new_n807), .B2(new_n618), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n807), .A2(KEYINPUT112), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n608), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n458), .A3(new_n249), .A4(new_n605), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n727), .A3(new_n600), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n737), .A2(new_n732), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n637), .A2(new_n673), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n635), .A2(new_n660), .A3(new_n655), .A4(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n784), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n458), .A2(new_n670), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n758), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n758), .A2(new_n818), .A3(new_n814), .A4(KEYINPUT113), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n813), .A2(new_n756), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n692), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n693), .A2(new_n673), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n500), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n458), .A2(new_n827), .A3(new_n684), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n704), .A2(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n731), .A2(new_n733), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(KEYINPUT114), .A3(new_n675), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n675), .B1(new_n731), .B2(new_n733), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n704), .A2(new_n828), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n833), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n839), .B2(new_n829), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n824), .A2(new_n838), .A3(KEYINPUT53), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n831), .A2(new_n835), .A3(KEYINPUT52), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n662), .A2(new_n715), .A3(new_n711), .A4(new_n719), .ZN(new_n846));
  INV_X1    g660(.A(new_n812), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n823), .A2(new_n756), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(new_n831), .B2(new_n835), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n845), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n842), .B(new_n843), .C1(new_n850), .C2(KEYINPUT53), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT115), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n824), .A2(new_n838), .A3(KEYINPUT53), .A4(new_n844), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n848), .A2(new_n849), .A3(new_n840), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(KEYINPUT53), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT54), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n824), .A2(new_n838), .A3(new_n844), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n843), .A4(new_n842), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n591), .B(KEYINPUT117), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n725), .A2(new_n779), .A3(new_n671), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n736), .A2(new_n593), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n685), .A2(new_n708), .A3(new_n249), .A4(new_n864), .ZN(new_n865));
  OAI221_X1 g679(.A(new_n862), .B1(new_n863), .B2(new_n731), .C1(new_n865), .C2(new_n620), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n708), .A2(new_n779), .A3(new_n864), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n752), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n868), .A2(KEYINPUT48), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(KEYINPUT48), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n863), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n730), .A2(new_n451), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n378), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT116), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT50), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n459), .B1(new_n688), .B2(new_n689), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n872), .A2(new_n874), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n708), .A2(new_n878), .A3(new_n710), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n875), .B(new_n876), .C1(new_n880), .C2(new_n863), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n724), .A2(new_n693), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n867), .A2(new_n883), .ZN(new_n884));
  OR3_X1    g698(.A1(new_n865), .A2(new_n691), .A3(new_n776), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n799), .B(new_n800), .C1(new_n710), .C2(new_n873), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n863), .A2(new_n784), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n871), .B1(new_n889), .B2(KEYINPUT51), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n891), .B(new_n886), .C1(new_n887), .C2(new_n888), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n852), .A2(new_n856), .A3(new_n861), .A4(new_n893), .ZN(new_n894));
  OR2_X1    g708(.A1(G952), .A2(G953), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n691), .A2(new_n617), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n249), .A3(new_n710), .A4(new_n459), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n873), .B2(KEYINPUT49), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT111), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n873), .A2(KEYINPUT49), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n685), .A3(new_n690), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT118), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n896), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n227), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n859), .A2(new_n842), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(G902), .ZN(new_n911));
  INV_X1    g725(.A(G210), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n489), .A2(new_n491), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n493), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT55), .Z(new_n916));
  AOI21_X1  g730(.A(new_n908), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n188), .B1(new_n859), .B2(new_n842), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT56), .B1(new_n918), .B2(G210), .ZN(new_n919));
  INV_X1    g733(.A(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n917), .A2(KEYINPUT119), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n923));
  INV_X1    g737(.A(new_n921), .ZN(new_n924));
  INV_X1    g738(.A(new_n908), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n919), .B2(new_n920), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n923), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n922), .A2(new_n927), .ZN(G51));
  NAND2_X1  g742(.A1(new_n910), .A2(KEYINPUT54), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(KEYINPUT120), .A3(new_n851), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n910), .A2(new_n931), .A3(KEYINPUT54), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n769), .B(KEYINPUT57), .Z(new_n933));
  NAND3_X1  g747(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n449), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n911), .A2(new_n768), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n908), .B1(new_n935), .B2(new_n936), .ZN(G54));
  AND3_X1   g751(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n938), .A2(new_n549), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n549), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n908), .ZN(G60));
  NOR2_X1   g755(.A1(new_n611), .A2(new_n613), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n616), .B(KEYINPUT59), .ZN(new_n943));
  AND4_X1   g757(.A1(new_n942), .A2(new_n930), .A3(new_n932), .A4(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n852), .A2(new_n856), .A3(new_n861), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n942), .B1(new_n945), .B2(new_n943), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n944), .A2(new_n908), .A3(new_n946), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n859), .B2(new_n842), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n652), .B(KEYINPUT122), .Z(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n952), .B(new_n925), .C1(new_n247), .C2(new_n950), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n953), .A2(KEYINPUT121), .A3(KEYINPUT61), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT61), .B1(new_n953), .B2(KEYINPUT121), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(G66));
  OAI21_X1  g770(.A(G953), .B1(new_n595), .B2(new_n462), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n813), .B2(G953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n914), .B1(G898), .B2(new_n227), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G69));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n784), .B1(new_n809), .B2(new_n808), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n375), .A2(new_n458), .A3(new_n962), .A4(new_n696), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n787), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n695), .A2(new_n698), .A3(new_n700), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n830), .A2(new_n675), .A3(new_n704), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n839), .A2(new_n701), .A3(KEYINPUT62), .A4(new_n704), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n802), .B1(new_n801), .B2(new_n789), .ZN(new_n971));
  INV_X1    g785(.A(new_n789), .ZN(new_n972));
  AOI211_X1 g786(.A(KEYINPUT110), .B(new_n972), .C1(new_n799), .C2(new_n800), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n970), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT124), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n970), .B(new_n976), .C1(new_n971), .C2(new_n973), .ZN(new_n977));
  AOI21_X1  g791(.A(G953), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI22_X1  g792(.A1(new_n343), .A2(new_n336), .B1(new_n333), .B2(new_n302), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(new_n542), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT123), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n961), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n977), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n976), .B1(new_n804), .B2(new_n970), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n227), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(KEYINPUT125), .A3(new_n981), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n227), .A2(G900), .ZN(new_n989));
  INV_X1    g803(.A(new_n758), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n967), .A2(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n752), .A2(new_n500), .A3(new_n825), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n992), .A2(new_n710), .A3(new_n696), .A4(new_n774), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n991), .A2(new_n993), .A3(new_n756), .A4(new_n787), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n804), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n989), .B1(new_n996), .B2(new_n227), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n980), .B1(new_n997), .B2(KEYINPUT127), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n994), .B1(new_n795), .B2(new_n803), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(G953), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n999), .B1(new_n1001), .B2(new_n989), .ZN(new_n1002));
  AOI21_X1  g816(.A(KEYINPUT126), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n227), .B1(G227), .B2(G900), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n988), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1004), .B1(new_n988), .B2(new_n1003), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1005), .A2(new_n1006), .ZN(G72));
  AND2_X1   g821(.A1(new_n1000), .A2(new_n813), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n679), .B(new_n362), .C1(new_n1008), .C2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n364), .B1(new_n344), .B2(new_n339), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n855), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1012), .A2(new_n925), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n975), .A2(new_n813), .A3(new_n977), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n1010), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1015), .B1(new_n680), .B2(new_n1017), .ZN(G57));
endmodule


