//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1302,
    new_n1303, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1397, new_n1398, new_n1399, new_n1400;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AND3_X1   g0015(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n216));
  AOI21_X1  g0016(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n203), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n227), .A2(new_n228), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n212), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n215), .B(new_n222), .C1(new_n234), .C2(KEYINPUT1), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n250), .B(new_n251), .Z(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n249), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT77), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G222), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G223), .A3(G1698), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n260), .B(new_n266), .C1(new_n225), .C2(new_n265), .ZN(new_n267));
  AND2_X1   g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n218), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G1), .A2(G13), .ZN(new_n271));
  OAI21_X1  g0071(.A(G274), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n276), .A2(new_n273), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n274), .B1(G226), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n270), .A2(G190), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(KEYINPUT68), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n218), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n210), .A2(new_n262), .A3(KEYINPUT69), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT69), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(G20), .B2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n210), .A2(G33), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n285), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n284), .A2(new_n218), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n209), .A2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G50), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT70), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n298), .ZN(new_n305));
  INV_X1    g0105(.A(G50), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n297), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT9), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n308), .A2(KEYINPUT9), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n255), .B(new_n279), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n270), .A2(new_n278), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G200), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n311), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n309), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n255), .B1(new_n317), .B2(new_n279), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT10), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT76), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT10), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n314), .A2(new_n322), .A3(new_n279), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n316), .A2(new_n309), .A3(KEYINPUT76), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n313), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(KEYINPUT71), .A3(new_n308), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(G179), .B2(new_n313), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT71), .B1(new_n328), .B2(new_n308), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n294), .A2(new_n225), .B1(new_n210), .B2(G68), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(G50), .B2(new_n289), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT64), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n271), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n282), .B2(new_n283), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT11), .ZN(new_n342));
  OR3_X1    g0142(.A1(new_n336), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n336), .B2(new_n341), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n305), .A2(new_n202), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT12), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n300), .A2(G68), .A3(new_n301), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n343), .A2(new_n344), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G274), .ZN(new_n349));
  AND2_X1   g0149(.A1(G1), .A2(G13), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n275), .ZN(new_n351));
  INV_X1    g0151(.A(new_n273), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n276), .A2(new_n273), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n224), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n357));
  INV_X1    g0157(.A(G232), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G1698), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n265), .B(new_n359), .C1(G226), .C2(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G97), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n340), .A2(new_n275), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n356), .B(new_n357), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n360), .B2(new_n361), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT13), .B1(new_n365), .B2(new_n355), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(G179), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n357), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n365), .B2(new_n355), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n327), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI211_X1 g0172(.A(KEYINPUT14), .B(new_n327), .C1(new_n364), .C2(new_n369), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n348), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n364), .B2(new_n369), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(new_n348), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n364), .A2(G190), .A3(new_n366), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n378), .A2(KEYINPUT79), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(KEYINPUT79), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n374), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G1698), .ZN(new_n383));
  OAI211_X1 g0183(.A(G223), .B(new_n383), .C1(new_n256), .C2(new_n257), .ZN(new_n384));
  OAI211_X1 g0184(.A(G226), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G87), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n269), .ZN(new_n388));
  INV_X1    g0188(.A(G179), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n277), .A2(G232), .B1(new_n351), .B2(new_n352), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(G169), .B1(new_n388), .B2(new_n390), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n265), .B2(G20), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n202), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(G58), .B(G68), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n289), .A2(G159), .B1(new_n399), .B2(G20), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n394), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n258), .B2(new_n210), .ZN(new_n403));
  NOR4_X1   g0203(.A1(new_n256), .A2(new_n257), .A3(new_n395), .A4(G20), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n400), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n402), .A2(new_n285), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n295), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n299), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n301), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n298), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT80), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT80), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n409), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n393), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT18), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n354), .A2(new_n358), .B1(new_n272), .B2(new_n273), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n269), .B2(new_n387), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n421), .B2(G169), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n409), .A2(new_n414), .A3(new_n411), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n414), .B1(new_n409), .B2(new_n411), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n402), .A2(new_n285), .A3(new_n406), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n388), .A2(G190), .A3(new_n390), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n375), .B1(new_n388), .B2(new_n390), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(new_n425), .A3(new_n426), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n432), .A2(new_n425), .A3(new_n426), .A4(KEYINPUT17), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n418), .A2(new_n429), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n265), .A2(G238), .A3(G1698), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n206), .B2(new_n265), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n259), .A2(G232), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT72), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT72), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n259), .A2(new_n442), .A3(G232), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n439), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(new_n363), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n274), .B1(G244), .B2(new_n277), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G200), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(G190), .B(new_n446), .C1(new_n444), .C2(new_n363), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n301), .A2(G77), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n299), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT75), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n305), .A2(new_n225), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT74), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n408), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n455));
  INV_X1    g0255(.A(G87), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT15), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G87), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT73), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT73), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n457), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n455), .B1(new_n464), .B2(new_n294), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n454), .B1(new_n465), .B2(new_n285), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n448), .A2(new_n449), .A3(new_n452), .A4(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n327), .B1(new_n445), .B2(new_n447), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n452), .A2(new_n466), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n389), .B(new_n446), .C1(new_n444), .C2(new_n363), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  OR3_X1    g0272(.A1(new_n382), .A2(new_n437), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n334), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT84), .ZN(new_n476));
  INV_X1    g0276(.A(G45), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G1), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n481), .A2(new_n276), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT83), .B1(new_n481), .B2(new_n272), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT5), .B(G41), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n351), .A2(new_n484), .A3(new_n485), .A4(new_n478), .ZN(new_n486));
  AOI22_X1  g0286(.A1(G257), .A2(new_n482), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(G244), .B(new_n383), .C1(new_n256), .C2(new_n257), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G283), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n262), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G250), .A2(G1698), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT4), .A2(G244), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(G1698), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n492), .B1(new_n265), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n490), .A2(new_n496), .A3(KEYINPUT82), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n269), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT82), .B1(new_n490), .B2(new_n496), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n487), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n327), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT6), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n502), .A2(new_n205), .A3(G107), .ZN(new_n503));
  XNOR2_X1  g0303(.A(G97), .B(G107), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n505), .A2(new_n210), .B1(new_n225), .B2(new_n290), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n206), .B1(new_n396), .B2(new_n397), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n285), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n209), .A2(G33), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n284), .A2(new_n218), .A3(new_n298), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G97), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n305), .A2(G97), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT81), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT81), .ZN(new_n515));
  AOI211_X1 g0315(.A(new_n515), .B(new_n512), .C1(new_n510), .C2(G97), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n508), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n490), .A2(new_n496), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT82), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(new_n269), .A3(new_n497), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(new_n389), .A3(new_n487), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n501), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n500), .A2(new_n375), .ZN(new_n524));
  INV_X1    g0324(.A(G190), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n487), .B(new_n525), .C1(new_n498), .C2(new_n499), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n517), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n476), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n504), .A2(new_n502), .ZN(new_n529));
  INV_X1    g0329(.A(new_n503), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(G20), .B1(G77), .B2(new_n289), .ZN(new_n532));
  OAI21_X1  g0332(.A(G107), .B1(new_n403), .B2(new_n404), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n341), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n514), .ZN(new_n535));
  INV_X1    g0335(.A(new_n516), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n526), .ZN(new_n538));
  AOI21_X1  g0338(.A(G200), .B1(new_n521), .B2(new_n487), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n501), .A2(new_n517), .A3(new_n522), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(KEYINPUT84), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G244), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n543));
  OAI211_X1 g0343(.A(G238), .B(new_n383), .C1(new_n256), .C2(new_n257), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G116), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n269), .ZN(new_n547));
  OAI221_X1 g0347(.A(G250), .B1(G1), .B2(new_n477), .C1(new_n268), .C2(new_n271), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n276), .A2(G274), .A3(new_n478), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n551), .A3(new_n389), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT85), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n510), .ZN(new_n555));
  INV_X1    g0355(.A(new_n463), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n462), .B1(new_n457), .B2(new_n459), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT86), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT86), .B1(new_n461), .B2(new_n463), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n210), .B1(new_n361), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(G87), .B2(new_n207), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n210), .B(G68), .C1(new_n256), .C2(new_n257), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n562), .B1(new_n294), .B2(new_n205), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(new_n285), .B1(new_n464), .B2(new_n305), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n550), .B1(new_n269), .B2(new_n546), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(KEYINPUT85), .A3(new_n389), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n547), .A2(new_n551), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n327), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n554), .A2(new_n569), .A3(new_n571), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n375), .B1(new_n547), .B2(new_n551), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n570), .A2(G190), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n555), .A2(G87), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n568), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n528), .A2(new_n542), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n482), .A2(G264), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n483), .A2(new_n486), .ZN(new_n584));
  OR2_X1    g0384(.A1(G250), .A2(G1698), .ZN(new_n585));
  INV_X1    g0385(.A(G257), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G1698), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n587), .C1(new_n256), .C2(new_n257), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT88), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n269), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n583), .B(new_n584), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n375), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n588), .A2(new_n590), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT88), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n269), .A3(new_n591), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n598), .A2(new_n525), .A3(new_n584), .A4(new_n583), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n545), .A2(G20), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT23), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n210), .B2(G107), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT22), .ZN(new_n606));
  AOI21_X1  g0406(.A(G20), .B1(new_n263), .B2(new_n264), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(G87), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n210), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(KEYINPUT22), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n605), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT24), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT24), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n613), .B(new_n605), .C1(new_n608), .C2(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n285), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n305), .A2(new_n206), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n617), .B(KEYINPUT25), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n510), .A2(new_n206), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n600), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n598), .A2(new_n389), .A3(new_n584), .A4(new_n583), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n594), .A2(new_n327), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n341), .B1(new_n612), .B2(new_n614), .ZN(new_n624));
  INV_X1    g0424(.A(new_n620), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n341), .A2(G116), .A3(new_n298), .A4(new_n509), .ZN(new_n628));
  INV_X1    g0428(.A(G116), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n305), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(G20), .B1(G33), .B2(G283), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n262), .A2(G97), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n631), .A2(new_n632), .B1(G20), .B2(new_n629), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n285), .A2(KEYINPUT20), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT20), .B1(new_n285), .B2(new_n633), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n628), .B(new_n630), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n256), .A2(new_n257), .A3(G303), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n586), .A2(new_n383), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(G264), .B2(new_n383), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n637), .B1(new_n265), .B2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n640), .A2(new_n269), .B1(new_n483), .B2(new_n486), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n481), .A2(G270), .A3(new_n276), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT87), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n481), .A2(KEYINPUT87), .A3(G270), .A4(new_n276), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n636), .A2(new_n647), .A3(KEYINPUT21), .A4(G169), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n636), .A2(G179), .A3(new_n646), .A4(new_n641), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n636), .A2(new_n647), .A3(G169), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT21), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(G200), .ZN(new_n654));
  INV_X1    g0454(.A(new_n636), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n641), .A2(G190), .A3(new_n646), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n650), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  NOR4_X1   g0458(.A1(new_n475), .A2(new_n582), .A3(new_n627), .A4(new_n658), .ZN(G372));
  XNOR2_X1  g0459(.A(new_n427), .B(KEYINPUT18), .ZN(new_n660));
  INV_X1    g0460(.A(new_n471), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n381), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(new_n374), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n435), .A2(new_n436), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n660), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n332), .B1(new_n666), .B2(new_n326), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n653), .A2(new_n649), .A3(new_n648), .ZN(new_n668));
  INV_X1    g0468(.A(new_n626), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n568), .A2(new_n578), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n575), .B1(G190), .B2(new_n570), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n561), .A2(new_n568), .B1(new_n572), .B2(new_n327), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n671), .A2(new_n672), .B1(new_n673), .B2(new_n552), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n540), .A2(new_n674), .A3(new_n621), .A4(new_n541), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n523), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT26), .B1(new_n580), .B2(new_n541), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n552), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n667), .B1(new_n475), .B2(new_n682), .ZN(G369));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT89), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT89), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n668), .A2(new_n636), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n636), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n650), .A2(new_n653), .A3(new_n657), .A4(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n684), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n669), .A2(new_n693), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n693), .B1(new_n624), .B2(new_n625), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n621), .A2(new_n626), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n693), .B1(new_n650), .B2(new_n653), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n621), .A2(new_n626), .ZN(new_n704));
  INV_X1    g0504(.A(new_n693), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n703), .A2(new_n704), .B1(new_n669), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n702), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n213), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n220), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n650), .A2(new_n626), .A3(new_n653), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n523), .A2(new_n527), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(new_n717), .A3(new_n621), .A4(new_n674), .ZN(new_n718));
  AOI211_X1 g0518(.A(KEYINPUT29), .B(new_n693), .C1(new_n715), .C2(new_n718), .ZN(new_n719));
  AND4_X1   g0519(.A1(new_n541), .A2(new_n540), .A3(new_n674), .A4(new_n621), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT92), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n668), .B2(new_n669), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n650), .A2(KEYINPUT92), .A3(new_n626), .A4(new_n653), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n677), .B1(new_n580), .B2(new_n541), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT91), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n523), .A2(new_n674), .A3(KEYINPUT26), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT91), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n728), .B(new_n677), .C1(new_n580), .C2(new_n541), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n724), .A2(new_n730), .A3(new_n680), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n705), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n719), .B1(new_n732), .B2(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n482), .A2(G257), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n584), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n497), .A2(new_n269), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(new_n520), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n641), .A2(G179), .A3(new_n646), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n598), .A2(new_n570), .A3(new_n583), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n737), .A2(new_n738), .A3(new_n739), .A4(KEYINPUT30), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n570), .B(KEYINPUT90), .ZN(new_n744));
  AOI21_X1  g0544(.A(G179), .B1(new_n641), .B2(new_n646), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n744), .A2(new_n500), .A3(new_n594), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n742), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n693), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n747), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n751));
  AND4_X1   g0551(.A1(new_n653), .A2(new_n657), .A3(new_n649), .A4(new_n648), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(new_n704), .A3(new_n705), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n750), .B(new_n751), .C1(new_n582), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G330), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n733), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n714), .B1(new_n756), .B2(G1), .ZN(G364));
  INV_X1    g0557(.A(new_n697), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n694), .A2(new_n696), .A3(new_n684), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n210), .A2(G13), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n209), .B1(new_n760), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n758), .B(new_n759), .C1(new_n709), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n694), .A2(new_n696), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n218), .B1(G20), .B2(new_n327), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n525), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n210), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G97), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n210), .A2(new_n389), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(new_n525), .A3(G200), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n773), .B1(new_n202), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT94), .ZN(new_n777));
  INV_X1    g0577(.A(new_n774), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n525), .A2(new_n375), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n779), .A2(G77), .B1(new_n782), .B2(G50), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT32), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n210), .A2(G179), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(new_n525), .A3(new_n375), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n784), .B1(new_n787), .B2(G159), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n786), .A2(KEYINPUT32), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n785), .A2(new_n525), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n206), .ZN(new_n792));
  NOR4_X1   g0592(.A1(new_n788), .A2(new_n790), .A3(new_n258), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n780), .A2(new_n785), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n456), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n778), .A2(new_n525), .A3(G200), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(G58), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n777), .A2(new_n783), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G303), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  OAI22_X1  g0601(.A1(new_n775), .A2(new_n801), .B1(new_n791), .B2(new_n491), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n800), .B(new_n802), .C1(G311), .C2(new_n779), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n772), .A2(G294), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n265), .B1(new_n782), .B2(G326), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n796), .A2(G322), .B1(G329), .B2(new_n787), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n769), .B1(new_n798), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n709), .A2(new_n762), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT93), .Z(new_n810));
  NOR2_X1   g0610(.A1(new_n708), .A2(new_n258), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G355), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(G116), .B2(new_n213), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n708), .A2(new_n265), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(new_n477), .B2(new_n221), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n253), .A2(G45), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n813), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n768), .A2(new_n766), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n810), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n808), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n767), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n763), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NAND4_X1  g0625(.A1(new_n468), .A2(new_n469), .A3(new_n470), .A4(new_n705), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n449), .A2(new_n452), .A3(new_n466), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n827), .A2(new_n448), .B1(new_n469), .B2(new_n693), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n826), .B1(new_n828), .B2(new_n661), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n682), .B2(new_n693), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n467), .A2(new_n471), .A3(new_n705), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n676), .B2(new_n681), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n809), .B1(new_n834), .B2(new_n755), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n755), .B2(new_n834), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n769), .A2(new_n765), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n810), .B1(G77), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n775), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n839), .A2(G150), .B1(new_n782), .B2(G137), .ZN(new_n840));
  INV_X1    g0640(.A(G143), .ZN(new_n841));
  INV_X1    g0641(.A(new_n796), .ZN(new_n842));
  INV_X1    g0642(.A(new_n779), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n840), .B1(new_n841), .B2(new_n842), .C1(new_n789), .C2(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT95), .Z(new_n845));
  OR2_X1    g0645(.A1(new_n845), .A2(KEYINPUT34), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(KEYINPUT34), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n202), .A2(new_n791), .B1(new_n794), .B2(new_n306), .ZN(new_n848));
  INV_X1    g0648(.A(G132), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n265), .B1(new_n786), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT96), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n848), .B(new_n851), .C1(G58), .C2(new_n772), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n846), .A2(new_n847), .A3(new_n852), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n775), .A2(new_n491), .B1(new_n791), .B2(new_n456), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n265), .B(new_n854), .C1(G311), .C2(new_n787), .ZN(new_n855));
  INV_X1    g0655(.A(new_n794), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G303), .A2(new_n782), .B1(new_n856), .B2(G107), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G116), .A2(new_n779), .B1(new_n796), .B2(G294), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n855), .A2(new_n773), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n838), .B1(new_n860), .B2(new_n768), .ZN(new_n861));
  INV_X1    g0661(.A(new_n826), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n469), .A2(new_n693), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n467), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n862), .B1(new_n864), .B2(new_n471), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n861), .B1(new_n765), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n836), .A2(new_n866), .ZN(G384));
  OR2_X1    g0667(.A1(new_n531), .A2(KEYINPUT35), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n531), .A2(KEYINPUT35), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n868), .A2(G116), .A3(new_n219), .A4(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(KEYINPUT97), .B(KEYINPUT36), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n870), .B(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n221), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n306), .A2(G68), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n209), .B(G13), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n374), .A2(new_n693), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n425), .A2(new_n426), .B1(new_n422), .B2(new_n691), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT37), .B1(new_n878), .B2(KEYINPUT99), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n432), .A2(new_n425), .A3(new_n426), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n878), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n691), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n407), .A2(new_n416), .B1(new_n393), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT99), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n884), .B(new_n433), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT100), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n691), .B1(new_n425), .B2(new_n426), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n437), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n884), .A2(new_n433), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n884), .A2(new_n885), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT37), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT100), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n887), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n889), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n880), .A2(new_n878), .A3(new_n886), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT37), .B1(new_n884), .B2(new_n433), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n891), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n904));
  NAND3_X1  g0704(.A1(new_n899), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n890), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n660), .B2(new_n664), .ZN(new_n907));
  INV_X1    g0707(.A(new_n901), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n898), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n903), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT39), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n877), .B1(new_n905), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n693), .A2(new_n348), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n382), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n374), .A2(new_n381), .A3(new_n916), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n831), .B1(new_n715), .B2(new_n718), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT98), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n921), .A2(new_n922), .A3(new_n862), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT98), .B1(new_n833), .B2(new_n826), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n912), .B(new_n920), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n660), .A2(new_n883), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n915), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT29), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n731), .B2(new_n705), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n474), .B1(new_n930), .B2(new_n719), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n667), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n928), .B(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n829), .B1(new_n919), .B2(new_n918), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT102), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n747), .A2(new_n935), .A3(new_n693), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(new_n747), .B2(new_n693), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT31), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n751), .B1(new_n582), .B2(new_n753), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n891), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n897), .B2(new_n898), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n747), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n528), .A2(new_n542), .A3(new_n581), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n658), .A2(new_n627), .A3(new_n693), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n748), .A2(KEYINPUT102), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n747), .A2(new_n935), .A3(new_n693), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n950), .A2(new_n749), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n912), .A3(new_n934), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n942), .A2(new_n945), .B1(new_n954), .B2(new_n941), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n474), .A2(new_n953), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n684), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n933), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n209), .B2(new_n760), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n933), .A2(new_n958), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n876), .B1(new_n960), .B2(new_n961), .ZN(G367));
  NAND4_X1  g0762(.A1(new_n668), .A2(new_n626), .A3(new_n621), .A4(new_n705), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n693), .A2(new_n517), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n540), .A2(new_n541), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n523), .A2(new_n693), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT42), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n964), .A2(KEYINPUT42), .A3(new_n968), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n541), .B1(new_n966), .B2(new_n626), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n970), .A2(new_n971), .B1(new_n705), .B2(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n705), .A2(new_n671), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(new_n680), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n674), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT103), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n973), .A2(KEYINPUT104), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n972), .A2(new_n705), .ZN(new_n983));
  INV_X1    g0783(.A(new_n971), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n981), .B(new_n983), .C1(new_n984), .C2(new_n969), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT104), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n989));
  OR3_X1    g0789(.A1(new_n973), .A2(new_n981), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n968), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n702), .A2(new_n991), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n988), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n992), .B1(new_n988), .B2(new_n990), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n709), .B(KEYINPUT41), .Z(new_n996));
  XNOR2_X1  g0796(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n706), .B2(new_n968), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n669), .A2(new_n705), .ZN(new_n1000));
  AND4_X1   g0800(.A1(new_n1000), .A2(new_n968), .A3(new_n963), .A4(new_n998), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n706), .B2(new_n968), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n963), .A2(new_n1000), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n991), .A2(new_n1006), .A3(new_n1003), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT107), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n702), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT108), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n668), .A2(new_n705), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(new_n698), .A3(new_n700), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n963), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n758), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n963), .B(new_n1013), .C1(new_n697), .C2(KEYINPUT108), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n997), .B1(new_n991), .B2(new_n1006), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n706), .A2(new_n968), .A3(new_n998), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1021), .A2(new_n1007), .A3(new_n1005), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n702), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(KEYINPUT107), .A3(new_n1023), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n756), .A2(new_n1010), .A3(new_n1018), .A4(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n996), .B1(new_n1025), .B2(new_n756), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n995), .B1(new_n1026), .B2(new_n762), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n819), .B1(new_n213), .B2(new_n464), .C1(new_n815), .C2(new_n243), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n810), .A2(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n842), .A2(new_n799), .B1(new_n843), .B2(new_n491), .ZN(new_n1030));
  INV_X1    g0830(.A(G311), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1031), .A2(new_n781), .B1(new_n791), .B2(new_n205), .ZN(new_n1032));
  INV_X1    g0832(.A(G317), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n258), .B1(new_n786), .B2(new_n1033), .C1(new_n771), .C2(new_n206), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT109), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n856), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT46), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n794), .B2(new_n629), .ZN(new_n1039));
  INV_X1    g0839(.A(G294), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1037), .B(new_n1039), .C1(new_n1040), .C2(new_n775), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1035), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1041), .A2(new_n1036), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n842), .A2(new_n291), .B1(new_n781), .B2(new_n841), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n225), .A2(new_n791), .B1(new_n794), .B2(new_n201), .ZN(new_n1045));
  INV_X1    g0845(.A(G137), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n265), .B1(new_n786), .B2(new_n1046), .C1(new_n771), .C2(new_n202), .ZN(new_n1047));
  OR3_X1    g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n779), .A2(G50), .B1(new_n839), .B2(G159), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT110), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1042), .A2(new_n1043), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT47), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1029), .B1(new_n1052), .B2(new_n768), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n975), .A2(new_n976), .A3(new_n766), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1027), .A2(new_n1055), .ZN(G387));
  NAND2_X1  g0856(.A1(new_n733), .A2(new_n755), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n1017), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n733), .A2(new_n755), .A3(new_n1018), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n709), .A3(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G150), .A2(new_n787), .B1(new_n856), .B2(G77), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1061), .B(new_n265), .C1(new_n205), .C2(new_n791), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT112), .Z(new_n1063));
  OAI21_X1  g0863(.A(new_n772), .B1(new_n559), .B2(new_n560), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n779), .A2(G68), .B1(new_n782), .B2(G159), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n796), .A2(G50), .B1(new_n839), .B2(new_n408), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n772), .A2(G283), .B1(new_n856), .B2(G294), .ZN(new_n1068));
  INV_X1    g0868(.A(G322), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n775), .A2(new_n1031), .B1(new_n781), .B2(new_n1069), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1070), .A2(KEYINPUT113), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(KEYINPUT113), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G303), .A2(new_n779), .B1(new_n796), .B2(G317), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT48), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1068), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT114), .Z(new_n1077));
  NAND2_X1  g0877(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1077), .A2(KEYINPUT49), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n265), .B1(new_n787), .B2(G326), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n629), .C2(new_n791), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT49), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1067), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n768), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n810), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n766), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n701), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n711), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n811), .A2(new_n1088), .B1(new_n206), .B2(new_n708), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n240), .A2(new_n477), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1091));
  OR3_X1    g0891(.A1(new_n1091), .A2(G50), .A3(new_n295), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1091), .B1(G50), .B2(new_n295), .ZN(new_n1093));
  AOI21_X1  g0893(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1092), .A2(new_n711), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n814), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1089), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1085), .B(new_n1087), .C1(new_n819), .C2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1084), .A2(new_n1098), .B1(new_n1018), .B2(new_n762), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1060), .A2(new_n1099), .ZN(G393));
  OAI21_X1  g0900(.A(new_n1023), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1021), .A2(new_n702), .A3(new_n1007), .A4(new_n1005), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1101), .A2(new_n762), .A3(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n796), .A2(G159), .B1(new_n782), .B2(G150), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT51), .Z(new_n1105));
  AOI22_X1  g0905(.A1(new_n779), .A2(new_n408), .B1(G68), .B2(new_n856), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G50), .A2(new_n839), .B1(new_n787), .B2(G143), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n771), .A2(new_n225), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n265), .B1(new_n791), .B2(new_n456), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n796), .A2(G311), .B1(new_n782), .B2(G317), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT52), .Z(new_n1113));
  AOI22_X1  g0913(.A1(new_n779), .A2(G294), .B1(G283), .B2(new_n856), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G303), .A2(new_n839), .B1(new_n787), .B2(G322), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n265), .B(new_n792), .C1(G116), .C2(new_n772), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n769), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n249), .A2(new_n814), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n820), .B1(G97), .B2(new_n708), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1085), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n968), .B2(new_n1086), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1103), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1059), .A2(new_n1125), .A3(KEYINPUT115), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT115), .B1(new_n1059), .B2(new_n1125), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1025), .A2(new_n709), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1124), .B1(new_n1128), .B2(new_n1129), .ZN(G390));
  AOI21_X1  g0930(.A(new_n684), .B1(new_n949), .B2(new_n952), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n474), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n931), .A2(new_n667), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n754), .A2(G330), .A3(new_n865), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n920), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n953), .A2(G330), .A3(new_n934), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n922), .B1(new_n921), .B2(new_n862), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n833), .A2(KEYINPUT98), .A3(new_n826), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(G330), .B(new_n865), .C1(new_n938), .C2(new_n939), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1135), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n864), .A2(new_n471), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n731), .A2(new_n705), .A3(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n754), .A2(G330), .A3(new_n865), .A4(new_n920), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1144), .A2(new_n826), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1133), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1135), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n877), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n913), .B(new_n905), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1146), .A2(new_n826), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n920), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n944), .A2(new_n1151), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1152), .A2(new_n1156), .A3(new_n1147), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n877), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n944), .A2(new_n904), .B1(KEYINPUT39), .B2(new_n912), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1159), .A2(new_n1160), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1149), .B(new_n1157), .C1(new_n1161), .C2(new_n1137), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1162), .A2(new_n709), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n934), .A2(new_n1131), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1141), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n920), .B1(new_n1131), .B2(new_n865), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1147), .A2(new_n826), .A3(new_n1146), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n1164), .A2(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n931), .A2(new_n667), .A3(new_n1132), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT116), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1170), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1157), .B1(new_n1161), .B2(new_n1137), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT117), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1149), .A2(new_n1170), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1167), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1144), .A2(new_n1177), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1178));
  OAI21_X1  g0978(.A(KEYINPUT116), .B1(new_n1178), .B2(new_n1133), .ZN(new_n1179));
  AND4_X1   g0979(.A1(KEYINPUT117), .A2(new_n1174), .A3(new_n1176), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1163), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1174), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n762), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1160), .A2(new_n764), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n810), .B1(new_n408), .B2(new_n837), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT118), .Z(new_n1186));
  NOR2_X1   g0986(.A1(new_n794), .A2(new_n291), .ZN(new_n1187));
  XOR2_X1   g0987(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1188));
  XNOR2_X1  g0988(.A(new_n1187), .B(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G128), .A2(new_n782), .B1(new_n787), .B2(G125), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n306), .C2(new_n791), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n779), .A2(new_n1193), .B1(new_n839), .B2(G137), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n258), .B1(new_n796), .B2(G132), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(new_n789), .C2(new_n771), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G107), .A2(new_n839), .B1(new_n787), .B2(G294), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n205), .B2(new_n843), .C1(new_n629), .C2(new_n842), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n491), .A2(new_n781), .B1(new_n791), .B2(new_n202), .ZN(new_n1199));
  OR4_X1    g0999(.A1(new_n265), .A2(new_n1199), .A3(new_n1108), .A4(new_n795), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n1191), .A2(new_n1196), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1186), .B1(new_n768), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1184), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1183), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1181), .A2(new_n1205), .ZN(G378));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1162), .B2(new_n1169), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT122), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n883), .A2(new_n308), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n334), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n326), .A2(new_n333), .A3(new_n1210), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1214), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1210), .B1(new_n326), .B2(new_n333), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1211), .B(new_n332), .C1(new_n319), .C2(new_n325), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n955), .B2(G330), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n374), .A2(new_n381), .A3(new_n916), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n916), .B1(new_n374), .B2(new_n381), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n865), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n949), .B2(new_n952), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n894), .A2(new_n887), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1226), .A2(KEYINPUT100), .B1(new_n437), .B2(new_n890), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT38), .B1(new_n1227), .B2(new_n896), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1225), .B(KEYINPUT40), .C1(new_n1228), .C2(new_n943), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT38), .B1(new_n891), .B2(new_n902), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n943), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n941), .B1(new_n940), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(new_n1232), .A3(G330), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1220), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n928), .B1(new_n1221), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n925), .A2(new_n926), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(new_n914), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1220), .A2(new_n1229), .A3(G330), .A4(new_n1232), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1209), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(KEYINPUT122), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1208), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT121), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1239), .A2(new_n1240), .B1(new_n915), .B2(new_n927), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1236), .A2(KEYINPUT121), .A3(new_n1241), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1248), .A2(new_n1249), .B1(new_n1169), .B2(new_n1162), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n709), .B(new_n1245), .C1(new_n1250), .C2(KEYINPUT57), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n809), .B1(new_n837), .B2(G50), .ZN(new_n1252));
  INV_X1    g1052(.A(G128), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n842), .A2(new_n1253), .B1(new_n775), .B2(new_n849), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n779), .A2(G137), .B1(new_n782), .B2(G125), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n794), .B2(new_n1192), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(G150), .C2(new_n772), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT59), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1260));
  INV_X1    g1060(.A(G41), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n262), .B(new_n1261), .C1(new_n791), .C2(new_n789), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G124), .B2(new_n787), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1259), .A2(new_n1260), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G50), .B1(new_n262), .B2(new_n1261), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n265), .B2(G41), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1261), .B(new_n258), .C1(new_n794), .C2(new_n225), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n775), .A2(new_n205), .B1(new_n791), .B2(new_n201), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1267), .B(new_n1268), .C1(G68), .C2(new_n772), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n779), .B1(new_n559), .B2(new_n560), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n782), .A2(G116), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n796), .A2(G107), .B1(G283), .B2(new_n787), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT58), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1264), .A2(new_n1266), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1252), .B1(new_n1275), .B2(new_n768), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1220), .B2(new_n765), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT120), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1279), .B2(new_n762), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1251), .A2(new_n1280), .ZN(G375));
  OAI21_X1  g1081(.A(new_n265), .B1(new_n791), .B2(new_n201), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n842), .A2(new_n1046), .B1(new_n843), .B2(new_n291), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1282), .B(new_n1283), .C1(G50), .C2(new_n772), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n775), .A2(new_n1192), .B1(new_n781), .B2(new_n849), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n1253), .A2(new_n786), .B1(new_n794), .B2(new_n789), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n842), .A2(new_n491), .B1(new_n794), .B2(new_n205), .ZN(new_n1288));
  OAI22_X1  g1088(.A1(new_n843), .A2(new_n206), .B1(new_n781), .B2(new_n1040), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n775), .A2(new_n629), .B1(new_n786), .B2(new_n799), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n258), .B1(new_n791), .B2(new_n225), .ZN(new_n1291));
  NOR4_X1   g1091(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1284), .A2(new_n1287), .B1(new_n1292), .B2(new_n1064), .ZN(new_n1293));
  OAI221_X1 g1093(.A(new_n810), .B1(G68), .B2(new_n837), .C1(new_n1293), .C2(new_n769), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n1135), .B2(new_n764), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1168), .B2(new_n762), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1178), .A2(new_n1133), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n996), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1296), .B1(new_n1297), .B2(new_n1300), .ZN(G381));
  NAND3_X1  g1101(.A1(new_n1060), .A2(new_n824), .A3(new_n1099), .ZN(new_n1302));
  OR4_X1    g1102(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1302), .ZN(new_n1303));
  OR4_X1    g1103(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1303), .ZN(G407));
  NAND2_X1  g1104(.A1(new_n692), .A2(G213), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(G375), .A2(G378), .A3(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT123), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1309));
  OAI211_X1 g1109(.A(G213), .B(G407), .C1(new_n1308), .C2(new_n1309), .ZN(G409));
  INV_X1    g1110(.A(KEYINPUT125), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1302), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n824), .B1(new_n1060), .B2(new_n1099), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1311), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1027), .A2(new_n1055), .A3(G390), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G390), .B1(new_n1027), .B2(new_n1055), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1314), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(G390), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n988), .A2(new_n990), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n992), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n988), .A2(new_n990), .A3(new_n992), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1010), .A2(new_n1024), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1324), .A2(new_n1059), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1299), .B1(new_n1325), .B2(new_n1057), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1323), .B1(new_n1326), .B2(new_n761), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1055), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1318), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G393), .A2(G396), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(KEYINPUT125), .A3(new_n1302), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1314), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1027), .A2(G390), .A3(new_n1055), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1329), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1317), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT60), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1298), .B1(new_n1149), .B2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1178), .A2(KEYINPUT60), .A3(new_n1133), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1338), .A2(new_n709), .A3(new_n1339), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(G384), .B(KEYINPUT124), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1296), .A3(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  AND2_X1   g1143(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1344), .B1(new_n1340), .B2(new_n1296), .ZN(new_n1345));
  INV_X1    g1145(.A(G2897), .ZN(new_n1346));
  OAI22_X1  g1146(.A1(new_n1343), .A2(new_n1345), .B1(new_n1346), .B2(new_n1305), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1305), .A2(new_n1346), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1340), .A2(new_n1296), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1342), .B(new_n1348), .C1(new_n1349), .C2(new_n1344), .ZN(new_n1350));
  AND2_X1   g1150(.A1(new_n1347), .A2(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1251), .A2(G378), .A3(new_n1280), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1353));
  NOR3_X1   g1153(.A1(new_n1243), .A2(new_n1247), .A3(new_n1246), .ZN(new_n1354));
  AOI21_X1  g1154(.A(KEYINPUT121), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1355));
  OAI211_X1 g1155(.A(new_n1299), .B(new_n1353), .C1(new_n1354), .C2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1278), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n762), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1356), .A2(new_n1357), .A3(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT117), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1360), .B1(new_n1297), .B2(new_n1182), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1173), .A2(KEYINPUT117), .A3(new_n1174), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1204), .B1(new_n1363), .B2(new_n1163), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1359), .A2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1352), .A2(new_n1365), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1351), .B1(new_n1366), .B2(new_n1305), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT61), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1305), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1370), .B1(new_n1352), .B2(new_n1365), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT62), .ZN(new_n1372));
  NOR2_X1   g1172(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1371), .A2(new_n1372), .A3(new_n1373), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1368), .A2(new_n1369), .A3(new_n1374), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1372), .B1(new_n1371), .B2(new_n1373), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1336), .B1(new_n1375), .B2(new_n1376), .ZN(new_n1377));
  INV_X1    g1177(.A(KEYINPUT127), .ZN(new_n1378));
  OAI211_X1 g1178(.A(KEYINPUT63), .B(new_n1342), .C1(new_n1349), .C2(new_n1344), .ZN(new_n1379));
  AOI211_X1 g1179(.A(new_n1370), .B(new_n1379), .C1(new_n1352), .C2(new_n1365), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT126), .ZN(new_n1381));
  AOI21_X1  g1181(.A(new_n1381), .B1(new_n1335), .B2(new_n1369), .ZN(new_n1382));
  AOI211_X1 g1182(.A(KEYINPUT126), .B(KEYINPUT61), .C1(new_n1317), .C2(new_n1334), .ZN(new_n1383));
  NOR2_X1   g1183(.A1(new_n1382), .A2(new_n1383), .ZN(new_n1384));
  NOR3_X1   g1184(.A1(new_n1367), .A2(new_n1380), .A3(new_n1384), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1366), .A2(new_n1305), .A3(new_n1373), .ZN(new_n1386));
  INV_X1    g1186(.A(KEYINPUT63), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1386), .A2(new_n1387), .ZN(new_n1388));
  AOI21_X1  g1188(.A(new_n1378), .B1(new_n1385), .B2(new_n1388), .ZN(new_n1389));
  INV_X1    g1189(.A(new_n1379), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1335), .A2(new_n1369), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1391), .A2(KEYINPUT126), .ZN(new_n1392));
  NAND3_X1  g1192(.A1(new_n1335), .A2(new_n1381), .A3(new_n1369), .ZN(new_n1393));
  AOI22_X1  g1193(.A1(new_n1371), .A2(new_n1390), .B1(new_n1392), .B2(new_n1393), .ZN(new_n1394));
  AND4_X1   g1194(.A1(new_n1378), .A2(new_n1394), .A3(new_n1388), .A4(new_n1368), .ZN(new_n1395));
  OAI21_X1  g1195(.A(new_n1377), .B1(new_n1389), .B2(new_n1395), .ZN(G405));
  INV_X1    g1196(.A(new_n1352), .ZN(new_n1397));
  AOI21_X1  g1197(.A(G378), .B1(new_n1251), .B2(new_n1280), .ZN(new_n1398));
  NOR2_X1   g1198(.A1(new_n1397), .A2(new_n1398), .ZN(new_n1399));
  XNOR2_X1  g1199(.A(new_n1399), .B(new_n1373), .ZN(new_n1400));
  XNOR2_X1  g1200(.A(new_n1400), .B(new_n1335), .ZN(G402));
endmodule


