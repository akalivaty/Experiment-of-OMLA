//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1142,
    new_n1143;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT64), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT65), .Z(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT66), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(new_n473), .A3(G125), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n470), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n472), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n477));
  OR2_X1    g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n476), .A2(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n468), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT67), .Z(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT68), .B1(new_n468), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n472), .A2(new_n485), .A3(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n483), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n482), .A2(new_n488), .A3(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n483), .ZN(new_n492));
  OR2_X1    g067(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n492), .A2(KEYINPUT69), .A3(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n465), .A2(new_n467), .A3(G126), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n483), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n464), .A2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G102), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(G166));
  AOI22_X1  g097(.A1(new_n516), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n509), .A2(new_n511), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n519), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n525), .B1(G51), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT7), .Z(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(G168));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n517), .A2(new_n532), .B1(new_n519), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n524), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n534), .B1(G651), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g113(.A(new_n538), .B(KEYINPUT70), .Z(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  XOR2_X1   g115(.A(KEYINPUT71), .B(G43), .Z(new_n541));
  AND2_X1   g116(.A1(new_n526), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n514), .ZN(new_n544));
  INV_X1    g119(.A(new_n517), .ZN(new_n545));
  AOI211_X1 g120(.A(new_n542), .B(new_n544), .C1(G81), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  INV_X1    g127(.A(G91), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n512), .A2(new_n516), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n553), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n512), .A2(G65), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n514), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n562), .A2(KEYINPUT72), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n562), .B2(KEYINPUT72), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND2_X1  g144(.A1(new_n554), .A2(new_n556), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G87), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT74), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n512), .A2(G74), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(G49), .B2(new_n526), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n570), .A2(new_n575), .A3(G87), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n572), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n572), .A2(new_n576), .A3(KEYINPUT75), .A4(new_n574), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n524), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  INV_X1    g161(.A(G48), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(new_n519), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n570), .B2(G86), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n526), .A2(G47), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI221_X1 g170(.A(new_n593), .B1(new_n594), .B2(new_n517), .C1(new_n514), .C2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n570), .A2(G92), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT10), .Z(new_n599));
  AOI22_X1  g174(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT77), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G54), .B2(new_n526), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n597), .B1(new_n604), .B2(G868), .ZN(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NOR2_X1   g187(.A1(new_n603), .A2(G559), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT78), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n472), .A2(new_n502), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT79), .B(KEYINPUT13), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n487), .A2(G123), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n480), .A2(G135), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(KEYINPUT80), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(KEYINPUT80), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n626), .B(new_n627), .C1(G111), .C2(new_n483), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n623), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2096), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT81), .Z(G156));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2435), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2438), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2451), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n645), .A2(G14), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2067), .B(G2678), .Z(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT17), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n648), .B2(new_n649), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n651), .B1(new_n650), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT84), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT20), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n670), .A2(new_n662), .A3(new_n665), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n668), .B(new_n671), .C1(new_n662), .C2(new_n670), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT22), .B(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G229));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G25), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n487), .A2(G119), .B1(G131), .B2(new_n480), .ZN(new_n682));
  OR2_X1    g257(.A1(G95), .A2(G2105), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n683), .B(G2104), .C1(G107), .C2(new_n483), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n681), .B1(new_n686), .B2(new_n680), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT35), .B(G1991), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT85), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G24), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT86), .Z(new_n694));
  XOR2_X1   g269(.A(G290), .B(KEYINPUT87), .Z(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(new_n692), .ZN(new_n696));
  INV_X1    g271(.A(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n591), .A2(G16), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G6), .B2(G16), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT32), .B(G1981), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n699), .B(new_n701), .C1(G6), .C2(G16), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G22), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G166), .B2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G1971), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n703), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n577), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G16), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G16), .B2(G23), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT33), .B(G1976), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(KEYINPUT34), .B1(new_n710), .B2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n713), .B(new_n714), .Z(new_n717));
  INV_X1    g292(.A(KEYINPUT34), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n717), .A2(new_n709), .A3(new_n718), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n691), .B(new_n698), .C1(new_n716), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT36), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n710), .A2(KEYINPUT34), .A3(new_n715), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n718), .B1(new_n717), .B2(new_n709), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n724), .A2(new_n725), .A3(new_n691), .A4(new_n698), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G29), .A2(G35), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G162), .B2(G29), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT29), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(G2090), .Z(new_n731));
  AND2_X1   g306(.A1(new_n692), .A2(G4), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n603), .B2(G16), .ZN(new_n733));
  INV_X1    g308(.A(G1348), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(G299), .A2(G16), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n692), .A2(KEYINPUT23), .A3(G20), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT23), .ZN(new_n738));
  INV_X1    g313(.A(G20), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(G16), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G1956), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G1961), .ZN(new_n744));
  NAND2_X1  g319(.A1(G301), .A2(G16), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n692), .A2(G5), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n743), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(G28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(G28), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n750), .A2(new_n751), .A3(new_n680), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n735), .A2(new_n748), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G29), .A2(G32), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n502), .A2(G105), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT26), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G141), .B2(new_n480), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n760));
  AND3_X1   g335(.A1(new_n487), .A2(new_n760), .A3(G129), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n760), .B1(new_n487), .B2(G129), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n756), .B(new_n759), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT92), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n755), .B1(new_n764), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT93), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT27), .B(G1996), .Z(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n692), .A2(G19), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n546), .B2(new_n692), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1341), .Z(new_n772));
  NAND2_X1  g347(.A1(G115), .A2(G2104), .ZN(new_n773));
  INV_X1    g348(.A(G127), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n468), .B2(new_n774), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n775), .A2(G2105), .B1(new_n480), .B2(G139), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n502), .A2(G103), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G33), .B(new_n780), .S(G29), .Z(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G2072), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n772), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G34), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(G29), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G160), .B2(G29), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(G2084), .ZN(new_n788));
  NOR2_X1   g363(.A1(G164), .A2(new_n680), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G27), .B2(new_n680), .ZN(new_n790));
  INV_X1    g365(.A(G2078), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT31), .B(G11), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n790), .B2(new_n791), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n783), .A2(new_n788), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n680), .A2(G26), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n480), .A2(G140), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT88), .ZN(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n483), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n487), .B2(G128), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n796), .B1(new_n804), .B2(new_n680), .ZN(new_n805));
  MUX2_X1   g380(.A(new_n796), .B(new_n805), .S(KEYINPUT28), .Z(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(G2067), .ZN(new_n807));
  NAND2_X1  g382(.A1(G168), .A2(G16), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G16), .B2(G21), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT94), .B(G1966), .Z(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n806), .A2(G2067), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n807), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n754), .A2(new_n769), .A3(new_n795), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n766), .A2(new_n768), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n747), .A2(new_n744), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n787), .A2(G2084), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OR3_X1    g395(.A1(new_n816), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n817), .B1(new_n816), .B2(new_n820), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n815), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n727), .A2(new_n731), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n809), .A2(new_n811), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n629), .A2(new_n680), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n825), .A2(KEYINPUT96), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n727), .A2(new_n827), .A3(new_n731), .A4(new_n823), .ZN(new_n830));
  INV_X1    g405(.A(new_n826), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n832), .ZN(G311));
  OR2_X1    g408(.A1(new_n830), .A2(new_n831), .ZN(G150));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n524), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT98), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(new_n514), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT99), .B(G55), .Z(new_n841));
  OAI22_X1  g416(.A1(new_n517), .A2(new_n840), .B1(new_n519), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n604), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT39), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n843), .B(new_n546), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n846), .B1(new_n852), .B2(G860), .ZN(G145));
  NAND2_X1  g428(.A1(new_n480), .A2(G142), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n487), .A2(G130), .ZN(new_n857));
  NOR2_X1   g432(.A1(G106), .A2(G2105), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(new_n483), .B2(G118), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n856), .B(new_n857), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n619), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n803), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n763), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n763), .A2(new_n863), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n780), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n764), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(new_n780), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n862), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(G160), .B(new_n629), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G162), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT100), .B1(new_n501), .B2(new_n504), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n873));
  INV_X1    g448(.A(new_n500), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n472), .B2(G126), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n873), .B(new_n503), .C1(new_n875), .C2(new_n483), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n872), .A2(new_n876), .B1(new_n497), .B2(new_n496), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n685), .B(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n871), .B(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n869), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(G37), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n869), .A2(new_n879), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g463(.A(new_n603), .B(G299), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(KEYINPUT105), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n889), .B(KEYINPUT41), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n893), .B2(KEYINPUT105), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n851), .B(KEYINPUT104), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n614), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n890), .B2(new_n896), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT42), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n591), .B(G166), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n577), .B(G290), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n901), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n897), .B(new_n907), .C1(new_n890), .C2(new_n896), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n899), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n906), .B1(new_n899), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(G868), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(G868), .B2(new_n843), .ZN(G295));
  OAI21_X1  g487(.A(new_n911), .B1(G868), .B2(new_n843), .ZN(G331));
  XNOR2_X1  g488(.A(new_n851), .B(G171), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n914), .A2(G286), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(G286), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n893), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n890), .B1(new_n915), .B2(new_n916), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n906), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n917), .B(new_n892), .C1(new_n893), .C2(KEYINPUT105), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n905), .A3(new_n919), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n923), .A3(new_n881), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n881), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n905), .B1(new_n922), .B2(new_n919), .ZN(new_n929));
  OR3_X1    g504(.A1(new_n928), .A2(KEYINPUT43), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n927), .A2(new_n930), .A3(KEYINPUT44), .A4(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n928), .B2(new_n929), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n921), .A2(new_n923), .A3(new_n934), .A4(new_n881), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n932), .A2(new_n938), .ZN(G397));
  NAND2_X1  g514(.A1(new_n872), .A2(new_n876), .ZN(new_n940));
  AOI21_X1  g515(.A(G1384), .B1(new_n940), .B2(new_n498), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT110), .B1(new_n941), .B2(KEYINPUT45), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  NOR4_X1   g519(.A1(new_n877), .A2(new_n943), .A3(new_n944), .A4(G1384), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n476), .A2(G40), .A3(new_n478), .ZN(new_n947));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n506), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n947), .B1(new_n949), .B2(new_n944), .ZN(new_n950));
  AOI21_X1  g525(.A(G1971), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n947), .ZN(new_n952));
  XOR2_X1   g527(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n952), .B1(new_n941), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n949), .A2(KEYINPUT50), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n955), .A2(G2090), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(G8), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G303), .A2(G8), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n959), .B(KEYINPUT55), .Z(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT112), .B(G1976), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(new_n579), .B2(new_n580), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n941), .A2(new_n952), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(G8), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n577), .A2(new_n967), .ZN(new_n968));
  NOR4_X1   g543(.A1(new_n964), .A2(KEYINPUT52), .A3(new_n966), .A4(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1981), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n589), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n545), .A2(G86), .ZN(new_n972));
  OAI21_X1  g547(.A(G1981), .B1(new_n588), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT49), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(KEYINPUT49), .A3(new_n973), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n976), .A2(G8), .A3(new_n965), .A4(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT52), .B1(new_n968), .B2(new_n966), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n969), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n947), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n982));
  INV_X1    g557(.A(new_n941), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(new_n953), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(G2090), .ZN(new_n985));
  OAI211_X1 g560(.A(G8), .B(new_n960), .C1(new_n951), .C2(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n962), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n946), .A2(new_n791), .A3(new_n950), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n989), .A2(new_n990), .B1(new_n744), .B2(new_n984), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n944), .B1(new_n877), .B2(G1384), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n992), .A2(new_n993), .A3(new_n952), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n992), .B2(new_n952), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n949), .A2(new_n944), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(KEYINPUT53), .A3(new_n791), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n991), .A2(new_n998), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n988), .A2(G301), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n997), .B2(new_n810), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n984), .A2(G2084), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n992), .A2(new_n952), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT114), .ZN(new_n1005));
  INV_X1    g580(.A(new_n996), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n992), .A2(new_n993), .A3(new_n952), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(KEYINPUT115), .A3(new_n811), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1002), .A2(new_n1003), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G286), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT51), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1002), .A2(G168), .A3(new_n1003), .A4(new_n1009), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(G8), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n1013), .B2(G8), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT62), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1010), .B2(G286), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(new_n1014), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT62), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n1018), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1000), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT126), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1018), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT125), .B(G2078), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n992), .A2(KEYINPUT53), .A3(new_n1029), .ZN(new_n1030));
  XOR2_X1   g605(.A(new_n947), .B(KEYINPUT124), .Z(new_n1031));
  NAND3_X1  g606(.A1(new_n946), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(G301), .B(KEYINPUT54), .Z(new_n1033));
  NAND3_X1  g608(.A1(new_n991), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n987), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n999), .A2(new_n1033), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1028), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n561), .A2(KEYINPUT57), .A3(new_n566), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT118), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n561), .A2(new_n566), .A3(new_n1040), .A4(KEYINPUT57), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  OR3_X1    g617(.A1(new_n557), .A2(KEYINPUT117), .A3(new_n560), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT117), .B1(new_n557), .B2(new_n560), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n566), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT56), .B(G2072), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n950), .B(new_n1049), .C1(new_n942), .C2(new_n945), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n742), .B1(new_n955), .B2(new_n956), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(new_n1051), .A3(new_n1050), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(KEYINPUT61), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT121), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1053), .A2(new_n1055), .A3(new_n1058), .A4(KEYINPUT61), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT61), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT58), .B(G1341), .Z(new_n1062));
  NAND2_X1  g637(.A1(new_n965), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT120), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n965), .A2(new_n1065), .A3(new_n1062), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT119), .B(G1996), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n950), .B(new_n1068), .C1(new_n942), .C2(new_n945), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n546), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT59), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n546), .C1(new_n1067), .C2(new_n1070), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1061), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1060), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n1060), .B2(new_n1075), .ZN(new_n1078));
  INV_X1    g653(.A(new_n965), .ZN(new_n1079));
  INV_X1    g654(.A(G2067), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n984), .A2(new_n734), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT60), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(new_n603), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1081), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1077), .A2(new_n1078), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1055), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n604), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(new_n1053), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1037), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n978), .A2(new_n581), .A3(new_n967), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n971), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(new_n966), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n986), .A2(new_n980), .A3(new_n969), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n1098));
  AND2_X1   g673(.A1(G168), .A2(G8), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1010), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1098), .B1(new_n1010), .B2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n987), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n981), .A2(new_n986), .ZN(new_n1105));
  OAI21_X1  g680(.A(G8), .B1(new_n951), .B2(new_n985), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1103), .B1(new_n1106), .B2(new_n961), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1105), .B(new_n1107), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n1096), .B(new_n1097), .C1(new_n1104), .C2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(KEYINPUT126), .B(new_n1000), .C1(new_n1020), .C2(new_n1024), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1027), .A2(new_n1091), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n992), .A2(new_n947), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1113), .A2(G1986), .A3(G290), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n697), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1114), .B1(G290), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT109), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n803), .B(new_n1080), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n763), .A2(G1996), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1118), .B(new_n1119), .C1(new_n867), .C2(G1996), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n690), .B2(new_n686), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n690), .B2(new_n686), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1122), .B2(new_n1112), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1111), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n686), .A2(new_n690), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1120), .A2(new_n1125), .B1(G2067), .B2(new_n803), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1126), .A2(new_n1112), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1113), .A2(G1996), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT127), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT46), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n1128), .B(new_n1130), .Z(new_n1131));
  INV_X1    g706(.A(new_n1118), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1112), .B1(new_n1132), .B2(new_n763), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1129), .B2(KEYINPUT46), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT47), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1122), .A2(new_n1112), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n1114), .B(KEYINPUT48), .Z(new_n1138));
  AOI211_X1 g713(.A(new_n1127), .B(new_n1136), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1124), .A2(new_n1139), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g715(.A(new_n462), .B1(new_n933), .B2(new_n935), .ZN(new_n1142));
  AOI211_X1 g716(.A(G401), .B(G227), .C1(new_n885), .C2(new_n886), .ZN(new_n1143));
  AND3_X1   g717(.A1(new_n1142), .A2(new_n1143), .A3(new_n678), .ZN(G308));
  NAND3_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(new_n678), .ZN(G225));
endmodule


