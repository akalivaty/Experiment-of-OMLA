//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n982, new_n983, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1039, new_n1040;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n204), .A2(G169gat), .A3(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n203), .A2(KEYINPUT66), .A3(new_n207), .A4(new_n205), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n210), .A2(new_n219), .A3(KEYINPUT25), .A4(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n212), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n225), .A3(new_n214), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n218), .A2(new_n215), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n226), .A2(new_n206), .A3(new_n203), .A4(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n218), .A2(KEYINPUT26), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT26), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n206), .B1(new_n202), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n223), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT27), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT67), .B1(new_n237), .B2(G183gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239));
  INV_X1    g038(.A(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT27), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(new_n237), .A3(G183gat), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(G183gat), .ZN(new_n245));
  AOI21_X1  g044(.A(G190gat), .B1(new_n245), .B2(KEYINPUT68), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT28), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT28), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(G190gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n240), .A2(KEYINPUT27), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT27), .B(G183gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(KEYINPUT69), .A3(new_n249), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n236), .B1(new_n247), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n231), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(G113gat), .B(G120gat), .Z(new_n259));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n260));
  XNOR2_X1  g059(.A(G127gat), .B(G134gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n259), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(G127gat), .B(G134gat), .Z(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n260), .ZN(new_n265));
  XNOR2_X1  g064(.A(G113gat), .B(G120gat), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n264), .B(new_n265), .C1(new_n266), .C2(KEYINPUT1), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n268), .A2(KEYINPUT71), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(KEYINPUT71), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n258), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n231), .A2(new_n257), .A3(KEYINPUT71), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT34), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n276), .B1(new_n274), .B2(KEYINPUT73), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n273), .B(new_n274), .C1(KEYINPUT73), .C2(new_n276), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G15gat), .B(G43gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G71gat), .B(G99gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n274), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n271), .A2(new_n285), .A3(new_n272), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n284), .B1(new_n286), .B2(KEYINPUT32), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT33), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n286), .A2(KEYINPUT72), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT72), .B1(new_n286), .B2(new_n288), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n287), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n286), .B(KEYINPUT32), .C1(new_n288), .C2(new_n284), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n281), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI211_X1 g094(.A(KEYINPUT74), .B(new_n280), .C1(new_n291), .C2(new_n292), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT36), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n293), .A2(new_n280), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n281), .B1(new_n292), .B2(new_n291), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT36), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT37), .ZN(new_n304));
  NAND2_X1  g103(.A1(G226gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n306), .B1(new_n258), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n305), .B1(new_n231), .B2(new_n257), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(G211gat), .A2(G218gat), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n311), .A2(KEYINPUT22), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(G211gat), .A2(G218gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n312), .B(new_n313), .C1(new_n311), .C2(new_n315), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n304), .B1(new_n310), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT69), .B1(new_n254), .B2(new_n249), .ZN(new_n322));
  AND4_X1   g121(.A1(KEYINPUT69), .A2(new_n249), .A3(new_n245), .A4(new_n250), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n245), .A2(KEYINPUT68), .ZN(new_n325));
  INV_X1    g124(.A(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n248), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n330), .A2(new_n236), .B1(new_n221), .B2(new_n230), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n305), .B1(new_n331), .B2(KEYINPUT29), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n220), .A2(new_n227), .A3(new_n226), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT25), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n208), .B2(new_n209), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n333), .A2(new_n335), .B1(new_n228), .B2(new_n229), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n235), .B1(new_n324), .B2(new_n329), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n306), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT75), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n308), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n321), .B1(new_n342), .B2(new_n320), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT88), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT38), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(G64gat), .B(G92gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(new_n231), .B2(new_n257), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n338), .B(new_n319), .C1(new_n349), .C2(new_n306), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n332), .A2(KEYINPUT76), .A3(new_n319), .A4(new_n338), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n320), .B1(new_n339), .B2(new_n341), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n304), .A3(new_n356), .ZN(new_n357));
  OAI211_X1 g156(.A(KEYINPUT88), .B(new_n321), .C1(new_n342), .C2(new_n320), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n345), .A2(new_n348), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  INV_X1    g159(.A(G148gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G141gat), .ZN(new_n362));
  INV_X1    g161(.A(G141gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G148gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT78), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT2), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G155gat), .ZN(new_n372));
  INV_X1    g171(.A(G162gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n371), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n366), .A2(new_n372), .A3(new_n373), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n380), .A2(new_n375), .B1(new_n362), .B2(new_n364), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n376), .B1(new_n365), .B2(new_n370), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT79), .B1(new_n384), .B2(new_n381), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n360), .B1(new_n386), .B2(new_n268), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n378), .A2(new_n388), .A3(new_n382), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT3), .B1(new_n384), .B2(new_n381), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n390), .A3(new_n268), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n263), .A2(new_n267), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n384), .A2(new_n381), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(KEYINPUT4), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(KEYINPUT5), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n387), .A2(new_n391), .A3(new_n394), .A4(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n394), .A2(new_n391), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n401), .A2(KEYINPUT80), .A3(new_n387), .A4(new_n397), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n391), .A2(KEYINPUT4), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n392), .A2(new_n393), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n386), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n407), .A3(new_n395), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n268), .B1(new_n381), .B2(new_n384), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n411), .B2(new_n396), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n400), .A2(new_n402), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414));
  INV_X1    g213(.A(G85gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT0), .B(G57gat), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n416), .B(new_n417), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT6), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n402), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n408), .A2(new_n412), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n418), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n418), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n340), .B1(new_n308), .B2(new_n309), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n332), .A2(KEYINPUT75), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n319), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT37), .B1(new_n430), .B2(new_n354), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n357), .A2(new_n431), .A3(new_n348), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT38), .ZN(new_n433));
  INV_X1    g232(.A(new_n348), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n355), .A2(new_n356), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT77), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n430), .A2(new_n354), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(KEYINPUT77), .A3(new_n434), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n359), .A2(new_n427), .A3(new_n433), .A4(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT39), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n404), .A2(new_n410), .A3(new_n395), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(KEYINPUT87), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(KEYINPUT87), .B2(new_n443), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n395), .B1(new_n401), .B2(new_n387), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT86), .B(KEYINPUT39), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n418), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n447), .A2(KEYINPUT40), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n424), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT40), .B1(new_n447), .B2(new_n449), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT30), .B1(new_n437), .B2(new_n439), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n438), .A2(KEYINPUT30), .A3(new_n434), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n348), .B1(new_n430), .B2(new_n354), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n453), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G78gat), .B(G106gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT83), .B(G50gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT31), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G22gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n314), .A2(KEYINPUT84), .A3(new_n316), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n307), .B(new_n466), .C1(new_n319), .C2(KEYINPUT84), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n406), .B1(new_n467), .B2(new_n388), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n319), .B1(new_n307), .B2(new_n389), .ZN(new_n469));
  INV_X1    g268(.A(G228gat), .ZN(new_n470));
  INV_X1    g269(.A(G233gat), .ZN(new_n471));
  OAI22_X1  g270(.A1(new_n468), .A2(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n470), .A2(new_n471), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT29), .B1(new_n393), .B2(new_n388), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT3), .B1(new_n319), .B2(new_n307), .ZN(new_n475));
  OAI221_X1 g274(.A(new_n473), .B1(new_n474), .B2(new_n319), .C1(new_n475), .C2(new_n393), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n465), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n464), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n467), .A2(new_n388), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n469), .B1(new_n480), .B2(new_n386), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n476), .B1(new_n481), .B2(new_n473), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G22gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n472), .A2(new_n465), .A3(new_n476), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n483), .A2(new_n478), .A3(new_n484), .A4(new_n464), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n459), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT30), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT77), .B1(new_n438), .B2(new_n434), .ZN(new_n492));
  NOR4_X1   g291(.A1(new_n430), .A2(new_n354), .A3(new_n436), .A4(new_n348), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n455), .A2(new_n456), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n420), .A2(new_n424), .A3(KEYINPUT81), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT81), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n423), .B(new_n418), .C1(new_n497), .C2(KEYINPUT6), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT82), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT82), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n494), .A2(new_n495), .A3(new_n502), .A4(new_n499), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n488), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n303), .B1(new_n490), .B2(new_n504), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n488), .A2(new_n299), .A3(new_n300), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n454), .A2(new_n457), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n427), .A2(KEYINPUT35), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n295), .ZN(new_n510));
  INV_X1    g309(.A(new_n296), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n488), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n501), .A2(new_n503), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n509), .B1(new_n513), .B2(KEYINPUT35), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G50gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G43gat), .ZN(new_n517));
  INV_X1    g316(.A(G43gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G50gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n519), .A3(KEYINPUT15), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(G29gat), .A2(G36gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(KEYINPUT14), .A3(new_n525), .ZN(new_n526));
  OR3_X1    g325(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT14), .ZN(new_n527));
  NAND2_X1  g326(.A1(G29gat), .A2(G36gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n518), .A2(KEYINPUT90), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G43gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n532), .A3(new_n516), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT91), .B1(new_n516), .B2(G43gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT15), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n530), .A2(new_n532), .A3(new_n538), .A4(new_n516), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n529), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n536), .A2(KEYINPUT92), .A3(new_n537), .A4(new_n539), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n521), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n529), .A2(new_n520), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT17), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G8gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n548));
  INV_X1    g347(.A(G15gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n465), .ZN(new_n550));
  NAND2_X1  g349(.A1(G15gat), .A2(G22gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(G1gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n550), .B2(new_n551), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n554), .A2(KEYINPUT16), .B1(new_n556), .B2(G1gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(G1gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OAI221_X1 g358(.A(new_n547), .B1(new_n548), .B2(new_n553), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n557), .A2(new_n559), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n547), .B1(new_n553), .B2(new_n548), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n539), .A2(new_n537), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT90), .B(G43gat), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n534), .B1(new_n566), .B2(new_n516), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n541), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n529), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n543), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n520), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572));
  INV_X1    g371(.A(new_n545), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n546), .A2(new_n564), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n564), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n545), .B1(new_n570), .B2(new_n520), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n575), .A2(KEYINPUT18), .A3(new_n576), .A4(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n576), .B(KEYINPUT13), .Z(new_n581));
  NOR2_X1   g380(.A1(new_n577), .A2(new_n578), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n571), .A2(new_n573), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(new_n564), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n581), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n564), .B1(new_n578), .B2(new_n572), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n544), .A2(KEYINPUT17), .A3(new_n545), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n579), .B(new_n576), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT18), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592));
  INV_X1    g391(.A(G197gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT11), .B(G169gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT12), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n586), .B(new_n591), .C1(KEYINPUT95), .C2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n591), .A2(new_n585), .A3(new_n580), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n580), .A2(KEYINPUT95), .A3(new_n585), .ZN(new_n600));
  INV_X1    g399(.A(new_n597), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n598), .A2(KEYINPUT96), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT96), .B1(new_n598), .B2(new_n602), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G64gat), .ZN(new_n607));
  INV_X1    g406(.A(G57gat), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n607), .B1(new_n608), .B2(KEYINPUT98), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT9), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n610), .A2(G71gat), .A3(G78gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n609), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n616), .A3(G57gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n608), .A2(KEYINPUT97), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n607), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n607), .A2(G57gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n608), .A2(G64gat), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n610), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G71gat), .B(G78gat), .ZN(new_n623));
  OAI22_X1  g422(.A1(new_n614), .A2(new_n619), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n577), .B1(KEYINPUT21), .B2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT99), .B(KEYINPUT19), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT20), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n628), .B(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n625), .A2(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n240), .ZN(new_n634));
  INV_X1    g433(.A(G211gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n632), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n631), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G232gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT100), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(KEYINPUT41), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(KEYINPUT41), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G85gat), .A2(G92gat), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT7), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G99gat), .B(G106gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(G99gat), .A2(G106gat), .ZN(new_n651));
  INV_X1    g450(.A(G92gat), .ZN(new_n652));
  AOI22_X1  g451(.A1(KEYINPUT8), .A2(new_n651), .B1(new_n415), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n649), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(KEYINPUT8), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n415), .A2(new_n652), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n655), .A2(new_n647), .A3(new_n656), .A4(new_n648), .ZN(new_n657));
  INV_X1    g456(.A(new_n650), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n654), .A2(new_n659), .A3(KEYINPUT101), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI211_X1 g463(.A(KEYINPUT102), .B(new_n644), .C1(new_n578), .C2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n571), .A2(new_n573), .A3(new_n664), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n667), .B2(new_n643), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n663), .B(new_n662), .C1(new_n578), .C2(new_n572), .ZN(new_n670));
  XOR2_X1   g469(.A(G190gat), .B(G218gat), .Z(new_n671));
  OAI22_X1  g470(.A1(new_n670), .A2(new_n588), .B1(KEYINPUT103), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n642), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n667), .A2(new_n643), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n667), .A2(new_n666), .A3(new_n643), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n664), .B1(new_n583), .B2(KEYINPUT17), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679));
  INV_X1    g478(.A(new_n671), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n678), .A2(new_n574), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n642), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n677), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(G134gat), .B(G162gat), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n673), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n673), .B2(new_n683), .ZN(new_n687));
  OAI22_X1  g486(.A1(new_n686), .A2(new_n687), .B1(new_n679), .B2(new_n680), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n683), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n684), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n680), .A2(new_n679), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n673), .A2(new_n683), .A3(new_n685), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n649), .B2(new_n653), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n624), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n660), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n660), .B(new_n695), .C1(new_n624), .C2(new_n697), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n625), .A2(KEYINPUT104), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(G230gat), .A2(G233gat), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT10), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n700), .A2(new_n708), .A3(new_n701), .A4(new_n702), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n664), .A2(KEYINPUT10), .A3(new_n625), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n704), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(G120gat), .B(G148gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(G176gat), .B(G204gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n713), .A2(new_n716), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n638), .A2(new_n694), .A3(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n515), .A2(new_n606), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n499), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G1gat), .ZN(G1324gat));
  INV_X1    g525(.A(new_n507), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT16), .B(G8gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n728), .A2(G8gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT106), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1325gat));
  NOR2_X1   g534(.A1(new_n299), .A2(new_n300), .ZN(new_n736));
  AOI21_X1  g535(.A(G15gat), .B1(new_n723), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n301), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT36), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT107), .B1(new_n298), .B2(new_n301), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n549), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n737), .B1(new_n723), .B2(new_n744), .ZN(G1326gat));
  NAND2_X1  g544(.A1(new_n723), .A2(new_n488), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G22gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n723), .A2(new_n465), .A3(new_n488), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n749), .B(new_n751), .ZN(G1327gat));
  AND2_X1   g551(.A1(new_n688), .A2(new_n693), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n631), .B(new_n637), .Z(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n721), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n606), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n753), .B(new_n756), .C1(new_n505), .C2(new_n514), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n757), .A2(G29gat), .A3(new_n499), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(KEYINPUT45), .Z(new_n759));
  AOI22_X1  g558(.A1(new_n490), .A2(new_n504), .B1(new_n741), .B2(new_n742), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n753), .B1(new_n760), .B2(new_n514), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g562(.A(KEYINPUT44), .B(new_n753), .C1(new_n505), .C2(new_n514), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n598), .A2(new_n602), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n755), .A2(new_n766), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n763), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n724), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G29gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n759), .A2(new_n770), .ZN(G1328gat));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n727), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G36gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n757), .A2(G36gat), .A3(new_n507), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT46), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1329gat));
  INV_X1    g575(.A(new_n743), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n763), .A2(new_n777), .A3(new_n764), .A4(new_n767), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n566), .ZN(new_n779));
  INV_X1    g578(.A(new_n736), .ZN(new_n780));
  OR3_X1    g579(.A1(new_n757), .A2(new_n780), .A3(new_n566), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1330gat));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n763), .A2(new_n488), .A3(new_n764), .A4(new_n767), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(G50gat), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n757), .A2(G50gat), .A3(new_n489), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n786), .B2(G50gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT48), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  AOI221_X4 g590(.A(new_n788), .B1(new_n785), .B2(KEYINPUT48), .C1(new_n786), .C2(G50gat), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(G1331gat));
  NAND2_X1  g592(.A1(new_n490), .A2(new_n504), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n743), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n513), .A2(KEYINPUT35), .ZN(new_n796));
  INV_X1    g595(.A(new_n509), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NOR4_X1   g598(.A1(new_n754), .A2(new_n753), .A3(new_n765), .A4(new_n721), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n724), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n615), .A2(G57gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n618), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n803), .B(new_n805), .ZN(G1332gat));
  AOI21_X1  g605(.A(new_n507), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT110), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n809), .B(new_n810), .Z(G1333gat));
  INV_X1    g610(.A(G71gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n801), .B2(new_n780), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n777), .A2(G71gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n801), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n815), .B(new_n816), .ZN(G1334gat));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n488), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(G78gat), .ZN(G1335gat));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n638), .A2(new_n765), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n799), .A2(new_n820), .A3(new_n753), .A4(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n753), .B(new_n821), .C1(new_n760), .C2(new_n514), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT51), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n822), .A2(new_n824), .A3(new_n720), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n415), .A3(new_n724), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n821), .A2(new_n720), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(KEYINPUT112), .Z(new_n828));
  NAND3_X1  g627(.A1(new_n763), .A2(new_n764), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(G85gat), .B1(new_n829), .B2(new_n499), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n830), .ZN(G1336gat));
  OAI21_X1  g630(.A(G92gat), .B1(new_n829), .B2(new_n507), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n507), .A2(G92gat), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n822), .A2(new_n824), .A3(new_n720), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n832), .B(new_n834), .C1(new_n837), .C2(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1337gat));
  INV_X1    g640(.A(G99gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n842), .A3(new_n736), .ZN(new_n843));
  OAI21_X1  g642(.A(G99gat), .B1(new_n829), .B2(new_n743), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1338gat));
  INV_X1    g644(.A(G106gat), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n489), .A2(new_n846), .ZN(new_n847));
  AND4_X1   g646(.A1(new_n763), .A2(new_n764), .A3(new_n828), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n822), .A2(new_n824), .A3(new_n488), .A4(new_n720), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT53), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n846), .ZN(new_n853));
  INV_X1    g652(.A(new_n848), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(KEYINPUT114), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n857), .ZN(G1339gat));
  NAND3_X1  g657(.A1(new_n709), .A2(new_n705), .A3(new_n710), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n709), .A2(KEYINPUT115), .A3(new_n710), .A4(new_n705), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n861), .A2(new_n712), .A3(KEYINPUT54), .A4(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n716), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n705), .B1(new_n709), .B2(new_n710), .ZN(new_n865));
  XNOR2_X1  g664(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n863), .A2(KEYINPUT55), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT117), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n863), .A2(new_n873), .A3(KEYINPUT55), .A4(new_n867), .ZN(new_n874));
  AND4_X1   g673(.A1(KEYINPUT118), .A2(new_n872), .A3(new_n718), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n717), .B1(new_n871), .B2(KEYINPUT117), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT118), .B1(new_n876), .B2(new_n874), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n765), .B(new_n870), .C1(new_n875), .C2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n599), .A2(new_n601), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n576), .B1(new_n575), .B2(new_n579), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n582), .A2(new_n584), .A3(new_n581), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n879), .B1(new_n596), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n720), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n753), .B1(new_n878), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n870), .B1(new_n875), .B2(new_n877), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n688), .A2(new_n883), .A3(new_n693), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n754), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n754), .A2(new_n753), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n766), .A3(new_n721), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n506), .A2(new_n507), .A3(new_n724), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G113gat), .B1(new_n895), .B2(new_n606), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n510), .A2(new_n511), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n892), .A2(new_n724), .A3(new_n489), .A4(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n488), .B1(new_n889), .B2(new_n891), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n901), .A2(KEYINPUT119), .A3(new_n724), .A4(new_n897), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n507), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n766), .A2(G113gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n896), .B1(new_n904), .B2(new_n905), .ZN(G1340gat));
  OAI21_X1  g705(.A(G120gat), .B1(new_n895), .B2(new_n721), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n721), .A2(G120gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n904), .B2(new_n908), .ZN(G1341gat));
  INV_X1    g708(.A(G127gat), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n895), .A2(new_n910), .A3(new_n754), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n507), .B(new_n638), .C1(new_n900), .C2(new_n903), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n910), .ZN(G1342gat));
  INV_X1    g712(.A(G134gat), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n894), .B2(new_n753), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n727), .A2(new_n694), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n914), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n899), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n902), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n917), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n900), .B2(new_n903), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT120), .B1(new_n923), .B2(KEYINPUT56), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n919), .A2(new_n925), .A3(new_n920), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n921), .B1(new_n924), .B2(new_n926), .ZN(G1343gat));
  AOI21_X1  g726(.A(new_n489), .B1(new_n889), .B2(new_n891), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n724), .A3(new_n743), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n727), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n606), .A2(G141gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT58), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT96), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n765), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n872), .A2(new_n870), .A3(new_n718), .A4(new_n874), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n598), .A2(new_n602), .A3(KEYINPUT96), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n753), .B1(new_n938), .B2(new_n884), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n754), .B1(new_n939), .B2(new_n888), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n940), .A2(new_n891), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT57), .B1(new_n941), .B2(new_n489), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n777), .A2(new_n499), .A3(new_n727), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT57), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n944), .A2(new_n947), .A3(new_n606), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n932), .B1(new_n948), .B2(new_n363), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n942), .A2(new_n946), .A3(new_n765), .A4(new_n943), .ZN(new_n950));
  AOI22_X1  g749(.A1(new_n950), .A2(G141gat), .B1(new_n930), .B2(new_n931), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT58), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1344gat));
  NAND3_X1  g752(.A1(new_n930), .A2(new_n361), .A3(new_n720), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT59), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n722), .A2(new_n605), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n489), .B1(new_n940), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT121), .B1(new_n957), .B2(KEYINPUT57), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n722), .A2(new_n605), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n603), .A2(new_n604), .A3(new_n935), .ZN(new_n961));
  INV_X1    g760(.A(new_n884), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n694), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n877), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n876), .A2(KEYINPUT118), .A3(new_n874), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n966), .A2(new_n753), .A3(new_n870), .A4(new_n883), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n960), .B1(new_n968), .B2(new_n754), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n959), .B(new_n945), .C1(new_n969), .C2(new_n489), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n928), .A2(KEYINPUT57), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n958), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n972), .A2(new_n720), .A3(new_n943), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n955), .B1(new_n973), .B2(G148gat), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n955), .A2(G148gat), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n944), .A2(new_n947), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n720), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n954), .B1(new_n974), .B2(new_n977), .ZN(G1345gat));
  AOI21_X1  g777(.A(G155gat), .B1(new_n930), .B2(new_n638), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n754), .A2(new_n372), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n976), .B2(new_n980), .ZN(G1346gat));
  NOR3_X1   g780(.A1(new_n944), .A2(new_n694), .A3(new_n947), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n916), .A2(new_n373), .ZN(new_n983));
  OAI22_X1  g782(.A1(new_n982), .A2(new_n373), .B1(new_n929), .B2(new_n983), .ZN(G1347gat));
  NOR2_X1   g783(.A1(new_n507), .A2(new_n724), .ZN(new_n985));
  AND4_X1   g784(.A1(new_n489), .A2(new_n892), .A3(new_n897), .A4(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n986), .A2(new_n216), .A3(new_n765), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n985), .A2(new_n736), .ZN(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n901), .A2(KEYINPUT122), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT122), .B1(new_n901), .B2(new_n989), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n990), .A2(new_n991), .A3(new_n606), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n987), .B1(new_n992), .B2(new_n216), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(KEYINPUT123), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT123), .ZN(new_n995));
  OAI211_X1 g794(.A(new_n987), .B(new_n995), .C1(new_n992), .C2(new_n216), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n996), .ZN(G1348gat));
  AOI21_X1  g796(.A(G176gat), .B1(new_n986), .B2(new_n720), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n990), .A2(new_n991), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n721), .A2(new_n217), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(G1349gat));
  NAND3_X1  g800(.A1(new_n892), .A2(new_n489), .A3(new_n989), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT122), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n901), .A2(KEYINPUT122), .A3(new_n989), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1004), .A2(new_n638), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(G183gat), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n986), .A2(new_n254), .A3(new_n638), .ZN(new_n1008));
  XNOR2_X1  g807(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1009), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n1010), .A2(new_n1011), .ZN(G1350gat));
  NAND3_X1  g811(.A1(new_n986), .A2(new_n326), .A3(new_n753), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1004), .A2(new_n753), .A3(new_n1005), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT61), .ZN(new_n1015));
  AND3_X1   g814(.A1(new_n1014), .A2(new_n1015), .A3(G190gat), .ZN(new_n1016));
  AOI21_X1  g815(.A(new_n1015), .B1(new_n1014), .B2(G190gat), .ZN(new_n1017));
  OAI21_X1  g816(.A(new_n1013), .B1(new_n1016), .B2(new_n1017), .ZN(G1351gat));
  AND2_X1   g817(.A1(new_n743), .A2(new_n985), .ZN(new_n1019));
  AND2_X1   g818(.A1(new_n972), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1020), .A2(new_n605), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1021), .A2(G197gat), .ZN(new_n1022));
  AND2_X1   g821(.A1(new_n928), .A2(new_n1019), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1023), .A2(new_n593), .A3(new_n765), .ZN(new_n1024));
  XOR2_X1   g823(.A(new_n1024), .B(KEYINPUT125), .Z(new_n1025));
  NAND2_X1  g824(.A1(new_n1022), .A2(new_n1025), .ZN(G1352gat));
  XOR2_X1   g825(.A(KEYINPUT126), .B(G204gat), .Z(new_n1027));
  NOR2_X1   g826(.A1(new_n721), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g828(.A(new_n1029), .B(KEYINPUT62), .Z(new_n1030));
  NAND3_X1  g829(.A1(new_n972), .A2(new_n720), .A3(new_n1019), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n1031), .A2(new_n1027), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1030), .A2(new_n1032), .ZN(G1353gat));
  NAND3_X1  g832(.A1(new_n1023), .A2(new_n635), .A3(new_n638), .ZN(new_n1034));
  NAND3_X1  g833(.A1(new_n972), .A2(new_n638), .A3(new_n1019), .ZN(new_n1035));
  AND3_X1   g834(.A1(new_n1035), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1036));
  AOI21_X1  g835(.A(KEYINPUT63), .B1(new_n1035), .B2(G211gat), .ZN(new_n1037));
  OAI21_X1  g836(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(G1354gat));
  AOI21_X1  g837(.A(G218gat), .B1(new_n1023), .B2(new_n753), .ZN(new_n1039));
  AND2_X1   g838(.A1(new_n753), .A2(G218gat), .ZN(new_n1040));
  AOI21_X1  g839(.A(new_n1039), .B1(new_n1020), .B2(new_n1040), .ZN(G1355gat));
endmodule


