//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT36), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G190gat), .Z(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT27), .B(G183gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT28), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n213), .B1(new_n216), .B2(KEYINPUT26), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(KEYINPUT26), .B2(new_n216), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n208), .A2(KEYINPUT28), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n209), .A2(new_n210), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n213), .B1(KEYINPUT23), .B2(new_n214), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT25), .B1(new_n214), .B2(KEYINPUT23), .ZN(new_n224));
  OR3_X1    g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT24), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n206), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT65), .B(G190gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(G183gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(KEYINPUT66), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n229), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT67), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(new_n232), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(KEYINPUT66), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n229), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n225), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n211), .B2(new_n212), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n229), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(KEYINPUT25), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n220), .B1(new_n244), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G113gat), .ZN(new_n253));
  INV_X1    g052(.A(G120gat), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT1), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G127gat), .B(G134gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n257));
  OAI221_X1 g056(.A(new_n255), .B1(new_n253), .B2(new_n254), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n257), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n258), .B(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n252), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n220), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n242), .B1(new_n241), .B2(new_n229), .ZN(new_n265));
  INV_X1    g064(.A(new_n229), .ZN(new_n266));
  AOI211_X1 g065(.A(KEYINPUT67), .B(new_n266), .C1(new_n239), .C2(new_n240), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n251), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n263), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n258), .B(new_n259), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n262), .A2(new_n272), .A3(G227gat), .A4(G233gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT32), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT33), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G15gat), .B(G43gat), .Z(new_n277));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n279), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n273), .B(KEYINPUT32), .C1(new_n275), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n262), .A2(new_n272), .ZN(new_n283));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284));
  AND2_X1   g083(.A1(KEYINPUT70), .A2(KEYINPUT34), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n262), .A2(new_n272), .B1(G227gat), .B2(G233gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n280), .A2(new_n282), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n280), .B2(new_n282), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n204), .B(new_n205), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n280), .A2(new_n282), .ZN(new_n293));
  INV_X1    g092(.A(new_n289), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n282), .A3(new_n289), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n295), .A2(new_n202), .A3(new_n203), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT3), .ZN(new_n299));
  XOR2_X1   g098(.A(G197gat), .B(G204gat), .Z(new_n300));
  NAND2_X1  g099(.A1(G211gat), .A2(G218gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(KEYINPUT22), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(G211gat), .A2(G218gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n304), .B2(new_n306), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n299), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G141gat), .B(G148gat), .Z(new_n311));
  NOR2_X1   g110(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n312));
  AND2_X1   g111(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G155gat), .B(G162gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT75), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(G155gat), .B2(G162gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT77), .B(G162gat), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT2), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n311), .A3(new_n315), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n310), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n304), .B(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n319), .A2(new_n299), .A3(new_n323), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n308), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G228gat), .ZN(new_n330));
  INV_X1    g129(.A(G233gat), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n325), .A2(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT81), .ZN(new_n333));
  INV_X1    g132(.A(new_n327), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT82), .B1(new_n334), .B2(KEYINPUT29), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n299), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n334), .A2(KEYINPUT82), .A3(KEYINPUT29), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n324), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G78gat), .B(G106gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT31), .B(G50gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G22gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(KEYINPUT83), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n345), .B1(new_n347), .B2(new_n343), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n333), .A2(new_n340), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n349), .B1(new_n333), .B2(new_n340), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G226gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(new_n331), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(KEYINPUT29), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n270), .A2(new_n355), .ZN(new_n356));
  AOI211_X1 g155(.A(new_n263), .B(new_n354), .C1(new_n268), .C2(new_n269), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n334), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n354), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n220), .B(new_n359), .C1(new_n244), .C2(new_n251), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n360), .B(new_n327), .C1(new_n270), .C2(new_n355), .ZN(new_n361));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  NAND3_X1  g163(.A1(new_n358), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(KEYINPUT74), .B(KEYINPUT30), .Z(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n364), .ZN(new_n369));
  INV_X1    g168(.A(new_n361), .ZN(new_n370));
  INV_X1    g169(.A(new_n355), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n252), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n327), .B1(new_n372), .B2(new_n360), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n369), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n358), .A2(KEYINPUT30), .A3(new_n361), .A4(new_n364), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT73), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT73), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n368), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT4), .B1(new_n271), .B2(new_n324), .ZN(new_n381));
  INV_X1    g180(.A(new_n324), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n261), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(new_n271), .A3(new_n328), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT78), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n385), .A2(new_n391), .A3(new_n386), .A4(new_n388), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT5), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n261), .A2(new_n382), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n271), .A2(new_n324), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n386), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n390), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n394), .A2(new_n400), .A3(KEYINPUT4), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n388), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n381), .A2(new_n384), .A3(KEYINPUT79), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n403), .A2(new_n393), .A3(new_n386), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G1gat), .B(G29gat), .Z(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(KEYINPUT0), .ZN(new_n408));
  XNOR2_X1  g207(.A(G57gat), .B(G85gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT80), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n406), .A2(new_n411), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT80), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n399), .A2(new_n405), .A3(new_n415), .A4(new_n410), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n412), .A2(new_n413), .A3(new_n414), .A4(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n406), .A2(KEYINPUT6), .A3(new_n411), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n352), .B1(new_n380), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n298), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n410), .B(KEYINPUT84), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n386), .B1(new_n403), .B2(new_n404), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT39), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n396), .A2(new_n397), .ZN(new_n426));
  OR3_X1    g225(.A1(new_n426), .A2(KEYINPUT85), .A3(new_n424), .ZN(new_n427));
  INV_X1    g226(.A(new_n404), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n397), .B1(new_n428), .B2(new_n402), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT85), .B1(new_n426), .B2(new_n424), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT40), .B1(new_n432), .B2(KEYINPUT86), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n406), .A2(new_n422), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n367), .A2(new_n374), .A3(new_n375), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT86), .B1(new_n425), .B2(new_n431), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT40), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n433), .A2(new_n434), .A3(new_n435), .A4(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT37), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n374), .B1(new_n440), .B2(new_n364), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n358), .A2(new_n361), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT37), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n440), .B1(new_n358), .B2(new_n361), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT38), .B1(new_n446), .B2(KEYINPUT87), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n441), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n369), .B1(new_n442), .B2(KEYINPUT37), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT38), .B1(new_n449), .B2(new_n446), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n450), .A3(new_n365), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n412), .A2(new_n434), .A3(new_n414), .A4(new_n416), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n418), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n352), .B(new_n439), .C1(new_n451), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n380), .A2(new_n419), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n295), .A2(new_n352), .A3(new_n296), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT35), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT35), .B1(new_n452), .B2(new_n418), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n290), .A2(new_n291), .ZN(new_n459));
  INV_X1    g258(.A(new_n435), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n352), .A4(new_n460), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n421), .A2(new_n454), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n344), .A2(G15gat), .ZN(new_n463));
  INV_X1    g262(.A(G15gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G22gat), .ZN(new_n465));
  INV_X1    g264(.A(G1gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT16), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(G1gat), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(new_n469), .B2(G1gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(G8gat), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G8gat), .ZN(new_n474));
  OAI221_X1 g273(.A(new_n468), .B1(new_n471), .B2(new_n474), .C1(G1gat), .C2(new_n469), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(G43gat), .A2(G50gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(G43gat), .A2(G50gat), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT15), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR4_X1   g279(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT89), .A4(KEYINPUT15), .ZN(new_n481));
  INV_X1    g280(.A(G29gat), .ZN(new_n482));
  INV_X1    g281(.A(G36gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT14), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT14), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(G29gat), .B2(G36gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(G29gat), .A2(G36gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n480), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n480), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n492));
  OR3_X1    g291(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT15), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n489), .A2(new_n494), .A3(KEYINPUT17), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT17), .B1(new_n489), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n477), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n489), .A2(new_n494), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n476), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT18), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n497), .A2(KEYINPUT18), .A3(new_n498), .A4(new_n501), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n499), .A2(new_n475), .A3(new_n473), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n498), .B(KEYINPUT13), .Z(new_n508));
  AOI21_X1  g307(.A(KEYINPUT91), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT91), .ZN(new_n510));
  INV_X1    g309(.A(new_n508), .ZN(new_n511));
  AOI211_X1 g310(.A(new_n510), .B(new_n511), .C1(new_n501), .C2(new_n506), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n504), .B(new_n505), .C1(new_n509), .C2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G113gat), .B(G141gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(G197gat), .ZN(new_n515));
  XOR2_X1   g314(.A(KEYINPUT11), .B(G169gat), .Z(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n517), .B(KEYINPUT12), .Z(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n513), .A2(KEYINPUT88), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n513), .B2(KEYINPUT88), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G218gat), .ZN(new_n524));
  INV_X1    g323(.A(G190gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n530));
  INV_X1    g329(.A(G92gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT8), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n533), .A2(KEYINPUT100), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT100), .B1(new_n533), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n529), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT101), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G99gat), .ZN(new_n542));
  INV_X1    g341(.A(G106gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT101), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n534), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n538), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT100), .ZN(new_n549));
  AND2_X1   g348(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n550), .A2(new_n551), .A3(G92gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n535), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n533), .A2(KEYINPUT100), .A3(new_n535), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n547), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(new_n529), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n499), .B1(new_n548), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT41), .ZN(new_n560));
  INV_X1    g359(.A(G232gat), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n560), .A2(new_n561), .A3(new_n331), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT102), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n557), .B1(new_n556), .B2(new_n529), .ZN(new_n564));
  AOI211_X1 g363(.A(new_n528), .B(new_n547), .C1(new_n554), .C2(new_n555), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n500), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT102), .ZN(new_n567));
  INV_X1    g366(.A(new_n562), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n495), .A2(new_n496), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n548), .A2(new_n558), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n525), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  AOI211_X1 g374(.A(G190gat), .B(new_n573), .C1(new_n563), .C2(new_n569), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n524), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n559), .A2(KEYINPUT102), .A3(new_n562), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n567), .B1(new_n566), .B2(new_n568), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n574), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(G190gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n570), .A2(new_n525), .A3(new_n574), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(G218gat), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n577), .A2(new_n583), .A3(KEYINPUT97), .ZN(new_n584));
  XNOR2_X1  g383(.A(G134gat), .B(G162gat), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n560), .B1(new_n561), .B2(new_n331), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G57gat), .ZN(new_n592));
  INV_X1    g391(.A(G64gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G57gat), .A2(G64gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(KEYINPUT9), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT92), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT92), .B1(G71gat), .B2(G78gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT93), .B1(new_n597), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT93), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n607), .A3(new_n596), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n599), .A2(new_n600), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT94), .B1(new_n609), .B2(KEYINPUT9), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n599), .B(new_n600), .C1(KEYINPUT94), .C2(KEYINPUT9), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n602), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n605), .A2(new_n608), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n476), .B1(new_n614), .B2(KEYINPUT21), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n614), .A2(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(G127gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n618), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n617), .B(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(G127gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n616), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(new_n624), .A3(new_n616), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(new_n321), .ZN(new_n629));
  XNOR2_X1  g428(.A(G183gat), .B(G211gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n629), .B(new_n630), .Z(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  INV_X1    g432(.A(new_n627), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n625), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n577), .A2(new_n583), .A3(KEYINPUT97), .A4(new_n589), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n614), .B1(new_n564), .B2(new_n565), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n613), .A2(new_n610), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n597), .A2(new_n604), .A3(KEYINPUT93), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n607), .B1(new_n606), .B2(new_n596), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n548), .A2(new_n643), .A3(new_n558), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n614), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n638), .A2(new_n644), .ZN(new_n650));
  INV_X1    g449(.A(new_n648), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n649), .A2(new_n652), .A3(new_n656), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n591), .A2(new_n636), .A3(new_n637), .A4(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n462), .A2(new_n523), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n419), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT104), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT103), .B(G1gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(G1324gat));
  INV_X1    g467(.A(new_n663), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n669), .A2(new_n460), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n474), .B1(new_n663), .B2(new_n435), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT42), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(KEYINPUT42), .B2(new_n671), .ZN(G1325gat));
  AND2_X1   g473(.A1(new_n292), .A2(new_n297), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT105), .ZN(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n669), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n663), .A2(new_n464), .A3(new_n459), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1326gat));
  NOR3_X1   g478(.A1(new_n462), .A2(new_n352), .A3(new_n523), .ZN(new_n680));
  INV_X1    g479(.A(new_n662), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  AND2_X1   g483(.A1(new_n591), .A2(new_n637), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n636), .A2(new_n660), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n522), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n462), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n482), .A3(new_n664), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  INV_X1    g489(.A(new_n352), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n455), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n454), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n457), .A2(new_n461), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n591), .A2(new_n637), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n685), .B1(new_n693), .B2(new_n694), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n696), .A3(KEYINPUT44), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(new_n419), .A3(new_n687), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n690), .B1(new_n482), .B2(new_n704), .ZN(G1328gat));
  NOR4_X1   g504(.A1(new_n462), .A2(KEYINPUT106), .A3(new_n699), .A4(new_n685), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT44), .B1(new_n701), .B2(new_n696), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709));
  INV_X1    g508(.A(new_n687), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n435), .A4(new_n710), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n700), .A2(new_n435), .A3(new_n702), .A4(new_n710), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT107), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n713), .A3(G36gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n688), .A2(new_n483), .A3(new_n435), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT46), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n714), .A2(new_n716), .A3(KEYINPUT108), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1329gat));
  INV_X1    g520(.A(G43gat), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n688), .A2(new_n722), .A3(new_n459), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n703), .A2(new_n687), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n298), .B(KEYINPUT105), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n723), .B1(new_n726), .B2(G43gat), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n722), .B1(new_n724), .B2(new_n298), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n727), .A2(KEYINPUT47), .B1(new_n728), .B2(new_n730), .ZN(G1330gat));
  INV_X1    g530(.A(G50gat), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n680), .A2(new_n732), .A3(new_n697), .A4(new_n686), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n703), .A2(new_n352), .A3(new_n687), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(new_n732), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1331gat));
  NAND4_X1  g536(.A1(new_n685), .A2(new_n523), .A3(new_n636), .A4(new_n660), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n462), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n664), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g540(.A1(new_n462), .A2(new_n460), .A3(new_n738), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(G1333gat));
  AOI21_X1  g545(.A(new_n599), .B1(new_n739), .B2(new_n725), .ZN(new_n747));
  INV_X1    g546(.A(new_n459), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(G71gat), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n747), .B1(new_n739), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n739), .A2(new_n691), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n636), .A2(new_n522), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n660), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT109), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n700), .A2(new_n702), .A3(new_n756), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n757), .A2(new_n664), .B1(new_n530), .B2(new_n532), .ZN(new_n758));
  NAND2_X1  g557(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n695), .A2(new_n697), .A3(new_n754), .A4(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n754), .ZN(new_n764));
  AOI211_X1 g563(.A(new_n685), .B(new_n764), .C1(new_n693), .C2(new_n694), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n763), .B(new_n660), .C1(new_n765), .C2(new_n759), .ZN(new_n766));
  NOR4_X1   g565(.A1(new_n766), .A2(new_n419), .A3(new_n551), .A4(new_n550), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n758), .A2(new_n767), .ZN(G1336gat));
  NAND4_X1  g567(.A1(new_n700), .A2(new_n435), .A3(new_n702), .A4(new_n756), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G92gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT111), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n772), .A3(G92gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n695), .A2(new_n697), .A3(new_n754), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n760), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n460), .A2(G92gat), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n775), .A2(new_n660), .A3(new_n763), .A4(new_n776), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n771), .A2(new_n773), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n780), .A2(new_n781), .A3(new_n770), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n780), .B2(new_n770), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n778), .A2(new_n779), .B1(new_n782), .B2(new_n783), .ZN(G1337gat));
  OR2_X1    g583(.A1(new_n766), .A2(new_n748), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n676), .A2(new_n542), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n785), .A2(new_n542), .B1(new_n757), .B2(new_n786), .ZN(G1338gat));
  OAI21_X1  g586(.A(new_n543), .B1(new_n766), .B2(new_n352), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n352), .A2(new_n543), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n700), .A2(new_n702), .A3(new_n756), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n791), .A2(KEYINPUT113), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n775), .A2(new_n691), .A3(new_n660), .A4(new_n763), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n757), .A2(new_n789), .B1(new_n795), .B2(new_n543), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n796), .B2(KEYINPUT53), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT114), .B1(new_n791), .B2(new_n792), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  AOI211_X1 g598(.A(new_n799), .B(KEYINPUT53), .C1(new_n788), .C2(new_n790), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n793), .A2(new_n797), .B1(new_n798), .B2(new_n800), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n507), .A2(new_n508), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n498), .B1(new_n497), .B2(new_n501), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n517), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n660), .B(new_n804), .C1(new_n513), .C2(new_n518), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n647), .B2(new_n648), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n645), .A2(new_n646), .A3(new_n651), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n651), .B1(new_n645), .B2(new_n646), .ZN(new_n811));
  XOR2_X1   g610(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n812));
  AOI211_X1 g611(.A(KEYINPUT117), .B(new_n656), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n647), .A2(new_n648), .A3(new_n812), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n657), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n810), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n522), .A2(new_n817), .A3(new_n659), .ZN(new_n818));
  INV_X1    g617(.A(new_n812), .ZN(new_n819));
  AOI211_X1 g618(.A(new_n651), .B(new_n819), .C1(new_n645), .C2(new_n646), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT117), .B1(new_n820), .B2(new_n656), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n815), .A2(new_n814), .A3(new_n657), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n809), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT55), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n805), .B1(new_n818), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n685), .ZN(new_n827));
  INV_X1    g626(.A(new_n825), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n804), .B1(new_n513), .B2(new_n518), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n649), .A2(new_n652), .A3(new_n656), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n697), .A2(new_n828), .A3(new_n817), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n636), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n681), .A2(new_n835), .A3(new_n523), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT115), .B1(new_n662), .B2(new_n522), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n833), .A2(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n419), .A2(new_n435), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n838), .A2(new_n456), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n523), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n833), .A2(new_n834), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n836), .A2(new_n837), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n664), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n847), .A2(new_n435), .A3(new_n456), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n522), .A2(new_n253), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT118), .Z(new_n851));
  OAI21_X1  g650(.A(new_n843), .B1(new_n849), .B2(new_n851), .ZN(G1340gat));
  AOI21_X1  g651(.A(G120gat), .B1(new_n848), .B2(new_n660), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n661), .A2(new_n254), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n841), .B2(new_n854), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n848), .A2(new_n623), .A3(new_n636), .ZN(new_n856));
  OAI21_X1  g655(.A(G127gat), .B1(new_n842), .B2(new_n834), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1342gat));
  OR3_X1    g657(.A1(new_n849), .A2(G134gat), .A3(new_n685), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n859), .A2(KEYINPUT56), .ZN(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n842), .B2(new_n685), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(KEYINPUT56), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n840), .A2(new_n298), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n691), .A2(KEYINPUT57), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n821), .A2(new_n822), .B1(new_n809), .B2(new_n808), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n831), .B(new_n817), .C1(new_n868), .C2(KEYINPUT55), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n637), .B2(new_n591), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n827), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n826), .A2(new_n685), .A3(KEYINPUT120), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n636), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n845), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n865), .B(new_n867), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n838), .B2(new_n352), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n520), .A2(new_n521), .A3(new_n830), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n880), .B(new_n817), .C1(KEYINPUT55), .C2(new_n868), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n697), .B1(new_n805), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n832), .B1(new_n882), .B2(KEYINPUT120), .ZN(new_n883));
  INV_X1    g682(.A(new_n873), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n834), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n845), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n865), .B1(new_n886), .B2(new_n867), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n522), .B(new_n864), .C1(new_n879), .C2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(G141gat), .ZN(new_n889));
  NOR4_X1   g688(.A1(new_n847), .A2(new_n725), .A3(new_n352), .A4(new_n435), .ZN(new_n890));
  INV_X1    g689(.A(G141gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n522), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT122), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT58), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n891), .B1(new_n888), .B2(KEYINPUT123), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n827), .A2(new_n871), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n832), .A3(new_n873), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n901), .A2(new_n834), .B1(new_n837), .B2(new_n836), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT121), .B1(new_n902), .B2(new_n866), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n878), .A3(new_n876), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n904), .A2(new_n905), .A3(new_n522), .A4(new_n864), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT124), .B(new_n898), .C1(new_n899), .C2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(G141gat), .A3(new_n906), .ZN(new_n910));
  INV_X1    g709(.A(new_n898), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n896), .B1(new_n907), .B2(new_n912), .ZN(G1344gat));
  INV_X1    g712(.A(G148gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n890), .A2(new_n914), .A3(new_n660), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n904), .A2(new_n864), .ZN(new_n916));
  AOI211_X1 g715(.A(KEYINPUT59), .B(new_n914), .C1(new_n916), .C2(new_n660), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n662), .A2(new_n522), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n844), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n923), .B2(new_n691), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n838), .A2(new_n352), .A3(new_n877), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n660), .A3(new_n864), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n918), .B1(new_n927), .B2(G148gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n915), .B1(new_n917), .B2(new_n928), .ZN(G1345gat));
  NAND3_X1  g728(.A1(new_n890), .A2(new_n321), .A3(new_n636), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n916), .A2(new_n636), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n930), .B1(new_n932), .B2(new_n321), .ZN(G1346gat));
  NOR2_X1   g732(.A1(new_n685), .A2(new_n320), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n890), .A2(new_n697), .ZN(new_n935));
  AOI22_X1  g734(.A1(new_n916), .A2(new_n934), .B1(new_n320), .B2(new_n935), .ZN(G1347gat));
  NOR3_X1   g735(.A1(new_n838), .A2(new_n664), .A3(new_n460), .ZN(new_n937));
  INV_X1    g736(.A(new_n456), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n522), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n660), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g742(.A1(new_n939), .A2(new_n636), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n230), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(new_n207), .B2(new_n944), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT60), .Z(G1350gat));
  NAND2_X1  g746(.A1(new_n939), .A2(new_n697), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G190gat), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT126), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n949), .A2(KEYINPUT126), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n949), .A2(KEYINPUT126), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(KEYINPUT61), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n206), .A3(new_n697), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n952), .A2(new_n955), .A3(new_n956), .ZN(G1351gat));
  INV_X1    g756(.A(G197gat), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n725), .A2(new_n664), .A3(new_n460), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n926), .A2(new_n522), .A3(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n962), .B1(new_n961), .B2(new_n960), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n937), .A2(new_n691), .A3(new_n676), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n958), .A3(new_n522), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1352gat));
  INV_X1    g765(.A(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n967), .A3(new_n660), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT62), .Z(new_n969));
  NAND3_X1  g768(.A1(new_n926), .A2(new_n660), .A3(new_n959), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n969), .B1(new_n971), .B2(new_n967), .ZN(G1353gat));
  INV_X1    g771(.A(G211gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n964), .A2(new_n973), .A3(new_n636), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n926), .A2(new_n636), .A3(new_n959), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  NAND3_X1  g777(.A1(new_n964), .A2(new_n524), .A3(new_n697), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n926), .A2(new_n697), .A3(new_n959), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n979), .B1(new_n981), .B2(new_n524), .ZN(G1355gat));
endmodule


