//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT79), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT0), .B(G128), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n193), .A2(new_n195), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(G128), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n193), .B(new_n195), .C1(KEYINPUT1), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  MUX2_X1   g023(.A(new_n201), .B(new_n208), .S(new_n209), .Z(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT81), .B(G224), .ZN(new_n211));
  INV_X1    g025(.A(G953), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT7), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n210), .B(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT77), .ZN(new_n216));
  XNOR2_X1  g030(.A(G104), .B(G107), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G107), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G104), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G107), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT77), .A3(G101), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT3), .B1(new_n222), .B2(G107), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n220), .A3(G104), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n226), .A2(new_n228), .A3(new_n223), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n219), .A2(new_n225), .B1(new_n229), .B2(new_n218), .ZN(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G116), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT2), .B(G113), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT80), .A2(KEYINPUT5), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT80), .A2(KEYINPUT5), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n233), .A2(G119), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n238), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n232), .B(new_n234), .C1(new_n240), .C2(new_n241), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n237), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT82), .B1(new_n230), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n219), .A2(new_n225), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n226), .A2(new_n228), .A3(new_n218), .A4(new_n223), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT82), .ZN(new_n251));
  OR2_X1    g065(.A1(KEYINPUT80), .A2(KEYINPUT5), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n243), .A2(new_n252), .A3(new_n239), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n245), .A2(new_n253), .A3(G113), .ZN(new_n254));
  OR2_X1    g068(.A1(new_n235), .A2(new_n236), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n250), .A2(new_n251), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n253), .B(G113), .C1(new_n258), .C2(new_n235), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n248), .A2(new_n255), .A3(new_n259), .A4(new_n249), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n247), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G110), .B(G122), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT8), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n261), .A2(KEYINPUT83), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT83), .B1(new_n261), .B2(new_n263), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n215), .B(KEYINPUT84), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n226), .A2(new_n228), .A3(new_n223), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G101), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n268), .A2(KEYINPUT4), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n235), .B(new_n236), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(KEYINPUT4), .A3(new_n249), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(new_n256), .B2(new_n250), .ZN(new_n273));
  INV_X1    g087(.A(new_n262), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n266), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n248), .A2(new_n249), .B1(new_n254), .B2(new_n255), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n260), .B1(new_n277), .B2(new_n251), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n230), .A2(new_n246), .A3(KEYINPUT82), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n263), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT83), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n261), .A2(KEYINPUT83), .A3(new_n263), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT84), .B1(new_n284), .B2(new_n215), .ZN(new_n285));
  OAI211_X1 g099(.A(KEYINPUT85), .B(new_n191), .C1(new_n276), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n275), .A2(KEYINPUT6), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n273), .A2(new_n274), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n210), .B(new_n213), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n215), .B1(new_n264), .B2(new_n265), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT84), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n275), .A3(new_n266), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT85), .B1(new_n296), .B2(new_n191), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n190), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n191), .B1(new_n276), .B2(new_n285), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT85), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n301), .A2(new_n189), .A3(new_n291), .A4(new_n286), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n188), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT86), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT11), .ZN(new_n306));
  INV_X1    g120(.A(G134), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(G137), .ZN(new_n308));
  INV_X1    g122(.A(G137), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT11), .A3(G134), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(G137), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G131), .ZN(new_n313));
  INV_X1    g127(.A(G131), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n308), .A2(new_n310), .A3(new_n314), .A4(new_n311), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n201), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n235), .A2(new_n236), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(new_n237), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT64), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n309), .A3(G134), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT64), .B1(new_n307), .B2(G137), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n309), .A2(G134), .ZN(new_n323));
  OAI211_X1 g137(.A(G131), .B(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n204), .A2(new_n324), .A3(new_n315), .A4(new_n206), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n317), .A2(new_n319), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(KEYINPUT28), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT67), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n317), .A2(new_n325), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(new_n270), .ZN(new_n331));
  AOI211_X1 g145(.A(KEYINPUT67), .B(new_n319), .C1(new_n317), .C2(new_n325), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n328), .B1(new_n333), .B2(KEYINPUT28), .ZN(new_n334));
  XOR2_X1   g148(.A(KEYINPUT26), .B(G101), .Z(new_n335));
  NOR2_X1   g149(.A1(G237), .A2(G953), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G210), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n335), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n305), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT30), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n342), .A2(KEYINPUT65), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(KEYINPUT65), .ZN(new_n344));
  INV_X1    g158(.A(new_n325), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n200), .B1(new_n315), .B2(new_n313), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n343), .B(new_n344), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n317), .A2(KEYINPUT65), .A3(new_n342), .A4(new_n325), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n270), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n340), .A3(new_n326), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT31), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n350), .A2(KEYINPUT31), .A3(new_n340), .A4(new_n326), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n328), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n270), .B1(new_n345), .B2(new_n346), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT67), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n330), .A2(new_n329), .A3(new_n270), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n327), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n356), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n340), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(KEYINPUT68), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n341), .A2(new_n355), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(G472), .A2(G902), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(KEYINPUT32), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT71), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n365), .A2(new_n369), .A3(KEYINPUT32), .A4(new_n366), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT69), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n366), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT32), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI211_X1 g188(.A(KEYINPUT69), .B(KEYINPUT32), .C1(new_n365), .C2(new_n366), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n368), .B(new_n370), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G472), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n334), .A2(new_n340), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n378), .A2(KEYINPUT70), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(KEYINPUT70), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n350), .A2(new_n326), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n363), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n379), .A2(new_n380), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n357), .A2(new_n326), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(new_n361), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(new_n328), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n363), .A2(new_n380), .ZN(new_n388));
  AOI21_X1  g202(.A(G902), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n377), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n376), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G125), .B(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT16), .ZN(new_n393));
  INV_X1    g207(.A(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G125), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n395), .A2(KEYINPUT16), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n393), .A2(G146), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n209), .A2(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT75), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT75), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n403), .A3(new_n192), .ZN(new_n404));
  XOR2_X1   g218(.A(KEYINPUT24), .B(G110), .Z(new_n405));
  NAND2_X1  g219(.A1(new_n231), .A2(G128), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n205), .A2(G119), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT73), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT73), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n405), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .ZN(new_n413));
  INV_X1    g227(.A(new_n407), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n406), .B(new_n413), .C1(new_n414), .C2(KEYINPUT23), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G110), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n398), .B(new_n404), .C1(new_n412), .C2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n409), .A2(new_n411), .A3(new_n405), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(G110), .ZN(new_n419));
  AOI21_X1  g233(.A(G146), .B1(new_n393), .B2(new_n396), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n418), .B(new_n419), .C1(new_n397), .C2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT74), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n421), .A2(new_n422), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n417), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT22), .B(G137), .ZN(new_n426));
  INV_X1    g240(.A(G221), .ZN(new_n427));
  INV_X1    g241(.A(G234), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n427), .A2(new_n428), .A3(G953), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n426), .B(new_n429), .Z(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n417), .B(new_n430), .C1(new_n423), .C2(new_n424), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n191), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT25), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT25), .A4(new_n191), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G217), .B1(new_n428), .B2(G902), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT72), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n432), .A2(new_n433), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n440), .A2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n441), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n391), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G469), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT10), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n250), .B2(new_n207), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n269), .A2(new_n201), .A3(new_n271), .ZN(new_n451));
  INV_X1    g265(.A(new_n316), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n230), .A2(KEYINPUT10), .A3(new_n208), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n212), .A2(G227), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT76), .ZN(new_n456));
  XNOR2_X1  g270(.A(G110), .B(G140), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT78), .B1(new_n230), .B2(new_n208), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT78), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n250), .A2(new_n461), .A3(new_n207), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n250), .A2(new_n207), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(KEYINPUT12), .A3(new_n316), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT12), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n464), .B1(new_n460), .B2(new_n462), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n468), .B1(new_n469), .B2(new_n452), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n459), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n316), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n458), .B1(new_n473), .B2(new_n454), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n448), .B(new_n191), .C1(new_n471), .C2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n448), .A2(new_n191), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n458), .A3(new_n454), .ZN(new_n478));
  INV_X1    g292(.A(new_n454), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n467), .B2(new_n470), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n478), .B1(new_n480), .B2(new_n458), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n475), .B(new_n477), .C1(new_n481), .C2(new_n448), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT9), .B(G234), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n427), .B1(new_n484), .B2(new_n191), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G113), .B(G122), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT93), .B(G104), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n488), .B(new_n489), .Z(new_n490));
  NOR2_X1   g304(.A1(new_n397), .A2(new_n420), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(new_n194), .ZN(new_n493));
  NOR2_X1   g307(.A1(KEYINPUT87), .A2(G143), .ZN(new_n494));
  OAI211_X1 g308(.A(G214), .B(new_n336), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n336), .A2(G214), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n492), .B2(new_n194), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n314), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT17), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n495), .A2(new_n497), .A3(new_n314), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n501), .A2(new_n498), .A3(KEYINPUT17), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n401), .A2(new_n403), .A3(new_n192), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n392), .B2(new_n192), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n400), .A2(KEYINPUT88), .A3(G146), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n505), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n508), .A2(new_n509), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(KEYINPUT89), .A3(new_n404), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT92), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT18), .A2(G131), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n495), .A2(new_n497), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT91), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n495), .A2(new_n497), .A3(new_n518), .A4(new_n521), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n520), .A2(new_n522), .B1(KEYINPUT18), .B2(new_n498), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n514), .A2(new_n515), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n515), .B1(new_n514), .B2(new_n523), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n490), .B(new_n504), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT19), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n401), .A2(new_n403), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n527), .B2(new_n392), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(G146), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n398), .B1(new_n501), .B2(new_n498), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT89), .B1(new_n512), .B2(new_n404), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n506), .A2(new_n510), .A3(new_n505), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n523), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT92), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n514), .A2(new_n515), .A3(new_n523), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n526), .B1(new_n538), .B2(new_n490), .ZN(new_n539));
  NOR2_X1   g353(.A1(G475), .A2(G902), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT20), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n536), .A2(new_n537), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n490), .B1(new_n545), .B2(new_n504), .ZN(new_n546));
  INV_X1    g360(.A(new_n490), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n547), .B(new_n503), .C1(new_n536), .C2(new_n537), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n191), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n542), .A2(new_n544), .B1(G475), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT94), .B1(new_n205), .B2(G143), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n194), .A3(G128), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT13), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n554), .A2(new_n555), .B1(new_n205), .B2(G143), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT95), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n554), .B2(new_n555), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n554), .A2(new_n557), .A3(new_n555), .ZN(new_n560));
  OAI21_X1  g374(.A(G134), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n554), .B(new_n307), .C1(G128), .C2(new_n194), .ZN(new_n562));
  XNOR2_X1  g376(.A(G116), .B(G122), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(new_n220), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT14), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n233), .A2(KEYINPUT14), .A3(G122), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(G107), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT96), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n554), .B1(G128), .B2(new_n194), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G134), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n573), .A2(new_n562), .B1(new_n220), .B2(new_n563), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n484), .A2(G217), .A3(new_n212), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n577), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n565), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G478), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(KEYINPUT15), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n581), .B(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n550), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(KEYINPUT97), .A2(G952), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(KEYINPUT97), .A2(G952), .ZN(new_n590));
  AOI21_X1  g404(.A(G953), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G237), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n591), .B1(new_n428), .B2(new_n592), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n191), .B(new_n212), .C1(G234), .C2(G237), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT21), .B(G898), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT98), .B1(new_n587), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n599));
  INV_X1    g413(.A(new_n597), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n550), .A2(new_n599), .A3(new_n600), .A4(new_n586), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n487), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n304), .A2(new_n447), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  OAI211_X1 g418(.A(KEYINPUT99), .B(new_n190), .C1(new_n292), .C2(new_n297), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n605), .A2(new_n187), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n298), .A2(new_n607), .A3(new_n302), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n365), .A2(new_n191), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n372), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n446), .A2(new_n487), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n600), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n549), .A2(G475), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n539), .A2(new_n543), .A3(new_n540), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n543), .B1(new_n539), .B2(new_n540), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n578), .A2(new_n580), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT33), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n578), .A2(new_n622), .A3(new_n580), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(G478), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n582), .A2(new_n191), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n581), .B2(new_n582), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n619), .A2(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n609), .A2(new_n615), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT34), .B(G104), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  INV_X1    g445(.A(new_n608), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n616), .B(new_n585), .C1(new_n617), .C2(new_n618), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n633), .B1(new_n634), .B2(new_n597), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n550), .A2(KEYINPUT100), .A3(new_n600), .A4(new_n585), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n605), .A2(new_n187), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n632), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n613), .A3(new_n614), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n431), .A2(KEYINPUT36), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n425), .A2(KEYINPUT101), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n425), .A2(KEYINPUT101), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n647), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(new_n643), .A3(new_n645), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n445), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n440), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n436), .B2(new_n437), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n612), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n304), .A2(new_n602), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT102), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(G12));
  NOR2_X1   g473(.A1(new_n487), .A2(new_n654), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n660), .B1(new_n376), .B2(new_n390), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n609), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n593), .B(KEYINPUT103), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n664), .B1(new_n665), .B2(new_n594), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n634), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  INV_X1    g483(.A(new_n487), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n666), .B(KEYINPUT39), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT40), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n673), .A2(KEYINPUT104), .ZN(new_n674));
  INV_X1    g488(.A(new_n382), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n363), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(G902), .B1(new_n385), .B2(new_n363), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n377), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n376), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n673), .B2(KEYINPUT104), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n298), .A2(KEYINPUT38), .A3(new_n302), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT38), .B1(new_n298), .B2(new_n302), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n550), .A2(new_n586), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n686), .A2(new_n187), .A3(new_n654), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n674), .A2(new_n681), .A3(new_n685), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G143), .ZN(G45));
  NOR2_X1   g503(.A1(new_n632), .A2(new_n638), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n372), .A2(new_n373), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT69), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n372), .A2(new_n371), .A3(new_n373), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n368), .A2(new_n370), .ZN(new_n695));
  INV_X1    g509(.A(new_n390), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n628), .A2(new_n666), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n690), .A2(new_n697), .A3(new_n660), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  NOR2_X1   g514(.A1(new_n609), .A2(new_n628), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n471), .A2(new_n474), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n191), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n448), .A2(KEYINPUT105), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n702), .B(new_n191), .C1(KEYINPUT105), .C2(new_n448), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n705), .A2(new_n486), .A3(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n701), .A2(new_n447), .A3(new_n600), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT41), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G113), .ZN(G15));
  NAND3_X1  g524(.A1(new_n447), .A2(new_n639), .A3(new_n707), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  AOI21_X1  g526(.A(new_n654), .B1(new_n598), .B2(new_n601), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n690), .A2(new_n697), .A3(new_n707), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  AOI21_X1  g529(.A(new_n653), .B1(new_n442), .B2(new_n444), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n355), .B1(new_n340), .B2(new_n387), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n366), .ZN(new_n718));
  AOI21_X1  g532(.A(KEYINPUT106), .B1(new_n610), .B2(G472), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n720));
  AOI211_X1 g534(.A(new_n720), .B(new_n377), .C1(new_n365), .C2(new_n191), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n716), .B(new_n718), .C1(new_n719), .C2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n707), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n597), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n690), .A2(new_n724), .A3(new_n686), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NAND4_X1  g540(.A1(new_n608), .A2(new_n187), .A3(new_n605), .A4(new_n707), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n611), .A2(new_n720), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n610), .A2(KEYINPUT106), .A3(G472), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n643), .B1(new_n649), .B2(new_n645), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n646), .A2(new_n647), .A3(new_n644), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n444), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n441), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n730), .A2(new_n698), .A3(new_n734), .A4(new_n718), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n727), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n209), .ZN(G27));
  NAND3_X1  g551(.A1(new_n696), .A2(new_n691), .A3(new_n367), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n716), .A3(new_n698), .ZN(new_n739));
  AND4_X1   g553(.A1(new_n298), .A2(new_n302), .A3(new_n187), .A4(new_n670), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT42), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n698), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(KEYINPUT42), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n697), .A3(new_n716), .A4(new_n740), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n314), .ZN(G33));
  NAND4_X1  g561(.A1(new_n697), .A2(new_n740), .A3(new_n716), .A4(new_n667), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  NAND3_X1  g563(.A1(new_n298), .A2(new_n302), .A3(new_n187), .ZN(new_n750));
  INV_X1    g564(.A(new_n627), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT43), .B1(new_n619), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n550), .A2(new_n753), .A3(new_n627), .ZN(new_n754));
  AND4_X1   g568(.A1(new_n612), .A2(new_n752), .A3(new_n754), .A4(new_n734), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n750), .B1(new_n755), .B2(KEYINPUT44), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n448), .B1(new_n481), .B2(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(KEYINPUT45), .B(new_n478), .C1(new_n480), .C2(new_n458), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n476), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n475), .B1(new_n760), .B2(KEYINPUT46), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n762), .B(new_n476), .C1(new_n758), .C2(new_n759), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n486), .B(new_n671), .C1(new_n761), .C2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n756), .B(new_n765), .C1(KEYINPUT44), .C2(new_n755), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  OAI21_X1  g581(.A(new_n486), .B1(new_n761), .B2(new_n763), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(KEYINPUT47), .B(new_n486), .C1(new_n761), .C2(new_n763), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n697), .A2(new_n716), .A3(new_n743), .ZN(new_n773));
  INV_X1    g587(.A(new_n750), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n736), .B1(new_n662), .B2(new_n667), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n734), .B2(new_n666), .ZN(new_n781));
  INV_X1    g595(.A(new_n666), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n654), .A2(KEYINPUT109), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n487), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n376), .B2(new_n679), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n606), .A2(new_n608), .A3(new_n686), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n778), .A2(new_n779), .A3(new_n699), .A4(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n697), .A2(new_n608), .A3(new_n606), .A4(new_n660), .ZN(new_n789));
  INV_X1    g603(.A(new_n667), .ZN(new_n790));
  OAI22_X1  g604(.A1(new_n789), .A2(new_n790), .B1(new_n727), .B2(new_n735), .ZN(new_n791));
  OAI22_X1  g605(.A1(new_n789), .A2(new_n743), .B1(new_n786), .B2(new_n785), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT52), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n587), .A2(new_n487), .A3(new_n654), .A4(new_n666), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n697), .A2(new_n774), .A3(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n734), .B(new_n718), .C1(new_n719), .C2(new_n721), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n740), .A3(new_n698), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n748), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n746), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n788), .A2(new_n793), .A3(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n711), .A2(new_n714), .ZN(new_n802));
  INV_X1    g616(.A(new_n615), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n634), .A2(KEYINPUT108), .B1(new_n619), .B2(new_n627), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(KEYINPUT108), .B2(new_n634), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n298), .A2(new_n302), .ZN(new_n806));
  INV_X1    g620(.A(new_n188), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT86), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT86), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n809), .B(new_n188), .C1(new_n298), .C2(new_n302), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n803), .B(new_n805), .C1(new_n808), .C2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n725), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n304), .B(new_n602), .C1(new_n447), .C2(new_n655), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n802), .A2(new_n708), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n777), .B1(new_n801), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n795), .A2(new_n798), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n742), .A3(new_n745), .A4(new_n748), .ZN(new_n817));
  INV_X1    g631(.A(new_n736), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n668), .A2(new_n787), .A3(new_n699), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n817), .B1(new_n819), .B2(KEYINPUT52), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n813), .A2(new_n708), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n711), .A2(new_n714), .A3(new_n811), .A4(new_n725), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n820), .A2(KEYINPUT53), .A3(new_n823), .A4(new_n788), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n815), .A2(KEYINPUT54), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT54), .B1(new_n815), .B2(new_n824), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n367), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n390), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n446), .B1(new_n829), .B2(new_n691), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n707), .A2(new_n298), .A3(new_n302), .A4(new_n187), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n752), .A2(new_n754), .A3(new_n664), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT48), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n446), .A2(new_n593), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n680), .A2(new_n832), .A3(KEYINPUT110), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT110), .ZN(new_n838));
  INV_X1    g652(.A(new_n679), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n694), .A2(new_n695), .A3(new_n839), .A4(new_n836), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n840), .B2(new_n831), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n837), .A2(new_n841), .A3(new_n619), .A4(new_n627), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n752), .A2(new_n754), .A3(new_n664), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n722), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n690), .A2(new_n707), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n845), .A2(new_n591), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n835), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n705), .A2(new_n706), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n485), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n770), .A2(new_n771), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n843), .A2(new_n722), .A3(new_n750), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n723), .A2(new_n187), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n684), .A2(new_n844), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n682), .B2(new_n683), .ZN(new_n857));
  INV_X1    g671(.A(new_n722), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n833), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT50), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n832), .A2(new_n797), .A3(new_n833), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n853), .A2(new_n856), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n550), .A2(new_n751), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n837), .A2(new_n841), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT111), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n837), .A2(new_n841), .A3(KEYINPUT111), .A4(new_n864), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n862), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n848), .B1(new_n869), .B2(KEYINPUT51), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n868), .ZN(new_n871));
  AND4_X1   g685(.A1(KEYINPUT51), .A2(new_n856), .A3(new_n860), .A4(new_n861), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n851), .A2(KEYINPUT112), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n851), .A2(KEYINPUT112), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n852), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n871), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT113), .B1(new_n870), .B2(new_n877), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n856), .A2(new_n853), .A3(new_n861), .A4(new_n860), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n871), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT51), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n847), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT113), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n882), .A2(new_n883), .A3(new_n876), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT114), .B1(new_n827), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n815), .A2(new_n824), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n815), .A2(new_n824), .A3(KEYINPUT54), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n870), .A2(KEYINPUT113), .A3(new_n877), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n883), .B1(new_n882), .B2(new_n876), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT114), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(G952), .A2(G953), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n886), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n446), .A2(new_n188), .A3(new_n485), .ZN(new_n899));
  INV_X1    g713(.A(new_n849), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n899), .A2(KEYINPUT107), .B1(new_n900), .B2(KEYINPUT49), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(KEYINPUT49), .B2(new_n900), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n550), .B(new_n627), .C1(new_n899), .C2(KEYINPUT107), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(new_n684), .A3(new_n680), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n898), .A2(new_n905), .ZN(G75));
  NOR2_X1   g720(.A1(new_n212), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n191), .B1(new_n815), .B2(new_n824), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT56), .B1(new_n909), .B2(G210), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n289), .B(KEYINPUT115), .Z(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT116), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n290), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n908), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n909), .A2(new_n916), .A3(G210), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n916), .B1(new_n909), .B2(G210), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT118), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n909), .A2(G210), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT117), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n924), .A2(new_n925), .A3(new_n917), .A4(new_n919), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n915), .B1(new_n922), .B2(new_n926), .ZN(G51));
  XOR2_X1   g741(.A(new_n476), .B(KEYINPUT57), .Z(new_n928));
  OAI21_X1  g742(.A(new_n702), .B1(new_n891), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n758), .A2(new_n759), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT119), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n909), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n907), .B1(new_n929), .B2(new_n932), .ZN(G54));
  AND2_X1   g747(.A1(KEYINPUT58), .A2(G475), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n909), .A2(new_n539), .A3(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(KEYINPUT120), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(KEYINPUT120), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n539), .B1(new_n909), .B2(new_n934), .ZN(new_n938));
  NOR4_X1   g752(.A1(new_n936), .A2(new_n937), .A3(new_n907), .A4(new_n938), .ZN(G60));
  NAND2_X1  g753(.A1(new_n621), .A2(new_n623), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n625), .B(KEYINPUT59), .Z(new_n941));
  AND3_X1   g755(.A1(new_n827), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n827), .B2(new_n941), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n907), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT60), .Z(new_n946));
  NAND2_X1  g760(.A1(new_n887), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n731), .A2(new_n732), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n907), .B1(new_n947), .B2(new_n443), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n949), .A2(KEYINPUT61), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(G66));
  INV_X1    g769(.A(new_n211), .ZN(new_n956));
  OAI21_X1  g770(.A(G953), .B1(new_n956), .B2(new_n595), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n823), .B(KEYINPUT121), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(G953), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n911), .B1(G898), .B2(new_n212), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT122), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT123), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n959), .B(new_n962), .ZN(G69));
  AOI21_X1  g777(.A(new_n791), .B1(new_n662), .B2(new_n698), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n688), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT62), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(new_n967), .A3(new_n688), .ZN(new_n968));
  INV_X1    g782(.A(new_n672), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n447), .A2(new_n969), .A3(new_n774), .A4(new_n805), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n766), .A2(new_n775), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n966), .A2(new_n968), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n212), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n349), .B(new_n529), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n974), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n212), .A2(G900), .ZN(new_n977));
  INV_X1    g791(.A(new_n746), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n690), .A2(new_n765), .A3(new_n686), .A4(new_n830), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(new_n748), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n971), .A2(new_n964), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n977), .B1(new_n981), .B2(new_n212), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT125), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n976), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n975), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT124), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n985), .B2(new_n984), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n212), .B1(G227), .B2(G900), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n986), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  OAI221_X1 g805(.A(new_n975), .B1(new_n987), .B2(new_n989), .C1(new_n984), .C2(new_n985), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n991), .A2(new_n992), .ZN(G72));
  XNOR2_X1  g807(.A(new_n814), .B(KEYINPUT121), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n994), .A2(new_n972), .ZN(new_n995));
  NAND2_X1  g809(.A1(G472), .A2(G902), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT63), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n676), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(new_n383), .B2(new_n351), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT127), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n887), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n981), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n997), .B1(new_n958), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n675), .A2(new_n363), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n908), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1006), .A2(KEYINPUT126), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(KEYINPUT126), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1002), .B1(new_n1007), .B2(new_n1008), .ZN(G57));
endmodule


