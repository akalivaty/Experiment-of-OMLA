

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U555 ( .A(G2105), .ZN(n526) );
  XOR2_X1 U556 ( .A(KEYINPUT64), .B(n527), .Z(n518) );
  AND2_X1 U557 ( .A1(n830), .A2(n829), .ZN(n519) );
  XOR2_X1 U558 ( .A(n822), .B(KEYINPUT96), .Z(n520) );
  AND2_X1 U559 ( .A1(n742), .A2(n741), .ZN(n745) );
  INV_X1 U560 ( .A(KEYINPUT94), .ZN(n743) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n761) );
  XNOR2_X1 U562 ( .A(n762), .B(n761), .ZN(n767) );
  NOR2_X1 U563 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U564 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U565 ( .A1(n731), .A2(n730), .ZN(n781) );
  NAND2_X1 U566 ( .A1(n797), .A2(n796), .ZN(n816) );
  NOR2_X1 U567 ( .A1(G651), .A2(n646), .ZN(n651) );
  NOR2_X1 U568 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U569 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U570 ( .A1(n531), .A2(n530), .ZN(G160) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n876) );
  NAND2_X1 U572 ( .A1(n876), .A2(G113), .ZN(n523) );
  NOR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XOR2_X1 U574 ( .A(KEYINPUT17), .B(n521), .Z(n867) );
  NAND2_X1 U575 ( .A1(n867), .A2(G137), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n523), .A2(n522), .ZN(n531) );
  NAND2_X1 U577 ( .A1(n526), .A2(G2104), .ZN(n524) );
  XNOR2_X2 U578 ( .A(n524), .B(KEYINPUT65), .ZN(n869) );
  NAND2_X1 U579 ( .A1(n869), .A2(G101), .ZN(n525) );
  XNOR2_X1 U580 ( .A(n525), .B(KEYINPUT23), .ZN(n528) );
  NOR2_X2 U581 ( .A1(G2104), .A2(n526), .ZN(n873) );
  NAND2_X1 U582 ( .A1(n873), .A2(G125), .ZN(n527) );
  NOR2_X1 U583 ( .A1(n528), .A2(n518), .ZN(n529) );
  XOR2_X1 U584 ( .A(KEYINPUT66), .B(n529), .Z(n530) );
  NOR2_X1 U585 ( .A1(G651), .A2(G543), .ZN(n637) );
  NAND2_X1 U586 ( .A1(G85), .A2(n637), .ZN(n533) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n646) );
  INV_X1 U588 ( .A(G651), .ZN(n534) );
  NOR2_X1 U589 ( .A1(n646), .A2(n534), .ZN(n640) );
  NAND2_X1 U590 ( .A1(G72), .A2(n640), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n533), .A2(n532), .ZN(n540) );
  NAND2_X1 U592 ( .A1(G47), .A2(n651), .ZN(n538) );
  XNOR2_X1 U593 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n536) );
  NOR2_X1 U594 ( .A1(G543), .A2(n534), .ZN(n535) );
  XNOR2_X1 U595 ( .A(n536), .B(n535), .ZN(n650) );
  NAND2_X1 U596 ( .A1(G60), .A2(n650), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n538), .A2(n537), .ZN(n539) );
  OR2_X1 U598 ( .A1(n540), .A2(n539), .ZN(G290) );
  XOR2_X1 U599 ( .A(G2438), .B(G2454), .Z(n542) );
  XNOR2_X1 U600 ( .A(G2435), .B(G2430), .ZN(n541) );
  XNOR2_X1 U601 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U602 ( .A(n543), .B(G2427), .Z(n545) );
  XNOR2_X1 U603 ( .A(G1348), .B(G1341), .ZN(n544) );
  XNOR2_X1 U604 ( .A(n545), .B(n544), .ZN(n549) );
  XOR2_X1 U605 ( .A(G2443), .B(G2446), .Z(n547) );
  XNOR2_X1 U606 ( .A(KEYINPUT100), .B(G2451), .ZN(n546) );
  XNOR2_X1 U607 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U608 ( .A(n549), .B(n548), .Z(n550) );
  AND2_X1 U609 ( .A1(G14), .A2(n550), .ZN(G401) );
  NAND2_X1 U610 ( .A1(G52), .A2(n651), .ZN(n552) );
  NAND2_X1 U611 ( .A1(G64), .A2(n650), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n552), .A2(n551), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n637), .A2(G90), .ZN(n553) );
  XNOR2_X1 U614 ( .A(n553), .B(KEYINPUT68), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G77), .A2(n640), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U617 ( .A(KEYINPUT69), .B(n556), .ZN(n557) );
  XNOR2_X1 U618 ( .A(KEYINPUT9), .B(n557), .ZN(n558) );
  NOR2_X1 U619 ( .A1(n559), .A2(n558), .ZN(G171) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G69), .ZN(G235) );
  NAND2_X1 U622 ( .A1(n637), .A2(G89), .ZN(n560) );
  XNOR2_X1 U623 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  NAND2_X1 U624 ( .A1(G76), .A2(n640), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U626 ( .A(KEYINPUT5), .B(n563), .ZN(n569) );
  NAND2_X1 U627 ( .A1(n650), .A2(G63), .ZN(n564) );
  XOR2_X1 U628 ( .A(KEYINPUT75), .B(n564), .Z(n566) );
  NAND2_X1 U629 ( .A1(n651), .A2(G51), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U631 ( .A(KEYINPUT6), .B(n567), .Z(n568) );
  NAND2_X1 U632 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U633 ( .A(KEYINPUT7), .B(n570), .ZN(G168) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n835) );
  NAND2_X1 U638 ( .A1(n835), .A2(G567), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n572), .Z(G234) );
  NAND2_X1 U640 ( .A1(G56), .A2(n650), .ZN(n573) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n573), .Z(n579) );
  NAND2_X1 U642 ( .A1(n637), .A2(G81), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n574), .B(KEYINPUT12), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G68), .A2(n640), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U646 ( .A(KEYINPUT13), .B(n577), .Z(n578) );
  NOR2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n651), .A2(G43), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n970) );
  INV_X1 U650 ( .A(G860), .ZN(n621) );
  OR2_X1 U651 ( .A1(n970), .A2(n621), .ZN(G153) );
  INV_X1 U652 ( .A(G868), .ZN(n662) );
  NOR2_X1 U653 ( .A1(n662), .A2(G171), .ZN(n582) );
  XNOR2_X1 U654 ( .A(n582), .B(KEYINPUT73), .ZN(n592) );
  NAND2_X1 U655 ( .A1(G92), .A2(n637), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G54), .A2(n651), .ZN(n584) );
  NAND2_X1 U657 ( .A1(G66), .A2(n650), .ZN(n583) );
  NAND2_X1 U658 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n640), .A2(G79), .ZN(n585) );
  XOR2_X1 U660 ( .A(KEYINPUT74), .B(n585), .Z(n586) );
  NOR2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT15), .ZN(n974) );
  OR2_X1 U664 ( .A1(G868), .A2(n974), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(G284) );
  NAND2_X1 U666 ( .A1(G91), .A2(n637), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G78), .A2(n640), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n650), .A2(G65), .ZN(n595) );
  XNOR2_X1 U670 ( .A(n595), .B(KEYINPUT70), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G53), .A2(n651), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U673 ( .A(KEYINPUT71), .B(n598), .Z(n599) );
  XOR2_X1 U674 ( .A(KEYINPUT72), .B(n601), .Z(G299) );
  NOR2_X1 U675 ( .A1(G286), .A2(n662), .ZN(n603) );
  NOR2_X1 U676 ( .A1(G299), .A2(G868), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n621), .A2(G559), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n604), .A2(n974), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n970), .ZN(n608) );
  NAND2_X1 U682 ( .A1(G868), .A2(n974), .ZN(n606) );
  NOR2_X1 U683 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U684 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G123), .A2(n873), .ZN(n609) );
  XNOR2_X1 U686 ( .A(n609), .B(KEYINPUT76), .ZN(n610) );
  XNOR2_X1 U687 ( .A(KEYINPUT18), .B(n610), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G135), .A2(n867), .ZN(n611) );
  XOR2_X1 U689 ( .A(KEYINPUT77), .B(n611), .Z(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U691 ( .A1(G99), .A2(n869), .ZN(n615) );
  NAND2_X1 U692 ( .A1(G111), .A2(n876), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n917) );
  XNOR2_X1 U695 ( .A(G2096), .B(n917), .ZN(n619) );
  INV_X1 U696 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U698 ( .A1(G559), .A2(n974), .ZN(n620) );
  XOR2_X1 U699 ( .A(n970), .B(n620), .Z(n660) );
  NAND2_X1 U700 ( .A1(n621), .A2(n660), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G93), .A2(n637), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G80), .A2(n640), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n650), .A2(G67), .ZN(n624) );
  XOR2_X1 U705 ( .A(KEYINPUT78), .B(n624), .Z(n625) );
  NOR2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n651), .A2(G55), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n663) );
  XNOR2_X1 U709 ( .A(n629), .B(n663), .ZN(G145) );
  NAND2_X1 U710 ( .A1(G88), .A2(n637), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G75), .A2(n640), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G50), .A2(n651), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G62), .A2(n650), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U716 ( .A1(n635), .A2(n634), .ZN(G166) );
  NAND2_X1 U717 ( .A1(G61), .A2(n650), .ZN(n636) );
  XNOR2_X1 U718 ( .A(n636), .B(KEYINPUT80), .ZN(n645) );
  NAND2_X1 U719 ( .A1(G48), .A2(n651), .ZN(n639) );
  NAND2_X1 U720 ( .A1(G86), .A2(n637), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n640), .A2(G73), .ZN(n641) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n641), .Z(n642) );
  NOR2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U726 ( .A1(G87), .A2(n646), .ZN(n648) );
  NAND2_X1 U727 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U730 ( .A1(G49), .A2(n651), .ZN(n652) );
  XOR2_X1 U731 ( .A(KEYINPUT79), .B(n652), .Z(n653) );
  NAND2_X1 U732 ( .A1(n654), .A2(n653), .ZN(G288) );
  XNOR2_X1 U733 ( .A(G166), .B(KEYINPUT19), .ZN(n659) );
  XNOR2_X1 U734 ( .A(G299), .B(G305), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n655), .B(n663), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(G288), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n657), .B(G290), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n659), .B(n658), .ZN(n885) );
  XOR2_X1 U739 ( .A(n885), .B(n660), .Z(n661) );
  NOR2_X1 U740 ( .A1(n662), .A2(n661), .ZN(n665) );
  NOR2_X1 U741 ( .A1(G868), .A2(n663), .ZN(n664) );
  NOR2_X1 U742 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XNOR2_X1 U744 ( .A(n666), .B(KEYINPUT81), .ZN(n667) );
  XNOR2_X1 U745 ( .A(n667), .B(KEYINPUT20), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n668), .A2(G2090), .ZN(n669) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U748 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(KEYINPUT82), .B(G44), .ZN(n671) );
  XNOR2_X1 U750 ( .A(n671), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U751 ( .A1(G120), .A2(G108), .ZN(n672) );
  NOR2_X1 U752 ( .A1(G235), .A2(n672), .ZN(n673) );
  NAND2_X1 U753 ( .A1(G57), .A2(n673), .ZN(n915) );
  NAND2_X1 U754 ( .A1(n915), .A2(G567), .ZN(n680) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(KEYINPUT83), .Z(n675) );
  NAND2_X1 U756 ( .A1(G132), .A2(G82), .ZN(n674) );
  XNOR2_X1 U757 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U758 ( .A1(n676), .A2(G218), .ZN(n677) );
  NAND2_X1 U759 ( .A1(G96), .A2(n677), .ZN(n678) );
  XNOR2_X1 U760 ( .A(KEYINPUT84), .B(n678), .ZN(n916) );
  NAND2_X1 U761 ( .A1(G2106), .A2(n916), .ZN(n679) );
  NAND2_X1 U762 ( .A1(n680), .A2(n679), .ZN(n839) );
  NAND2_X1 U763 ( .A1(G661), .A2(G483), .ZN(n681) );
  NOR2_X1 U764 ( .A1(n839), .A2(n681), .ZN(n838) );
  NAND2_X1 U765 ( .A1(n838), .A2(G36), .ZN(n682) );
  XOR2_X1 U766 ( .A(KEYINPUT85), .B(n682), .Z(G176) );
  NAND2_X1 U767 ( .A1(G114), .A2(n876), .ZN(n683) );
  XNOR2_X1 U768 ( .A(n683), .B(KEYINPUT86), .ZN(n685) );
  NAND2_X1 U769 ( .A1(n867), .A2(G138), .ZN(n684) );
  NAND2_X1 U770 ( .A1(n685), .A2(n684), .ZN(n689) );
  NAND2_X1 U771 ( .A1(G126), .A2(n873), .ZN(n687) );
  NAND2_X1 U772 ( .A1(G102), .A2(n869), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U774 ( .A1(n689), .A2(n688), .ZN(G164) );
  INV_X1 U775 ( .A(G166), .ZN(G303) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n730) );
  NAND2_X1 U777 ( .A1(G160), .A2(G40), .ZN(n729) );
  NOR2_X1 U778 ( .A1(n730), .A2(n729), .ZN(n728) );
  NAND2_X1 U779 ( .A1(G105), .A2(n869), .ZN(n690) );
  XNOR2_X1 U780 ( .A(n690), .B(KEYINPUT38), .ZN(n697) );
  NAND2_X1 U781 ( .A1(G141), .A2(n867), .ZN(n692) );
  NAND2_X1 U782 ( .A1(G117), .A2(n876), .ZN(n691) );
  NAND2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U784 ( .A1(G129), .A2(n873), .ZN(n693) );
  XNOR2_X1 U785 ( .A(KEYINPUT89), .B(n693), .ZN(n694) );
  NOR2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n859) );
  NOR2_X1 U788 ( .A1(G1996), .A2(n859), .ZN(n937) );
  NAND2_X1 U789 ( .A1(G119), .A2(n873), .ZN(n699) );
  NAND2_X1 U790 ( .A1(G107), .A2(n876), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n704) );
  NAND2_X1 U792 ( .A1(G131), .A2(n867), .ZN(n700) );
  XNOR2_X1 U793 ( .A(n700), .B(KEYINPUT88), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n869), .A2(G95), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n860) );
  INV_X1 U797 ( .A(G1991), .ZN(n952) );
  NOR2_X1 U798 ( .A1(n860), .A2(n952), .ZN(n706) );
  AND2_X1 U799 ( .A1(n859), .A2(G1996), .ZN(n705) );
  NOR2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n921) );
  INV_X1 U801 ( .A(n728), .ZN(n707) );
  NOR2_X1 U802 ( .A1(n921), .A2(n707), .ZN(n800) );
  AND2_X1 U803 ( .A1(n952), .A2(n860), .ZN(n918) );
  NOR2_X1 U804 ( .A1(G1986), .A2(G290), .ZN(n708) );
  XOR2_X1 U805 ( .A(n708), .B(KEYINPUT97), .Z(n709) );
  NOR2_X1 U806 ( .A1(n918), .A2(n709), .ZN(n710) );
  NOR2_X1 U807 ( .A1(n800), .A2(n710), .ZN(n711) );
  NOR2_X1 U808 ( .A1(n937), .A2(n711), .ZN(n712) );
  XNOR2_X1 U809 ( .A(n712), .B(KEYINPUT39), .ZN(n723) );
  NAND2_X1 U810 ( .A1(G104), .A2(n869), .ZN(n714) );
  NAND2_X1 U811 ( .A1(G140), .A2(n867), .ZN(n713) );
  NAND2_X1 U812 ( .A1(n714), .A2(n713), .ZN(n716) );
  XOR2_X1 U813 ( .A(KEYINPUT87), .B(KEYINPUT34), .Z(n715) );
  XNOR2_X1 U814 ( .A(n716), .B(n715), .ZN(n721) );
  NAND2_X1 U815 ( .A1(G128), .A2(n873), .ZN(n718) );
  NAND2_X1 U816 ( .A1(G116), .A2(n876), .ZN(n717) );
  NAND2_X1 U817 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U818 ( .A(KEYINPUT35), .B(n719), .Z(n720) );
  NOR2_X1 U819 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U820 ( .A(KEYINPUT36), .B(n722), .ZN(n849) );
  XNOR2_X1 U821 ( .A(G2067), .B(KEYINPUT37), .ZN(n724) );
  NOR2_X1 U822 ( .A1(n849), .A2(n724), .ZN(n928) );
  NAND2_X1 U823 ( .A1(n728), .A2(n928), .ZN(n801) );
  NAND2_X1 U824 ( .A1(n723), .A2(n801), .ZN(n725) );
  NAND2_X1 U825 ( .A1(n849), .A2(n724), .ZN(n929) );
  NAND2_X1 U826 ( .A1(n725), .A2(n929), .ZN(n726) );
  NAND2_X1 U827 ( .A1(n728), .A2(n726), .ZN(n727) );
  XNOR2_X1 U828 ( .A(KEYINPUT98), .B(n727), .ZN(n814) );
  XNOR2_X1 U829 ( .A(G1986), .B(G290), .ZN(n984) );
  NAND2_X1 U830 ( .A1(n984), .A2(n728), .ZN(n827) );
  INV_X1 U831 ( .A(n827), .ZN(n812) );
  INV_X1 U832 ( .A(n729), .ZN(n731) );
  NAND2_X1 U833 ( .A1(G8), .A2(n781), .ZN(n825) );
  NOR2_X1 U834 ( .A1(G1966), .A2(n825), .ZN(n776) );
  INV_X1 U835 ( .A(n781), .ZN(n732) );
  XNOR2_X1 U836 ( .A(G1996), .B(KEYINPUT92), .ZN(n948) );
  NAND2_X1 U837 ( .A1(n732), .A2(n948), .ZN(n733) );
  XNOR2_X1 U838 ( .A(n733), .B(KEYINPUT26), .ZN(n735) );
  AND2_X1 U839 ( .A1(n781), .A2(G1341), .ZN(n734) );
  NAND2_X1 U840 ( .A1(KEYINPUT26), .A2(n734), .ZN(n738) );
  NAND2_X1 U841 ( .A1(n735), .A2(n738), .ZN(n737) );
  INV_X1 U842 ( .A(KEYINPUT93), .ZN(n736) );
  NAND2_X1 U843 ( .A1(n737), .A2(n736), .ZN(n742) );
  INV_X1 U844 ( .A(n970), .ZN(n740) );
  NAND2_X1 U845 ( .A1(n738), .A2(KEYINPUT93), .ZN(n739) );
  AND2_X1 U846 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U847 ( .A1(n745), .A2(n974), .ZN(n744) );
  XNOR2_X1 U848 ( .A(n744), .B(n743), .ZN(n751) );
  NAND2_X1 U849 ( .A1(n745), .A2(n974), .ZN(n749) );
  NOR2_X1 U850 ( .A1(G2067), .A2(n781), .ZN(n747) );
  INV_X1 U851 ( .A(n781), .ZN(n763) );
  NOR2_X1 U852 ( .A1(n763), .A2(G1348), .ZN(n746) );
  NOR2_X1 U853 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U854 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U855 ( .A1(n751), .A2(n750), .ZN(n756) );
  NAND2_X1 U856 ( .A1(n763), .A2(G2072), .ZN(n752) );
  XNOR2_X1 U857 ( .A(n752), .B(KEYINPUT27), .ZN(n754) );
  INV_X1 U858 ( .A(G1956), .ZN(n999) );
  NOR2_X1 U859 ( .A1(n999), .A2(n763), .ZN(n753) );
  NOR2_X1 U860 ( .A1(n754), .A2(n753), .ZN(n757) );
  INV_X1 U861 ( .A(G299), .ZN(n975) );
  NAND2_X1 U862 ( .A1(n757), .A2(n975), .ZN(n755) );
  NAND2_X1 U863 ( .A1(n756), .A2(n755), .ZN(n760) );
  NOR2_X1 U864 ( .A1(n757), .A2(n975), .ZN(n758) );
  XOR2_X1 U865 ( .A(n758), .B(KEYINPUT28), .Z(n759) );
  NAND2_X1 U866 ( .A1(n760), .A2(n759), .ZN(n762) );
  INV_X1 U867 ( .A(G1961), .ZN(n971) );
  NAND2_X1 U868 ( .A1(n781), .A2(n971), .ZN(n765) );
  XNOR2_X1 U869 ( .A(G2078), .B(KEYINPUT25), .ZN(n946) );
  NAND2_X1 U870 ( .A1(n763), .A2(n946), .ZN(n764) );
  NAND2_X1 U871 ( .A1(n765), .A2(n764), .ZN(n771) );
  NAND2_X1 U872 ( .A1(n771), .A2(G171), .ZN(n766) );
  NAND2_X1 U873 ( .A1(n767), .A2(n766), .ZN(n789) );
  NOR2_X1 U874 ( .A1(G2084), .A2(n781), .ZN(n777) );
  NOR2_X1 U875 ( .A1(n776), .A2(n777), .ZN(n768) );
  NAND2_X1 U876 ( .A1(G8), .A2(n768), .ZN(n769) );
  XNOR2_X1 U877 ( .A(KEYINPUT30), .B(n769), .ZN(n770) );
  NOR2_X1 U878 ( .A1(G168), .A2(n770), .ZN(n773) );
  NOR2_X1 U879 ( .A1(G171), .A2(n771), .ZN(n772) );
  NOR2_X1 U880 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U881 ( .A(KEYINPUT31), .B(n774), .Z(n787) );
  AND2_X1 U882 ( .A1(n789), .A2(n787), .ZN(n775) );
  NOR2_X1 U883 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U884 ( .A1(G8), .A2(n777), .ZN(n778) );
  XOR2_X1 U885 ( .A(KEYINPUT91), .B(n778), .Z(n779) );
  NAND2_X1 U886 ( .A1(n780), .A2(n779), .ZN(n797) );
  INV_X1 U887 ( .A(G8), .ZN(n786) );
  NOR2_X1 U888 ( .A1(G1971), .A2(n825), .ZN(n783) );
  NOR2_X1 U889 ( .A1(G2090), .A2(n781), .ZN(n782) );
  NOR2_X1 U890 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U891 ( .A1(n784), .A2(G303), .ZN(n785) );
  OR2_X1 U892 ( .A1(n786), .A2(n785), .ZN(n790) );
  AND2_X1 U893 ( .A1(n787), .A2(n790), .ZN(n788) );
  NAND2_X1 U894 ( .A1(n789), .A2(n788), .ZN(n794) );
  INV_X1 U895 ( .A(n790), .ZN(n792) );
  AND2_X1 U896 ( .A1(G286), .A2(G8), .ZN(n791) );
  OR2_X1 U897 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U898 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U899 ( .A(KEYINPUT32), .B(n795), .ZN(n796) );
  NOR2_X1 U900 ( .A1(G2090), .A2(G303), .ZN(n798) );
  NAND2_X1 U901 ( .A1(G8), .A2(n798), .ZN(n799) );
  NAND2_X1 U902 ( .A1(n816), .A2(n799), .ZN(n805) );
  INV_X1 U903 ( .A(n800), .ZN(n802) );
  NAND2_X1 U904 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U905 ( .A(n803), .B(KEYINPUT90), .Z(n826) );
  AND2_X1 U906 ( .A1(n825), .A2(n826), .ZN(n804) );
  AND2_X1 U907 ( .A1(n805), .A2(n804), .ZN(n810) );
  NOR2_X1 U908 ( .A1(G1981), .A2(G305), .ZN(n806) );
  XOR2_X1 U909 ( .A(n806), .B(KEYINPUT24), .Z(n807) );
  NOR2_X1 U910 ( .A1(n825), .A2(n807), .ZN(n808) );
  AND2_X1 U911 ( .A1(n826), .A2(n808), .ZN(n809) );
  NOR2_X1 U912 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U913 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U914 ( .A1(n814), .A2(n813), .ZN(n832) );
  NOR2_X1 U915 ( .A1(G1976), .A2(G288), .ZN(n823) );
  NOR2_X1 U916 ( .A1(G1971), .A2(G303), .ZN(n815) );
  NOR2_X1 U917 ( .A1(n823), .A2(n815), .ZN(n979) );
  NAND2_X1 U918 ( .A1(n816), .A2(n979), .ZN(n817) );
  XNOR2_X1 U919 ( .A(KEYINPUT95), .B(n817), .ZN(n820) );
  NAND2_X1 U920 ( .A1(G1976), .A2(G288), .ZN(n978) );
  INV_X1 U921 ( .A(n825), .ZN(n818) );
  NAND2_X1 U922 ( .A1(n978), .A2(n818), .ZN(n819) );
  NOR2_X1 U923 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U924 ( .A1(n821), .A2(KEYINPUT33), .ZN(n822) );
  NAND2_X1 U925 ( .A1(n823), .A2(KEYINPUT33), .ZN(n824) );
  OR2_X1 U926 ( .A1(n825), .A2(n824), .ZN(n830) );
  XOR2_X1 U927 ( .A(G1981), .B(G305), .Z(n991) );
  AND2_X1 U928 ( .A1(n991), .A2(n826), .ZN(n828) );
  AND2_X1 U929 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U930 ( .A1(n520), .A2(n519), .ZN(n831) );
  NAND2_X1 U931 ( .A1(n832), .A2(n831), .ZN(n834) );
  XOR2_X1 U932 ( .A(KEYINPUT99), .B(KEYINPUT40), .Z(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U936 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U938 ( .A1(n838), .A2(n837), .ZN(G188) );
  XNOR2_X1 U939 ( .A(G120), .B(KEYINPUT101), .ZN(G236) );
  INV_X1 U940 ( .A(n839), .ZN(G319) );
  XOR2_X1 U941 ( .A(KEYINPUT104), .B(KEYINPUT44), .Z(n841) );
  NAND2_X1 U942 ( .A1(G124), .A2(n873), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n848) );
  NAND2_X1 U944 ( .A1(G100), .A2(n869), .ZN(n843) );
  NAND2_X1 U945 ( .A1(G112), .A2(n876), .ZN(n842) );
  NAND2_X1 U946 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n844), .B(KEYINPUT105), .ZN(n846) );
  NAND2_X1 U948 ( .A1(G136), .A2(n867), .ZN(n845) );
  NAND2_X1 U949 ( .A1(n846), .A2(n845), .ZN(n847) );
  NOR2_X1 U950 ( .A1(n848), .A2(n847), .ZN(G162) );
  XNOR2_X1 U951 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n849), .B(KEYINPUT108), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n864) );
  NAND2_X1 U954 ( .A1(G103), .A2(n869), .ZN(n853) );
  NAND2_X1 U955 ( .A1(G139), .A2(n867), .ZN(n852) );
  NAND2_X1 U956 ( .A1(n853), .A2(n852), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G127), .A2(n873), .ZN(n855) );
  NAND2_X1 U958 ( .A1(G115), .A2(n876), .ZN(n854) );
  NAND2_X1 U959 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U960 ( .A(KEYINPUT47), .B(n856), .Z(n857) );
  NOR2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n922) );
  XOR2_X1 U962 ( .A(n917), .B(n922), .Z(n862) );
  XOR2_X1 U963 ( .A(n860), .B(n859), .Z(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U965 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U966 ( .A(G164), .B(G162), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n882) );
  NAND2_X1 U968 ( .A1(n867), .A2(G142), .ZN(n868) );
  XOR2_X1 U969 ( .A(KEYINPUT107), .B(n868), .Z(n871) );
  NAND2_X1 U970 ( .A1(n869), .A2(G106), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n872), .B(KEYINPUT45), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G130), .A2(n873), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U975 ( .A1(n876), .A2(G118), .ZN(n877) );
  XOR2_X1 U976 ( .A(KEYINPUT106), .B(n877), .Z(n878) );
  NOR2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U978 ( .A(G160), .B(n880), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U980 ( .A1(G37), .A2(n883), .ZN(n884) );
  XOR2_X1 U981 ( .A(KEYINPUT109), .B(n884), .Z(G395) );
  XNOR2_X1 U982 ( .A(n970), .B(n885), .ZN(n887) );
  XNOR2_X1 U983 ( .A(G171), .B(n974), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U985 ( .A(G286), .B(n888), .Z(n889) );
  NOR2_X1 U986 ( .A1(G37), .A2(n889), .ZN(G397) );
  XOR2_X1 U987 ( .A(G1986), .B(G1971), .Z(n891) );
  XNOR2_X1 U988 ( .A(G1966), .B(G1961), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n895) );
  XOR2_X1 U990 ( .A(G1991), .B(G1976), .Z(n893) );
  XNOR2_X1 U991 ( .A(G1996), .B(G1956), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U993 ( .A(n895), .B(n894), .Z(n897) );
  XNOR2_X1 U994 ( .A(G2474), .B(KEYINPUT41), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n899) );
  XOR2_X1 U996 ( .A(G1981), .B(KEYINPUT103), .Z(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(G229) );
  XOR2_X1 U998 ( .A(G2096), .B(KEYINPUT43), .Z(n901) );
  XNOR2_X1 U999 ( .A(G2067), .B(G2678), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1001 ( .A(n902), .B(KEYINPUT42), .Z(n904) );
  XNOR2_X1 U1002 ( .A(G2072), .B(G2090), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U1004 ( .A(KEYINPUT102), .B(G2100), .Z(n906) );
  XNOR2_X1 U1005 ( .A(G2078), .B(G2084), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(G227) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n909), .B(KEYINPUT110), .ZN(n910) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n910), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n911), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n912) );
  XOR2_X1 U1013 ( .A(KEYINPUT49), .B(n912), .Z(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(G225) );
  XNOR2_X1 U1015 ( .A(KEYINPUT111), .B(G225), .ZN(G308) );
  XOR2_X1 U1016 ( .A(G108), .B(KEYINPUT112), .Z(G238) );
  INV_X1 U1018 ( .A(G132), .ZN(G219) );
  INV_X1 U1019 ( .A(G96), .ZN(G221) );
  INV_X1 U1020 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1021 ( .A1(n916), .A2(n915), .ZN(G325) );
  INV_X1 U1022 ( .A(G325), .ZN(G261) );
  INV_X1 U1023 ( .A(G171), .ZN(G301) );
  INV_X1 U1024 ( .A(G57), .ZN(G237) );
  NOR2_X1 U1025 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1026 ( .A(n919), .B(KEYINPUT114), .ZN(n920) );
  NAND2_X1 U1027 ( .A1(n921), .A2(n920), .ZN(n927) );
  XOR2_X1 U1028 ( .A(G2072), .B(n922), .Z(n924) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n923) );
  NOR2_X1 U1030 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n925), .Z(n926) );
  NOR2_X1 U1032 ( .A1(n927), .A2(n926), .ZN(n935) );
  INV_X1 U1033 ( .A(n928), .ZN(n930) );
  NAND2_X1 U1034 ( .A1(n930), .A2(n929), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(G2084), .B(G160), .ZN(n931) );
  XNOR2_X1 U1036 ( .A(KEYINPUT113), .B(n931), .ZN(n932) );
  NOR2_X1 U1037 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1038 ( .A1(n935), .A2(n934), .ZN(n940) );
  XOR2_X1 U1039 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1040 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1041 ( .A(KEYINPUT51), .B(n938), .ZN(n939) );
  NOR2_X1 U1042 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1043 ( .A(KEYINPUT52), .B(n941), .ZN(n943) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n942) );
  NAND2_X1 U1045 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1046 ( .A1(n944), .A2(G29), .ZN(n945) );
  XNOR2_X1 U1047 ( .A(KEYINPUT115), .B(n945), .ZN(n1033) );
  XNOR2_X1 U1048 ( .A(n946), .B(G27), .ZN(n950) );
  XOR2_X1 U1049 ( .A(KEYINPUT118), .B(G32), .Z(n947) );
  XNOR2_X1 U1050 ( .A(n948), .B(n947), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(n951), .B(KEYINPUT119), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(G25), .B(n952), .ZN(n953) );
  NAND2_X1 U1054 ( .A1(n953), .A2(G28), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(G2072), .B(KEYINPUT116), .ZN(n954) );
  XNOR2_X1 U1056 ( .A(n954), .B(G33), .ZN(n956) );
  XNOR2_X1 U1057 ( .A(G26), .B(G2067), .ZN(n955) );
  NOR2_X1 U1058 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1059 ( .A(n957), .B(KEYINPUT117), .ZN(n958) );
  NOR2_X1 U1060 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1062 ( .A(n962), .B(KEYINPUT53), .ZN(n965) );
  XOR2_X1 U1063 ( .A(G2084), .B(G34), .Z(n963) );
  XNOR2_X1 U1064 ( .A(KEYINPUT54), .B(n963), .ZN(n964) );
  NAND2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1066 ( .A(G35), .B(G2090), .ZN(n966) );
  NOR2_X1 U1067 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1068 ( .A(KEYINPUT55), .B(n968), .Z(n969) );
  NOR2_X1 U1069 ( .A1(G29), .A2(n969), .ZN(n1029) );
  INV_X1 U1070 ( .A(G1341), .ZN(n1004) );
  XNOR2_X1 U1071 ( .A(n970), .B(n1004), .ZN(n973) );
  XNOR2_X1 U1072 ( .A(G301), .B(n971), .ZN(n972) );
  NAND2_X1 U1073 ( .A1(n973), .A2(n972), .ZN(n989) );
  XNOR2_X1 U1074 ( .A(G1348), .B(n974), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(n975), .B(G1956), .ZN(n977) );
  NAND2_X1 U1076 ( .A1(G1971), .A2(G303), .ZN(n976) );
  NAND2_X1 U1077 ( .A1(n977), .A2(n976), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1079 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1080 ( .A(KEYINPUT120), .B(n982), .Z(n983) );
  XOR2_X1 U1081 ( .A(KEYINPUT121), .B(n985), .Z(n986) );
  NAND2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(KEYINPUT122), .B(n990), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G168), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(KEYINPUT57), .B(n993), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(G16), .B(KEYINPUT56), .ZN(n996) );
  NAND2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n1027) );
  INV_X1 U1090 ( .A(G16), .ZN(n1025) );
  XNOR2_X1 U1091 ( .A(KEYINPUT123), .B(G1961), .ZN(n998) );
  XNOR2_X1 U1092 ( .A(n998), .B(G5), .ZN(n1014) );
  XNOR2_X1 U1093 ( .A(n999), .B(G20), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(G1981), .B(G6), .Z(n1003) );
  XOR2_X1 U1095 ( .A(G1348), .B(G4), .Z(n1000) );
  XNOR2_X1 U1096 ( .A(KEYINPUT125), .B(n1000), .ZN(n1001) );
  XNOR2_X1 U1097 ( .A(n1001), .B(KEYINPUT59), .ZN(n1002) );
  NAND2_X1 U1098 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  XOR2_X1 U1099 ( .A(KEYINPUT124), .B(n1004), .Z(n1005) );
  XNOR2_X1 U1100 ( .A(G19), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1101 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1102 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1103 ( .A(n1010), .B(KEYINPUT60), .ZN(n1012) );
  XNOR2_X1 U1104 ( .A(G1966), .B(G21), .ZN(n1011) );
  NOR2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1106 ( .A1(n1014), .A2(n1013), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(G1971), .B(G22), .ZN(n1016) );
  XNOR2_X1 U1108 ( .A(G24), .B(G1986), .ZN(n1015) );
  NOR2_X1 U1109 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XOR2_X1 U1110 ( .A(G1976), .B(G23), .Z(n1017) );
  NAND2_X1 U1111 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1112 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1113 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1114 ( .A(n1022), .B(KEYINPUT126), .ZN(n1023) );
  XNOR2_X1 U1115 ( .A(n1023), .B(KEYINPUT61), .ZN(n1024) );
  NAND2_X1 U1116 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1117 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1119 ( .A1(G11), .A2(n1030), .ZN(n1031) );
  XOR2_X1 U1120 ( .A(KEYINPUT127), .B(n1031), .Z(n1032) );
  XNOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1034), .ZN(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

