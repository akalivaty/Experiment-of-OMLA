//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G137), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(KEYINPUT11), .A3(G134), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G134), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n191), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n192), .B(KEYINPUT66), .C1(new_n193), .C2(new_n194), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G131), .Z(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n190), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n192), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n190), .A2(new_n202), .ZN(new_n205));
  OAI21_X1  g019(.A(G131), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n213), .A2(new_n215), .B1(new_n217), .B2(G128), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n212), .B1(new_n209), .B2(new_n211), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  INV_X1    g034(.A(new_n216), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n218), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n207), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT64), .B(G143), .ZN(new_n226));
  OAI211_X1 g040(.A(G128), .B(new_n216), .C1(new_n226), .C2(new_n212), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT0), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n214), .B1(new_n226), .B2(new_n212), .ZN(new_n229));
  XOR2_X1   g043(.A(KEYINPUT0), .B(G128), .Z(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI22_X1  g045(.A1(new_n227), .A2(new_n228), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n195), .A2(new_n196), .ZN(new_n233));
  INV_X1    g047(.A(new_n191), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n198), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n232), .B1(new_n236), .B2(new_n201), .ZN(new_n237));
  XOR2_X1   g051(.A(G116), .B(G119), .Z(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT69), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT2), .B(G113), .Z(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n239), .B(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n225), .A2(new_n237), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n213), .A2(new_n215), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n222), .A2(KEYINPUT0), .B1(new_n245), .B2(new_n230), .ZN(new_n246));
  AND4_X1   g060(.A1(new_n198), .A2(new_n233), .A3(new_n200), .A4(new_n234), .ZN(new_n247));
  INV_X1    g061(.A(G131), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n197), .B2(new_n198), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n246), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n201), .B(new_n206), .C1(new_n251), .C2(new_n218), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n242), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT28), .B1(new_n244), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n242), .A3(new_n252), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT74), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G953), .ZN(new_n262));
  OR2_X1    g076(.A1(KEYINPUT70), .A2(G237), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT70), .A2(G237), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n260), .A2(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G210), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G101), .ZN(new_n267));
  INV_X1    g081(.A(G101), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n268), .A3(G210), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n267), .B2(new_n269), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n255), .A2(new_n274), .A3(new_n256), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n254), .A2(new_n258), .A3(new_n273), .A4(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(G902), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT30), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n225), .B2(new_n237), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n250), .A2(KEYINPUT30), .A3(new_n252), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n243), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n255), .ZN(new_n284));
  INV_X1    g098(.A(new_n273), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n276), .A3(new_n277), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G472), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n254), .A2(new_n258), .A3(new_n275), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n285), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n255), .A2(new_n273), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n255), .A2(KEYINPUT72), .A3(new_n273), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n283), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(KEYINPUT31), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n298), .A2(KEYINPUT31), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n295), .A2(new_n299), .A3(new_n283), .A4(new_n296), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n292), .A2(new_n301), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G472), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n304), .A2(KEYINPUT32), .A3(new_n305), .A4(new_n306), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n311), .A2(new_n310), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n290), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G217), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(G234), .B2(new_n306), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n318));
  AOI21_X1  g132(.A(G902), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n260), .A2(new_n262), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(G221), .A3(G234), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT76), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT22), .B(G137), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT16), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(KEYINPUT16), .B2(new_n328), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(G146), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n220), .A2(G119), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n336), .A2(KEYINPUT23), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(KEYINPUT23), .ZN(new_n338));
  INV_X1    g152(.A(G119), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n337), .A2(new_n338), .B1(new_n339), .B2(G128), .ZN(new_n340));
  INV_X1    g154(.A(G110), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(G128), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT24), .B(G110), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n335), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n334), .A2(new_n212), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n340), .A2(new_n341), .B1(new_n344), .B2(new_n345), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n331), .A2(G146), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n326), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n334), .B(new_n212), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n346), .A3(new_n342), .ZN(new_n355));
  INV_X1    g169(.A(new_n352), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(new_n325), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n320), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n317), .A2(new_n318), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n316), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n360), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n353), .A2(new_n357), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n316), .A2(G902), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n314), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT79), .B(G469), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n371));
  INV_X1    g185(.A(G107), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(G104), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT3), .B1(new_n374), .B2(G107), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n374), .A2(G107), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n268), .B(new_n373), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT4), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G101), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n378), .B(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n219), .A2(new_n221), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n223), .A3(G128), .ZN(new_n383));
  INV_X1    g197(.A(new_n218), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n372), .A2(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(G101), .B1(new_n376), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n377), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n381), .A2(new_n246), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n223), .B1(new_n226), .B2(new_n212), .ZN(new_n392));
  OAI22_X1  g206(.A1(new_n392), .A2(new_n220), .B1(new_n221), .B2(new_n219), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n383), .ZN(new_n394));
  INV_X1    g208(.A(new_n388), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n389), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n236), .A2(new_n201), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n391), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n251), .A2(new_n395), .A3(new_n218), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n388), .B1(new_n393), .B2(new_n383), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n398), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT12), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT12), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n405), .B(new_n398), .C1(new_n401), .C2(new_n402), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n321), .A2(G227), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT78), .ZN(new_n408));
  XNOR2_X1  g222(.A(G110), .B(G140), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n400), .A2(new_n404), .A3(new_n406), .A4(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n378), .A2(G101), .A3(new_n379), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n377), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n246), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n385), .A2(new_n390), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n402), .A2(KEYINPUT10), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n398), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n411), .B1(new_n420), .B2(new_n400), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n306), .B(new_n370), .C1(new_n413), .C2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT80), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n418), .A2(new_n419), .A3(new_n398), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n399), .B1(new_n391), .B2(new_n397), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n410), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(G902), .B1(new_n427), .B2(new_n412), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT80), .A3(new_n370), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n400), .A2(new_n404), .A3(new_n406), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n410), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n420), .A2(new_n400), .A3(new_n411), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n306), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n424), .A2(new_n429), .B1(G469), .B2(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT9), .B(G234), .Z(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G221), .B1(new_n437), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G113), .B(G122), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(new_n374), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n226), .B1(new_n265), .B2(G214), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT70), .B(G237), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n321), .A2(new_n444), .A3(G143), .A4(G214), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n199), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT84), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n321), .A2(new_n444), .A3(G214), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n209), .A2(new_n211), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n445), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT84), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n199), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n200), .A3(new_n445), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n448), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n331), .A2(KEYINPUT19), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n331), .B(KEYINPUT83), .Z(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(KEYINPUT19), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n349), .B1(new_n459), .B2(new_n212), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT18), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n452), .A2(new_n462), .A3(new_n248), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n248), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n451), .B2(new_n445), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n331), .B(KEYINPUT83), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(new_n212), .ZN(new_n467));
  OAI22_X1  g281(.A1(new_n463), .A2(new_n465), .B1(new_n351), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n442), .B1(new_n461), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n468), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n448), .A2(new_n454), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n354), .B1(new_n471), .B2(KEYINPUT17), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT17), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n448), .A2(new_n473), .A3(new_n454), .A4(new_n455), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n470), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n469), .B1(new_n475), .B2(new_n442), .ZN(new_n476));
  OR2_X1    g290(.A1(G475), .A2(G902), .ZN(new_n477));
  OAI211_X1 g291(.A(KEYINPUT85), .B(KEYINPUT20), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n479));
  INV_X1    g293(.A(new_n442), .ZN(new_n480));
  INV_X1    g294(.A(new_n457), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT19), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n212), .B(new_n481), .C1(new_n466), .C2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n212), .B2(new_n334), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n453), .B1(new_n452), .B2(new_n199), .ZN(new_n485));
  AOI211_X1 g299(.A(KEYINPUT84), .B(new_n200), .C1(new_n451), .C2(new_n445), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n484), .B1(new_n487), .B2(new_n455), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n480), .B1(new_n488), .B2(new_n470), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT17), .B1(new_n485), .B2(new_n486), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n474), .A2(new_n490), .A3(new_n335), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n442), .A3(new_n468), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n477), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n479), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n478), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n475), .A2(new_n442), .ZN(new_n498));
  INV_X1    g312(.A(new_n492), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n306), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G475), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n259), .A2(G952), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(G234), .B2(G237), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT21), .B(G898), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n504), .B(KEYINPUT90), .Z(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI211_X1 g320(.A(new_n306), .B(new_n321), .C1(G234), .C2(G237), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n208), .A2(G128), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n189), .B(new_n511), .C1(new_n226), .C2(new_n220), .ZN(new_n512));
  INV_X1    g326(.A(G122), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT86), .B1(new_n513), .B2(G116), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT86), .ZN(new_n515));
  INV_X1    g329(.A(G116), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(G122), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(G116), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n518), .A2(new_n372), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n372), .B1(new_n518), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n512), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g336(.A(KEYINPUT13), .B(new_n511), .C1(new_n226), .C2(new_n220), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n220), .B1(new_n209), .B2(new_n211), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n523), .A2(new_n526), .A3(G134), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT87), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n518), .A2(new_n519), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G107), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n518), .A2(new_n372), .A3(new_n519), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n523), .A2(new_n526), .A3(G134), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n512), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT14), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n514), .A2(new_n517), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n514), .B2(new_n517), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n519), .B(new_n538), .C1(new_n539), .C2(KEYINPUT88), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n539), .A2(KEYINPUT88), .ZN(new_n541));
  OAI21_X1  g355(.A(G107), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G134), .B1(new_n524), .B2(new_n510), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n520), .B1(new_n512), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n542), .A2(KEYINPUT89), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT89), .B1(new_n542), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n536), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n437), .A2(new_n315), .A3(G953), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n536), .B(new_n548), .C1(new_n545), .C2(new_n546), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n306), .ZN(new_n553));
  INV_X1    g367(.A(G478), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(KEYINPUT15), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n553), .B(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n497), .A2(new_n501), .A3(new_n509), .A4(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G214), .B1(G237), .B2(G902), .ZN(new_n559));
  INV_X1    g373(.A(G224), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(G953), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n224), .A2(new_n329), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n232), .A2(G125), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT7), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT5), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n339), .A3(G116), .ZN(new_n568));
  OAI211_X1 g382(.A(G113), .B(new_n568), .C1(new_n238), .C2(new_n567), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n238), .B2(new_n241), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(new_n388), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G122), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  AOI211_X1 g387(.A(new_n565), .B(new_n566), .C1(new_n571), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n243), .A2(new_n381), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n570), .A2(new_n388), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n572), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n563), .A2(KEYINPUT7), .A3(new_n562), .A4(new_n564), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n563), .A2(new_n564), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(new_n561), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n572), .B(KEYINPUT81), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n575), .B2(new_n576), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n584), .A2(KEYINPUT6), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n577), .B1(new_n584), .B2(KEYINPUT6), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G210), .B1(G237), .B2(G902), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n580), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n588), .B(KEYINPUT82), .Z(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n580), .B2(new_n587), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n559), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n440), .A2(new_n558), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n369), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  NAND2_X1  g410(.A1(new_n497), .A2(new_n501), .ZN(new_n597));
  AOI21_X1  g411(.A(G478), .B1(new_n552), .B2(new_n306), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n550), .A2(KEYINPUT91), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n552), .A2(new_n599), .A3(KEYINPUT33), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n550), .B(new_n551), .C1(KEYINPUT91), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n554), .A2(G902), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n598), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n559), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n580), .A2(new_n587), .ZN(new_n608));
  INV_X1    g422(.A(new_n588), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n607), .B1(new_n610), .B2(new_n589), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n597), .A2(new_n509), .A3(new_n606), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT92), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n605), .B1(new_n497), .B2(new_n501), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT92), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n614), .A2(new_n615), .A3(new_n509), .A4(new_n611), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n304), .A2(new_n306), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(G472), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n619), .A2(new_n307), .ZN(new_n620));
  INV_X1    g434(.A(new_n363), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n367), .B(new_n438), .C1(new_n621), .C2(new_n361), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n424), .A2(new_n429), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n434), .A2(G469), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n617), .A2(new_n620), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NAND4_X1  g442(.A1(new_n625), .A2(new_n307), .A3(new_n509), .A4(new_n619), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n553), .B(new_n555), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n497), .A2(new_n630), .A3(new_n501), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n611), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT35), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NAND2_X1  g452(.A1(new_n355), .A2(new_n356), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n325), .A2(KEYINPUT36), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n366), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n364), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n619), .A2(new_n643), .A3(new_n307), .ZN(new_n644));
  INV_X1    g458(.A(new_n558), .ZN(new_n645));
  INV_X1    g459(.A(new_n593), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n435), .A2(new_n439), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n644), .A2(new_n645), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT37), .B(G110), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n651));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n503), .B1(new_n507), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n631), .A2(new_n651), .A3(new_n611), .A4(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n497), .A2(new_n501), .A3(new_n630), .A4(new_n654), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT95), .B1(new_n656), .B2(new_n633), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n643), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n312), .A2(new_n313), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n659), .B1(new_n660), .B2(new_n289), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n658), .A2(new_n661), .A3(new_n647), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  NOR2_X1   g477(.A1(new_n590), .A2(new_n592), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT38), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n665), .A2(new_n607), .A3(new_n643), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n557), .B1(new_n497), .B2(new_n501), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n653), .B(KEYINPUT39), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n647), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n668), .B1(KEYINPUT40), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n285), .B1(new_n244), .B2(new_n253), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n297), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n674), .B2(G902), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n660), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n672), .B(new_n676), .C1(KEYINPUT40), .C2(new_n671), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n226), .ZN(G45));
  AND3_X1   g492(.A1(new_n614), .A2(KEYINPUT96), .A3(new_n654), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT96), .B1(new_n614), .B2(new_n654), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n661), .A2(new_n681), .A3(new_n647), .A4(new_n611), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT97), .B(G146), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G48));
  NAND2_X1  g498(.A1(new_n660), .A2(new_n289), .ZN(new_n685));
  INV_X1    g499(.A(new_n368), .ZN(new_n686));
  INV_X1    g500(.A(G469), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n428), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n422), .A2(new_n423), .ZN(new_n689));
  AOI21_X1  g503(.A(KEYINPUT80), .B1(new_n428), .B2(new_n370), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n438), .B(new_n688), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT98), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT98), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n623), .A2(new_n693), .A3(new_n438), .A4(new_n688), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n617), .A2(new_n685), .A3(new_n686), .A4(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT41), .B(G113), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT99), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n697), .B(new_n699), .ZN(G15));
  NOR2_X1   g514(.A1(new_n695), .A2(new_n633), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n632), .A2(new_n508), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n685), .A2(new_n701), .A3(new_n686), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  NAND4_X1  g518(.A1(new_n685), .A2(new_n701), .A3(new_n645), .A4(new_n643), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  NOR2_X1   g520(.A1(G472), .A2(G902), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT100), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n304), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT101), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n304), .A2(KEYINPUT101), .A3(new_n708), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n619), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n368), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n667), .A2(new_n611), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n696), .A2(new_n714), .A3(new_n509), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  NAND4_X1  g531(.A1(new_n619), .A2(new_n711), .A3(new_n643), .A4(new_n712), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n681), .A2(new_n701), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  NAND3_X1  g535(.A1(new_n309), .A2(new_n289), .A3(new_n311), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n432), .A2(KEYINPUT103), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n420), .A2(new_n400), .A3(new_n724), .A4(new_n411), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT102), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n431), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n430), .A2(KEYINPUT102), .A3(new_n410), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(G469), .B1(new_n730), .B2(G902), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n439), .B1(new_n731), .B2(new_n623), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n722), .A2(new_n732), .A3(new_n686), .ZN(new_n733));
  INV_X1    g547(.A(new_n680), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n614), .A2(KEYINPUT96), .A3(new_n654), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n664), .A2(new_n559), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n733), .A2(new_n734), .A3(new_n735), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n732), .A2(new_n737), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n314), .A2(new_n368), .A3(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT42), .ZN(new_n741));
  AOI22_X1  g555(.A1(KEYINPUT42), .A2(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  INV_X1    g557(.A(new_n739), .ZN(new_n744));
  INV_X1    g558(.A(new_n656), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n685), .A2(new_n744), .A3(new_n686), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  NAND2_X1  g561(.A1(new_n730), .A2(KEYINPUT45), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n687), .B1(new_n433), .B2(new_n749), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n748), .A2(new_n750), .B1(G469), .B2(G902), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(KEYINPUT46), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n751), .A2(KEYINPUT46), .B1(new_n424), .B2(new_n429), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n439), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n670), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT104), .Z(new_n757));
  INV_X1    g571(.A(new_n597), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n606), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT43), .B1(new_n759), .B2(KEYINPUT105), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n761), .A2(new_n762), .A3(new_n620), .A4(new_n659), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n757), .B1(KEYINPUT44), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(KEYINPUT44), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n736), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT106), .B(G137), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G39));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n755), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n755), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n314), .A2(new_n681), .A3(new_n368), .A4(new_n737), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT108), .B(G140), .Z(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G42));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n665), .A2(new_n686), .A3(new_n559), .A4(new_n438), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n623), .A2(new_n688), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(KEYINPUT49), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(KEYINPUT49), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n676), .ZN(new_n789));
  INV_X1    g603(.A(new_n759), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT109), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n685), .A2(new_n686), .A3(new_n594), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n620), .A2(new_n509), .A3(new_n646), .A4(new_n625), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n631), .A2(new_n614), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n648), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n792), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n629), .A2(new_n593), .ZN(new_n798));
  INV_X1    g612(.A(new_n795), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n595), .A2(KEYINPUT109), .A3(new_n648), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n497), .A2(new_n501), .A3(new_n557), .A4(new_n654), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT110), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n737), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n803), .A2(KEYINPUT110), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n661), .A2(new_n807), .A3(new_n647), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n744), .A2(new_n734), .A3(new_n719), .A4(new_n735), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n746), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT111), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n697), .A2(new_n703), .A3(new_n705), .A4(new_n716), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n802), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n808), .A2(new_n746), .A3(new_n814), .A4(new_n809), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n742), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n653), .B(KEYINPUT112), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n732), .A2(new_n659), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n676), .A2(new_n715), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n682), .A2(new_n662), .A3(new_n720), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n314), .A2(new_n440), .A3(new_n659), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n679), .A2(new_n680), .A3(new_n718), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n824), .A2(new_n658), .B1(new_n825), .B2(new_n701), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(KEYINPUT52), .A3(new_n682), .A4(new_n820), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(new_n827), .A3(KEYINPUT113), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n821), .A2(new_n829), .A3(new_n822), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n817), .A2(KEYINPUT53), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n697), .A2(new_n703), .A3(new_n705), .A4(new_n716), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n797), .B2(new_n801), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n815), .A2(new_n742), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n836), .A3(new_n811), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n823), .A2(new_n827), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n831), .A2(new_n832), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n835), .A2(new_n836), .A3(new_n830), .A4(new_n811), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n823), .A2(KEYINPUT113), .A3(new_n827), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n833), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(KEYINPUT114), .B(new_n833), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n837), .A2(new_n838), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n840), .B1(new_n849), .B2(KEYINPUT54), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  INV_X1    g665(.A(new_n762), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n503), .A3(new_n714), .A4(new_n760), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n695), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n665), .A2(new_n607), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT50), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n856), .B(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n695), .A2(new_n736), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n789), .A2(new_n686), .A3(new_n503), .A4(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n597), .A3(new_n606), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n852), .A2(new_n503), .A3(new_n760), .A4(new_n859), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n861), .B1(new_n866), .B2(new_n719), .ZN(new_n867));
  INV_X1    g681(.A(new_n853), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n737), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n777), .A2(KEYINPUT115), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n785), .A2(new_n438), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n777), .B2(KEYINPUT115), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT116), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n858), .B(new_n867), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n851), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n614), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n860), .A2(new_n878), .ZN(new_n879));
  AOI211_X1 g693(.A(new_n502), .B(new_n879), .C1(new_n611), .C2(new_n854), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT48), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n722), .A2(new_n686), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n881), .B1(new_n866), .B2(new_n883), .ZN(new_n884));
  AOI211_X1 g698(.A(KEYINPUT48), .B(new_n882), .C1(new_n864), .C2(new_n865), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n858), .A2(new_n867), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n777), .B1(new_n438), .B2(new_n785), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n869), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n851), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n886), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n877), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n850), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(G952), .A2(G953), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n783), .B(new_n791), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n896), .B1(new_n850), .B2(new_n894), .ZN(new_n898));
  INV_X1    g712(.A(new_n791), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT119), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(G75));
  NOR2_X1   g715(.A1(new_n585), .A2(new_n586), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n582), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n831), .A2(new_n839), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(G902), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(G210), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n321), .A2(G952), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n906), .A2(new_n591), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n904), .A2(new_n909), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n910), .A2(new_n915), .ZN(G51));
  NAND2_X1  g730(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n831), .A2(new_n832), .A3(new_n839), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(G469), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT57), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n421), .B2(new_n413), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n907), .A2(new_n748), .A3(new_n750), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n911), .B1(new_n923), .B2(new_n924), .ZN(G54));
  NAND3_X1  g739(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n926), .A2(new_n476), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n476), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n927), .A2(new_n928), .A3(new_n911), .ZN(G60));
  INV_X1    g743(.A(new_n603), .ZN(new_n930));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n850), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n930), .A2(new_n932), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n911), .B1(new_n919), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n933), .A2(new_n935), .A3(KEYINPUT120), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT121), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n365), .B1(new_n905), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n905), .A2(new_n641), .A3(new_n943), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n912), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  OAI22_X1  g761(.A1(new_n944), .A2(new_n946), .B1(KEYINPUT122), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G66));
  INV_X1    g764(.A(new_n835), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n321), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n259), .B1(new_n505), .B2(G224), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT124), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n902), .B1(G898), .B2(new_n321), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G69));
  NAND2_X1  g774(.A1(new_n281), .A2(new_n282), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(new_n459), .Z(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(G227), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n963), .A2(new_n652), .A3(new_n321), .ZN(new_n964));
  AOI22_X1  g778(.A1(new_n764), .A2(new_n766), .B1(new_n778), .B2(new_n779), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n826), .A2(new_n682), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n883), .A2(new_n715), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n746), .B1(new_n757), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n742), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n965), .A2(new_n966), .A3(new_n970), .ZN(new_n971));
  AOI22_X1  g785(.A1(new_n971), .A2(new_n962), .B1(new_n260), .B2(new_n262), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n677), .A2(new_n966), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT62), .Z(new_n974));
  NOR3_X1   g788(.A1(new_n795), .A2(new_n671), .A3(new_n736), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n369), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n976), .A3(new_n965), .ZN(new_n977));
  INV_X1    g791(.A(new_n962), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n964), .B1(new_n972), .B2(new_n979), .ZN(G72));
  NOR2_X1   g794(.A1(new_n284), .A2(new_n273), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT127), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n965), .A2(new_n966), .A3(new_n970), .A4(new_n835), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT126), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT63), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT125), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n983), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n984), .B1(new_n983), .B2(new_n987), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n987), .B1(new_n977), .B2(new_n951), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n285), .B1(new_n283), .B2(new_n255), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n911), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n986), .B1(new_n286), .B2(new_n297), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n849), .B2(new_n995), .ZN(G57));
endmodule


