//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n209), .A2(KEYINPUT0), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(KEYINPUT0), .B2(new_n209), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT66), .B(G77), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n222), .A2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G58), .A2(G232), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT67), .Z(new_n231));
  AOI211_X1 g0031(.A(new_n220), .B(new_n231), .C1(KEYINPUT1), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND2_X1  g0048(.A1(new_n214), .A2(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n211), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  INV_X1    g0051(.A(G50), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n211), .A2(new_n253), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n249), .B1(new_n250), .B2(new_n251), .C1(new_n252), .C2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(new_n206), .B2(new_n253), .ZN(new_n257));
  NAND4_X1  g0057(.A1(KEYINPUT68), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(new_n210), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g0060(.A(new_n260), .B(KEYINPUT11), .Z(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n214), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT12), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n211), .A2(G1), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n266), .B1(new_n269), .B2(new_n214), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G238), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  OAI211_X1 g0078(.A(G1), .B(G13), .C1(new_n253), .C2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n275), .A2(new_n279), .A3(G274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n234), .A2(G1698), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n282), .B(new_n283), .C1(G226), .C2(G1698), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G97), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n279), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OR3_X1    g0086(.A1(new_n281), .A2(new_n286), .A3(KEYINPUT13), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT13), .B1(new_n281), .B2(new_n286), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT14), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n290), .A3(G169), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n287), .A2(G179), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n290), .B1(new_n289), .B2(G169), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n272), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(G200), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n296), .B(new_n271), .C1(new_n297), .C2(new_n289), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(KEYINPUT71), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n213), .A2(KEYINPUT8), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT8), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G58), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n254), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT15), .B(G87), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n306), .B1(new_n211), .B2(new_n221), .C1(new_n250), .C2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n308), .A2(new_n259), .B1(new_n221), .B2(new_n264), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n268), .A2(G77), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G1698), .ZN(new_n312));
  OR2_X1    g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(KEYINPUT3), .A2(G33), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n315), .A2(G238), .B1(new_n318), .B2(G107), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n282), .A2(G232), .A3(new_n312), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n273), .ZN(new_n322));
  INV_X1    g0122(.A(new_n280), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(G244), .B2(new_n276), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n311), .B1(G190), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n326), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n325), .A2(new_n332), .B1(new_n309), .B2(new_n310), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n299), .B2(KEYINPUT71), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT75), .ZN(new_n337));
  OAI211_X1 g0137(.A(G226), .B(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT73), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT73), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n282), .A2(new_n340), .A3(G226), .A4(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G87), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n282), .A2(G223), .A3(new_n312), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n339), .A2(new_n341), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n273), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n279), .A2(G232), .A3(new_n274), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n280), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(G200), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  AOI211_X1 g0149(.A(G190), .B(new_n347), .C1(new_n344), .C2(new_n273), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n337), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n345), .A2(new_n297), .A3(new_n348), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n347), .B1(new_n344), .B2(new_n273), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n352), .B(KEYINPUT75), .C1(G200), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT72), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G58), .A2(G68), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n211), .B1(new_n215), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G159), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n254), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(G58), .A2(G68), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n363), .B2(new_n202), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(KEYINPUT72), .C1(new_n360), .C2(new_n254), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n282), .B2(G20), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n318), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n214), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n356), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT7), .B1(new_n318), .B2(new_n211), .ZN(new_n372));
  NOR4_X1   g0172(.A1(new_n316), .A2(new_n317), .A3(new_n367), .A4(G20), .ZN(new_n373));
  OAI21_X1  g0173(.A(G68), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n374), .A2(KEYINPUT16), .A3(new_n362), .A4(new_n365), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n371), .A2(new_n375), .A3(new_n259), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT69), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n301), .A2(new_n303), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT70), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n302), .A2(KEYINPUT69), .A3(G58), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n379), .B1(new_n378), .B2(new_n380), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n264), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n383), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(new_n268), .A3(new_n381), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n376), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  XOR2_X1   g0189(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n390));
  NAND3_X1  g0190(.A1(new_n355), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  OR2_X1    g0191(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n351), .B2(new_n354), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n353), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n332), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n353), .A2(KEYINPUT74), .A3(new_n330), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT74), .B1(new_n353), .B2(new_n330), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT18), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n399), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n353), .A2(KEYINPUT74), .A3(new_n330), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n376), .A2(new_n387), .B1(new_n332), .B2(new_n395), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n394), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n323), .B1(G226), .B2(new_n276), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n222), .A2(new_n318), .B1(new_n315), .B2(G223), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n282), .A2(G222), .A3(new_n312), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n410), .B1(new_n413), .B2(new_n279), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n332), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(G179), .B2(new_n414), .ZN(new_n416));
  INV_X1    g0216(.A(new_n259), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n382), .A2(new_n383), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(new_n211), .A3(G33), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n305), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n264), .A2(new_n252), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n269), .B2(new_n252), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n414), .A2(new_n297), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(G200), .B2(new_n414), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT9), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n421), .A2(KEYINPUT9), .A3(new_n423), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT10), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT10), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n433), .B(new_n427), .C1(new_n429), .C2(new_n430), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n425), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n300), .A2(new_n336), .A3(new_n409), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT21), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n282), .A2(G264), .A3(G1698), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n282), .A2(G257), .A3(new_n312), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n318), .A2(G303), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT81), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT81), .A4(new_n441), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n273), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT5), .B(G41), .ZN(new_n447));
  INV_X1    g0247(.A(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G1), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n447), .A2(new_n279), .A3(G274), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n449), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n279), .ZN(new_n452));
  INV_X1    g0252(.A(G270), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n446), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G169), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT82), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT79), .B(G116), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n458), .B1(new_n460), .B2(new_n263), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n264), .A3(KEYINPUT82), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n263), .B1(G1), .B2(new_n253), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n259), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G116), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n470), .B(new_n211), .C1(G33), .C2(new_n471), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT83), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n459), .A2(G20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n259), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n469), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT83), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n472), .B(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n478), .A2(KEYINPUT20), .A3(new_n259), .A4(new_n474), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n468), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n438), .B1(new_n457), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n279), .B1(new_n442), .B2(new_n443), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n454), .B1(new_n482), .B2(new_n445), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G190), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n484), .B(new_n480), .C1(new_n328), .C2(new_n483), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n476), .A2(new_n479), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n465), .A2(G116), .B1(new_n461), .B2(new_n462), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(G179), .A3(new_n483), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n488), .A2(new_n456), .A3(KEYINPUT21), .A4(G169), .ZN(new_n490));
  AND4_X1   g0290(.A1(new_n481), .A2(new_n485), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G257), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n450), .B1(new_n452), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(G244), .B(new_n312), .C1(new_n316), .C2(new_n317), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT77), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n315), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n493), .B1(new_n501), .B2(new_n273), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n332), .ZN(new_n503));
  AOI211_X1 g0303(.A(new_n330), .B(new_n493), .C1(new_n501), .C2(new_n273), .ZN(new_n504));
  OAI21_X1  g0304(.A(G107), .B1(new_n372), .B2(new_n373), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT6), .ZN(new_n506));
  AND2_X1   g0306(.A1(G97), .A2(G107), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G107), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(KEYINPUT6), .A3(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n512), .A2(G20), .B1(G77), .B2(new_n305), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n417), .B1(new_n505), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n464), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n258), .A2(new_n210), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(G97), .A4(new_n257), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(G97), .B2(new_n263), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n514), .A2(KEYINPUT78), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT78), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n305), .A2(G77), .ZN(new_n521));
  INV_X1    g0321(.A(new_n511), .ZN(new_n522));
  XNOR2_X1  g0322(.A(G97), .B(G107), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(new_n506), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n521), .B1(new_n524), .B2(new_n211), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n510), .B1(new_n368), .B2(new_n369), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n259), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n263), .A2(G97), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n465), .B2(G97), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n520), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n503), .A2(new_n504), .B1(new_n519), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n529), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n502), .A2(G190), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n534), .C1(new_n328), .C2(new_n502), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(G238), .B(new_n312), .C1(new_n316), .C2(new_n317), .ZN(new_n537));
  OAI211_X1 g0337(.A(G244), .B(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n538), .C1(new_n253), .C2(new_n459), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n273), .ZN(new_n540));
  INV_X1    g0340(.A(new_n449), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n279), .A2(new_n541), .A3(G250), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n279), .A2(G274), .A3(new_n449), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n540), .A2(new_n297), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n544), .B1(new_n273), .B2(new_n539), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(G200), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n307), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n263), .ZN(new_n550));
  INV_X1    g0350(.A(G87), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n259), .A2(new_n551), .A3(new_n464), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n282), .A2(new_n211), .A3(G68), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n250), .B2(new_n471), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n211), .B1(new_n285), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n508), .A2(new_n551), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n556), .A2(KEYINPUT80), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT80), .B1(new_n556), .B2(new_n557), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n553), .B(new_n555), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  AOI211_X1 g0360(.A(new_n550), .B(new_n552), .C1(new_n560), .C2(new_n259), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n548), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n259), .ZN(new_n563));
  INV_X1    g0363(.A(new_n550), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n465), .A2(new_n549), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n547), .A2(new_n330), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n540), .A2(new_n545), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n332), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n282), .A2(G257), .A3(G1698), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n282), .A2(G250), .A3(new_n312), .ZN(new_n573));
  INV_X1    g0373(.A(G294), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n572), .B(new_n573), .C1(new_n253), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n273), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n451), .A2(G264), .A3(new_n279), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(new_n330), .A3(new_n450), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n450), .A3(new_n577), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n332), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n211), .B(G87), .C1(new_n316), .C2(new_n317), .ZN(new_n582));
  XNOR2_X1  g0382(.A(new_n582), .B(KEYINPUT22), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n459), .A2(new_n253), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT23), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n211), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n510), .A2(KEYINPUT23), .A3(G20), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n584), .A2(new_n211), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT24), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT24), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n583), .A2(new_n591), .A3(new_n588), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n417), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT25), .ZN(new_n595));
  AOI211_X1 g0395(.A(G107), .B(new_n263), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  OR2_X1    g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n598), .A2(new_n599), .B1(G107), .B2(new_n465), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n579), .B(new_n581), .C1(new_n593), .C2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n578), .A2(G190), .A3(new_n450), .ZN(new_n603));
  INV_X1    g0403(.A(new_n592), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n591), .B1(new_n583), .B2(new_n588), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n259), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n580), .A2(G200), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n603), .A2(new_n606), .A3(new_n600), .A4(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n571), .A2(new_n602), .A3(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n437), .A2(new_n491), .A3(new_n536), .A4(new_n609), .ZN(G372));
  AND2_X1   g0410(.A1(new_n490), .A2(new_n489), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(new_n481), .A3(new_n602), .ZN(new_n612));
  AOI21_X1  g0412(.A(G169), .B1(new_n540), .B2(new_n545), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n613), .A2(KEYINPUT85), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(KEYINPUT85), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n614), .A2(new_n566), .A3(new_n567), .A4(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n608), .A2(new_n616), .A3(new_n562), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n612), .A2(new_n617), .A3(new_n536), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n501), .A2(new_n273), .ZN(new_n619));
  INV_X1    g0419(.A(new_n493), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G169), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n502), .A2(G179), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n532), .A2(KEYINPUT78), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n527), .A2(new_n520), .A3(new_n529), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n624), .A2(new_n627), .A3(new_n570), .A4(new_n562), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT26), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n533), .B1(new_n622), .B2(new_n623), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(new_n616), .A4(new_n562), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n629), .A2(new_n632), .A3(new_n616), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n436), .B1(new_n618), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n298), .A2(new_n331), .A3(new_n333), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n295), .ZN(new_n636));
  INV_X1    g0436(.A(new_n390), .ZN(new_n637));
  AOI211_X1 g0437(.A(new_n637), .B(new_n388), .C1(new_n351), .C2(new_n354), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n392), .B1(new_n355), .B2(new_n389), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n408), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n432), .A2(new_n434), .ZN(new_n642));
  OAI22_X1  g0442(.A1(new_n641), .A2(new_n642), .B1(new_n424), .B2(new_n416), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n634), .A2(new_n643), .ZN(G369));
  NAND2_X1  g0444(.A1(new_n611), .A2(new_n481), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n262), .A2(new_n211), .A3(G13), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G343), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n488), .A2(new_n651), .ZN(new_n652));
  MUX2_X1   g0452(.A(new_n645), .B(new_n491), .S(new_n652), .Z(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G330), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n602), .A2(new_n651), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n651), .B1(new_n593), .B2(new_n601), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n608), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n657), .B1(new_n602), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n651), .B1(new_n611), .B2(new_n481), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n657), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n207), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n557), .A2(G116), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G1), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n216), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n651), .B1(new_n633), .B2(new_n618), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT29), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n612), .A2(new_n617), .A3(new_n536), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT87), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n562), .A2(new_n570), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n676), .B(new_n631), .C1(new_n531), .C2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n630), .A2(new_n616), .A3(KEYINPUT26), .A4(new_n562), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n676), .B1(new_n628), .B2(new_n631), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n616), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT88), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n675), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI211_X1 g0484(.A(KEYINPUT88), .B(new_n616), .C1(new_n680), .C2(new_n681), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n651), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n674), .B1(new_n686), .B2(new_n673), .ZN(new_n687));
  INV_X1    g0487(.A(new_n651), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n491), .A2(new_n609), .A3(new_n536), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT31), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n483), .A2(G179), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n547), .A2(new_n577), .A3(new_n576), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(KEYINPUT30), .A3(new_n502), .A4(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n502), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n691), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n547), .A2(G179), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n456), .A2(new_n621), .A3(new_n580), .A4(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT86), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n700), .B(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n688), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n690), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n700), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n687), .B1(G330), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n671), .B1(new_n709), .B2(G1), .ZN(G364));
  AND2_X1   g0510(.A1(new_n211), .A2(G13), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n262), .B1(new_n711), .B2(G45), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n666), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n656), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(G330), .B2(new_n653), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G13), .A2(G33), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n654), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n211), .A2(new_n330), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n328), .A2(G190), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G317), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT33), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n725), .A2(KEYINPUT33), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G311), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n330), .A2(G200), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(G20), .A3(new_n297), .ZN(new_n731));
  INV_X1    g0531(.A(G322), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(G20), .A3(G190), .ZN(new_n733));
  OAI221_X1 g0533(.A(new_n728), .B1(new_n729), .B2(new_n731), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n297), .A2(new_n328), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(G20), .A3(new_n330), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n282), .B(new_n734), .C1(G303), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n330), .A2(new_n328), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT91), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n740), .A2(new_n211), .A3(G190), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT90), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n735), .A2(new_n721), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n742), .B1(new_n735), .B2(new_n721), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(G329), .A2(new_n741), .B1(new_n746), .B2(G326), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n738), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G283), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n722), .A2(G20), .A3(new_n330), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT93), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT94), .Z(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(G20), .B1(new_n740), .B2(new_n297), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n748), .B1(new_n749), .B2(new_n756), .C1(new_n574), .C2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n741), .ZN(new_n760));
  OR3_X1    g0560(.A1(new_n760), .A2(KEYINPUT32), .A3(new_n360), .ZN(new_n761));
  OAI21_X1  g0561(.A(KEYINPUT32), .B1(new_n760), .B2(new_n360), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n757), .A2(G97), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n755), .A2(G107), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n213), .A2(new_n733), .B1(new_n723), .B2(new_n214), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n318), .B1(new_n737), .B2(G87), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(KEYINPUT92), .ZN(new_n768));
  INV_X1    g0568(.A(new_n731), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n766), .B(new_n768), .C1(new_n222), .C2(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n746), .A2(G50), .B1(new_n767), .B2(KEYINPUT92), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n765), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n759), .B1(new_n764), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n210), .B1(G20), .B2(new_n332), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n318), .A2(new_n207), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n448), .B2(new_n217), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n247), .B2(new_n448), .ZN(new_n778));
  INV_X1    g0578(.A(G355), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n665), .A2(new_n318), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT89), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n778), .B1(G116), .B2(new_n207), .C1(new_n779), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n719), .A2(new_n774), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n720), .A2(new_n714), .A3(new_n775), .A4(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n716), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(G396));
  INV_X1    g0587(.A(new_n774), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n756), .A2(new_n214), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT34), .ZN(new_n790));
  INV_X1    g0590(.A(new_n733), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n791), .A2(G143), .B1(new_n769), .B2(G159), .ZN(new_n792));
  INV_X1    g0592(.A(G150), .ZN(new_n793));
  INV_X1    g0593(.A(G137), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n792), .B1(new_n793), .B2(new_n723), .C1(new_n745), .C2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n789), .B1(new_n790), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G132), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n282), .B1(new_n252), .B2(new_n736), .C1(new_n760), .C2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n757), .B2(G58), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n796), .B(new_n799), .C1(new_n790), .C2(new_n795), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n755), .A2(G87), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n318), .B1(new_n723), .B2(new_n749), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n736), .A2(new_n510), .B1(new_n731), .B2(new_n459), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(G294), .C2(new_n791), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G311), .A2(new_n741), .B1(new_n746), .B2(G303), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n801), .A2(new_n763), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n800), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n788), .B1(new_n807), .B2(KEYINPUT95), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(KEYINPUT95), .B2(new_n807), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n774), .A2(new_n717), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n809), .B(new_n714), .C1(G77), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n334), .A2(new_n651), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n311), .A2(new_n651), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n329), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n813), .B1(new_n815), .B2(new_n334), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n812), .B1(new_n717), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n672), .B(new_n816), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n708), .A2(G330), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n714), .B1(new_n819), .B2(new_n820), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G384));
  OR2_X1    g0624(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n825), .A2(new_n826), .A3(G116), .A4(new_n212), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT36), .Z(new_n828));
  NAND3_X1  g0628(.A1(new_n217), .A2(new_n222), .A3(new_n358), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n201), .A2(G68), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n262), .B(G13), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n295), .A2(new_n651), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  INV_X1    g0635(.A(new_n649), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n388), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n397), .A2(new_n400), .A3(KEYINPUT18), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n406), .B1(new_n404), .B2(new_n405), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n837), .B1(new_n640), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n404), .A2(new_n405), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n837), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n842), .B1(new_n844), .B2(new_n393), .ZN(new_n845));
  INV_X1    g0645(.A(new_n393), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n846), .A2(KEYINPUT37), .A3(new_n843), .A4(new_n837), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n835), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT97), .ZN(new_n850));
  INV_X1    g0650(.A(new_n837), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n394), .B2(new_n408), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT96), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n842), .B1(new_n837), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n844), .B2(new_n393), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n846), .A2(new_n854), .A3(new_n843), .A4(new_n837), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n852), .A2(KEYINPUT38), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT39), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n849), .A2(new_n850), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n849), .A2(new_n859), .A3(new_n858), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT97), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n856), .A2(new_n857), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n835), .B1(new_n841), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n859), .B1(new_n864), .B2(new_n858), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n834), .B(new_n860), .C1(new_n862), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n272), .A2(new_n651), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n295), .A2(new_n298), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(new_n295), .B2(new_n298), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n672), .A2(new_n816), .ZN(new_n871));
  INV_X1    g0671(.A(new_n813), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n864), .A2(new_n858), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n873), .A2(new_n874), .B1(new_n408), .B2(new_n649), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n866), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n643), .B1(new_n687), .B2(new_n437), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n876), .B(new_n877), .Z(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n816), .B1(new_n868), .B2(new_n869), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n703), .A2(KEYINPUT31), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(new_n705), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n849), .A2(new_n858), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(new_n874), .A3(new_n879), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n703), .B1(new_n689), .B2(KEYINPUT31), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n703), .A2(KEYINPUT31), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n436), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n655), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n891), .B2(new_n887), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n878), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n262), .B2(new_n711), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n878), .A2(new_n893), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n832), .B1(new_n895), .B2(new_n896), .ZN(G367));
  OAI221_X1 g0697(.A(new_n783), .B1(new_n207), .B2(new_n307), .C1(new_n240), .C2(new_n776), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n714), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n758), .A2(new_n214), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(G150), .B2(new_n791), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT101), .Z(new_n902));
  OAI22_X1  g0702(.A1(new_n201), .A2(new_n731), .B1(new_n723), .B2(new_n360), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n318), .B(new_n903), .C1(G58), .C2(new_n737), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n741), .A2(G137), .ZN(new_n905));
  INV_X1    g0705(.A(new_n754), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n222), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n746), .A2(G143), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n904), .A2(new_n905), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT46), .B1(new_n736), .B2(new_n467), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n459), .A2(KEYINPUT46), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(new_n736), .B2(new_n911), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n912), .B1(new_n729), .B2(new_n745), .C1(new_n760), .C2(new_n725), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n731), .A2(new_n749), .B1(new_n723), .B2(new_n574), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n282), .B(new_n914), .C1(G303), .C2(new_n791), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n915), .B1(new_n471), .B2(new_n754), .C1(new_n510), .C2(new_n758), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n902), .A2(new_n909), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT47), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n899), .B1(new_n918), .B2(new_n774), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n561), .A2(new_n688), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n616), .B2(new_n562), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n616), .B2(new_n920), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT98), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n719), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n709), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n531), .B(new_n535), .C1(new_n533), .C2(new_n688), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT99), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n630), .A2(new_n651), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n663), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT45), .Z(new_n932));
  NOR2_X1   g0732(.A1(new_n930), .A2(new_n663), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT44), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n661), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n661), .B1(new_n932), .B2(new_n934), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n660), .B(new_n662), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n656), .B(new_n939), .Z(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n926), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n666), .B(KEYINPUT41), .Z(new_n943));
  OAI21_X1  g0743(.A(new_n712), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n930), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n661), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT100), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n923), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT100), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n947), .B(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n950), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n946), .A2(new_n602), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n651), .B1(new_n957), .B2(new_n531), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n930), .A2(new_n660), .A3(new_n662), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT42), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n923), .A2(new_n949), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n951), .A2(new_n955), .A3(new_n963), .A4(new_n961), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n925), .B1(new_n945), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT102), .ZN(new_n969));
  INV_X1    g0769(.A(new_n967), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n944), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT102), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n972), .A3(new_n925), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n969), .A2(new_n973), .ZN(G387));
  NAND2_X1  g0774(.A1(new_n926), .A2(new_n940), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n709), .A2(new_n941), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n976), .A3(new_n666), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n781), .A2(new_n668), .B1(G107), .B2(new_n207), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n237), .A2(new_n448), .ZN(new_n979));
  INV_X1    g0779(.A(new_n668), .ZN(new_n980));
  AOI211_X1 g0780(.A(G45), .B(new_n980), .C1(G68), .C2(G77), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n304), .A2(new_n252), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT50), .Z(new_n983));
  AOI21_X1  g0783(.A(new_n776), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n978), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT103), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n783), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n714), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n282), .B1(new_n736), .B2(new_n221), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT104), .B(G150), .Z(new_n991));
  AOI21_X1  g0791(.A(new_n990), .B1(new_n741), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n756), .B2(new_n471), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT105), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n757), .A2(new_n549), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n791), .A2(G50), .B1(new_n769), .B2(G68), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(new_n360), .C2(new_n745), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n418), .B2(new_n724), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(G303), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n731), .A2(new_n1000), .B1(new_n733), .B2(new_n725), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT106), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n729), .B2(new_n723), .C1(new_n732), .C2(new_n745), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT48), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT107), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n757), .A2(G283), .B1(G294), .B2(new_n737), .ZN(new_n1008));
  AND3_X1   g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1007), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1005), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT108), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT108), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1013), .B(new_n1005), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(KEYINPUT49), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n318), .B1(new_n754), .B2(new_n459), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G326), .B2(new_n741), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT49), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n999), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n989), .B1(new_n1020), .B2(new_n774), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1021), .A2(KEYINPUT109), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n660), .A2(G20), .A3(new_n718), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n1021), .B2(KEYINPUT109), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1022), .A2(new_n1024), .B1(new_n713), .B2(new_n941), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT110), .B1(new_n977), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n977), .A2(new_n1025), .A3(KEYINPUT110), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(G393));
  NAND2_X1  g0829(.A1(new_n946), .A2(new_n719), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT111), .Z(new_n1031));
  OAI22_X1  g0831(.A1(new_n745), .A2(new_n725), .B1(new_n729), .B2(new_n733), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT52), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n760), .A2(new_n732), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n318), .B1(new_n723), .B2(new_n1000), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n736), .A2(new_n749), .B1(new_n731), .B2(new_n574), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n757), .A2(new_n460), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n765), .A2(new_n1033), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n741), .A2(G143), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n201), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n318), .B1(new_n1041), .B2(new_n724), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n737), .A2(G68), .B1(new_n769), .B2(new_n304), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G77), .B2(new_n757), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n745), .A2(new_n793), .B1(new_n360), .B2(new_n733), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT51), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n801), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1039), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n774), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n783), .B1(new_n471), .B2(new_n207), .C1(new_n244), .C2(new_n776), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1031), .A2(new_n714), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n938), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n712), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n976), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n667), .B1(new_n938), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1053), .A2(new_n976), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(G390));
  INV_X1    g0859(.A(new_n880), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1060), .B(G330), .C1(new_n888), .C2(new_n889), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n860), .B1(new_n862), .B2(new_n865), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n871), .A2(new_n872), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n870), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n833), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n833), .B(KEYINPUT112), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n883), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n815), .A2(new_n334), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n813), .B1(new_n686), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1069), .B1(new_n1071), .B2(new_n870), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1061), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n708), .A2(G330), .A3(new_n816), .A4(new_n1064), .ZN(new_n1075));
  OAI211_X1 g0875(.A(G330), .B(new_n816), .C1(new_n888), .C2(new_n889), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n870), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n707), .ZN(new_n1079));
  OAI211_X1 g0879(.A(G330), .B(new_n816), .C1(new_n888), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1061), .B1(new_n1081), .B2(new_n1064), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1078), .A2(new_n1071), .B1(new_n1082), .B2(new_n1063), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n890), .A2(new_n436), .A3(new_n655), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n877), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  AND4_X1   g0887(.A1(KEYINPUT113), .A2(new_n1067), .A3(new_n1072), .A4(new_n1075), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1075), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT113), .B1(new_n1090), .B2(new_n1072), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1074), .B(new_n1087), .C1(new_n1088), .C2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1067), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT113), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1090), .A2(KEYINPUT113), .A3(new_n1072), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1073), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT114), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1082), .A2(new_n1063), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1071), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n643), .B(new_n1084), .C1(new_n687), .C2(new_n437), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1103), .A3(KEYINPUT114), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1092), .B(new_n666), .C1(new_n1097), .C2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1062), .A2(new_n717), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n714), .B1(new_n418), .B2(new_n811), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G294), .A2(new_n741), .B1(new_n746), .B2(G283), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n318), .B1(new_n736), .B2(new_n551), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n731), .A2(new_n471), .B1(new_n733), .B2(new_n467), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(G107), .C2(new_n724), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1109), .B(new_n1112), .C1(new_n251), .C2(new_n758), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n737), .A2(new_n991), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT53), .Z(new_n1115));
  NAND2_X1  g0915(.A1(new_n741), .A2(G125), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(new_n201), .C2(new_n754), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n797), .A2(new_n733), .B1(new_n731), .B2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n318), .B(new_n1119), .C1(G137), .C2(new_n724), .ZN(new_n1120));
  INV_X1    g0920(.A(G128), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n745), .C1(new_n360), .C2(new_n758), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n789), .A2(new_n1113), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1108), .B1(new_n1123), .B2(new_n774), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1097), .A2(new_n713), .B1(new_n1107), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1106), .A2(new_n1125), .ZN(G378));
  AOI21_X1  g0926(.A(new_n1086), .B1(new_n1097), .B2(new_n1087), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n886), .ZN(new_n1128));
  OAI21_X1  g0928(.A(G330), .B1(new_n1128), .B2(new_n884), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n866), .A3(new_n875), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n655), .B1(new_n885), .B2(new_n886), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n876), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT118), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT116), .B(KEYINPUT117), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n435), .B(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n424), .A2(new_n649), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1135), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n1134), .A3(new_n1140), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1133), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1130), .A2(new_n1132), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT57), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n666), .B1(new_n1127), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1092), .A2(new_n1103), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1148), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1130), .A2(new_n1132), .A3(new_n1146), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT57), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n717), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n906), .A2(G58), .B1(G283), .B2(new_n741), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n467), .B2(new_n745), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n278), .B(new_n318), .C1(new_n736), .C2(new_n221), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G107), .A2(new_n791), .B1(new_n724), .B2(G97), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n307), .B2(new_n731), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1160), .A2(new_n900), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT58), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n736), .A2(new_n1118), .B1(new_n733), .B2(new_n1121), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n731), .A2(new_n794), .B1(new_n723), .B2(new_n797), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n746), .C2(G125), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n793), .B2(new_n758), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n253), .B(new_n278), .C1(new_n754), .C2(new_n360), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G124), .B2(new_n741), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1164), .A2(KEYINPUT58), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G50), .B1(new_n253), .B2(new_n278), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n282), .B2(G41), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1165), .A2(new_n1174), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n774), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT115), .Z(new_n1180));
  OAI21_X1  g0980(.A(new_n714), .B1(new_n811), .B2(new_n1041), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1154), .A2(new_n713), .B1(new_n1158), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1156), .A2(new_n1183), .ZN(G375));
  AND2_X1   g0984(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n943), .B(KEYINPUT119), .Z(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n714), .B1(new_n811), .B2(G68), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n906), .A2(G58), .B1(G128), .B2(new_n741), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n282), .B1(new_n723), .B2(new_n1118), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n736), .A2(new_n360), .B1(new_n733), .B2(new_n794), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(G150), .C2(new_n769), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n746), .A2(G132), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n757), .A2(G50), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1190), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n318), .B1(new_n723), .B2(new_n459), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n736), .A2(new_n471), .B1(new_n731), .B2(new_n510), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n746), .C2(G294), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n1000), .B2(new_n760), .C1(new_n756), .C2(new_n251), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n995), .B1(new_n749), .B2(new_n733), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT120), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1196), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1189), .B1(new_n1203), .B2(new_n774), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1064), .B2(new_n718), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1083), .B2(new_n712), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1188), .A2(new_n1207), .ZN(G381));
  NAND3_X1  g1008(.A1(new_n1027), .A2(new_n786), .A3(new_n1028), .ZN(new_n1209));
  OR4_X1    g1009(.A1(G384), .A2(new_n1209), .A3(G390), .A4(G381), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1210), .A2(G387), .A3(G375), .A4(G378), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT121), .ZN(G407));
  NAND2_X1  g1012(.A1(new_n1107), .A2(new_n1124), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1074), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(new_n712), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n667), .B1(new_n1185), .B2(new_n1214), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n1092), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n650), .ZN(new_n1218));
  OAI211_X1 g1018(.A(G407), .B(G213), .C1(G375), .C2(new_n1218), .ZN(G409));
  OAI211_X1 g1019(.A(G378), .B(new_n1183), .C1(new_n1150), .C2(new_n1155), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1151), .A2(new_n1154), .A3(new_n1187), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1158), .A2(new_n1182), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1222), .B1(new_n1223), .B2(new_n712), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1217), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1220), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n650), .A2(G213), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1083), .A2(new_n1086), .A3(KEYINPUT60), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT122), .Z(new_n1230));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n667), .B(new_n1087), .C1(new_n1231), .C2(new_n1186), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G384), .B1(new_n1233), .B2(new_n1207), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n823), .B(new_n1206), .C1(new_n1230), .C2(new_n1232), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n650), .A2(G213), .A3(G2897), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1235), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1238), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1228), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n969), .A2(new_n973), .A3(new_n1058), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n786), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n970), .A2(new_n944), .B1(new_n924), .B2(new_n919), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1245), .A2(new_n1209), .B1(new_n1246), .B2(G390), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1209), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT124), .B1(new_n1249), .B2(new_n1244), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT124), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1245), .A2(new_n1251), .A3(new_n1209), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n968), .A2(new_n1058), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1246), .A2(G390), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1250), .B(new_n1252), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1248), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1220), .A2(new_n1225), .B1(G213), .B2(new_n650), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1242), .A2(new_n1256), .A3(new_n1257), .A4(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1226), .A2(new_n1227), .A3(new_n1259), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT123), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1258), .A2(KEYINPUT123), .A3(new_n1259), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1262), .A2(KEYINPUT125), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT125), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1268), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1270), .B1(new_n1271), .B2(new_n1261), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1257), .B1(new_n1274), .B2(new_n1258), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT126), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1242), .A2(new_n1277), .A3(new_n1257), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT62), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1265), .A2(KEYINPUT127), .A3(new_n1280), .A4(new_n1267), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1258), .A2(KEYINPUT62), .A3(new_n1259), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1265), .A2(new_n1280), .A3(new_n1267), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT127), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1279), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1273), .B1(new_n1287), .B2(new_n1256), .ZN(G405));
  AOI21_X1  g1088(.A(G378), .B1(new_n1156), .B2(new_n1183), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1220), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1259), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(new_n1256), .ZN(G402));
endmodule


