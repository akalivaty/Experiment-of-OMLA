//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(G8gat), .Z(new_n207));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208));
  INV_X1    g007(.A(G57gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G64gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT96), .ZN(new_n211));
  INV_X1    g010(.A(G64gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(G57gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT95), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G71gat), .A2(G78gat), .ZN(new_n216));
  OR2_X1    g015(.A1(G71gat), .A2(G78gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT9), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT9), .B1(new_n210), .B2(new_n213), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(new_n216), .A3(new_n217), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(G211gat), .ZN(new_n225));
  XOR2_X1   g024(.A(G127gat), .B(G155gat), .Z(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n208), .ZN(new_n228));
  NAND2_X1  g027(.A1(G231gat), .A2(G233gat), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n228), .B(new_n229), .Z(new_n230));
  OR2_X1    g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n230), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT97), .B(G183gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n234), .B(new_n235), .Z(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n231), .A2(new_n236), .A3(new_n232), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(G190gat), .B(G218gat), .Z(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n242), .A2(KEYINPUT99), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(KEYINPUT99), .ZN(new_n244));
  NAND2_X1  g043(.A1(G85gat), .A2(G92gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT7), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT8), .ZN(new_n247));
  AND2_X1   g046(.A1(G99gat), .A2(G106gat), .ZN(new_n248));
  OAI221_X1 g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .C1(G85gat), .C2(G92gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(G99gat), .A2(G106gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n251), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT98), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n252), .A2(KEYINPUT98), .A3(new_n253), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G43gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G50gat), .ZN(new_n260));
  INV_X1    g059(.A(G50gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G43gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n262), .A3(KEYINPUT15), .ZN(new_n263));
  OR3_X1    g062(.A1(new_n259), .A2(KEYINPUT90), .A3(G50gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(KEYINPUT90), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n264), .A2(new_n260), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT89), .B(KEYINPUT15), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G29gat), .ZN(new_n269));
  INV_X1    g068(.A(G36gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT14), .ZN(new_n272));
  NAND2_X1  g071(.A1(G29gat), .A2(G36gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n273), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n263), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT17), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n277), .A2(KEYINPUT17), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n258), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(G232gat), .A2(G233gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT41), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(new_n258), .B2(new_n277), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n243), .B(new_n244), .C1(new_n281), .C2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n284), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n286), .A2(KEYINPUT99), .A3(new_n280), .A4(new_n242), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT100), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n282), .A2(KEYINPUT41), .ZN(new_n291));
  XNOR2_X1  g090(.A(G134gat), .B(G162gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT100), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n288), .A2(new_n289), .A3(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n220), .A2(new_n222), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n256), .A2(KEYINPUT10), .A3(new_n299), .A4(new_n257), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n254), .A2(new_n223), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n252), .A3(new_n253), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT10), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G230gat), .ZN(new_n306));
  INV_X1    g105(.A(G233gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n301), .A2(new_n302), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G120gat), .B(G148gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(G176gat), .B(G204gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n316), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n310), .A2(new_n312), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n240), .A2(new_n298), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  INV_X1    g122(.A(G169gat), .ZN(new_n324));
  INV_X1    g123(.A(G176gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT26), .ZN(new_n326));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT26), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n323), .B(new_n326), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT68), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT27), .B(G183gat), .ZN(new_n334));
  INV_X1    g133(.A(G190gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT28), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n324), .A2(new_n325), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(new_n328), .A3(new_n327), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n339), .A2(KEYINPUT68), .A3(new_n323), .A4(new_n326), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT28), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n334), .A2(new_n341), .A3(new_n335), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n333), .A2(new_n337), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345));
  INV_X1    g144(.A(G113gat), .ZN(new_n346));
  OR2_X1    g145(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n350));
  INV_X1    g149(.A(G120gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n351), .B2(G113gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n346), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n344), .B(new_n345), .C1(new_n349), .C2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n345), .ZN(new_n356));
  XNOR2_X1  g155(.A(G113gat), .B(G120gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n356), .B1(KEYINPUT1), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT24), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n323), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n362));
  INV_X1    g161(.A(G183gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n335), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT65), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n327), .A2(KEYINPUT23), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n338), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT66), .B(G176gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(KEYINPUT23), .A3(new_n324), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT65), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n361), .A2(new_n364), .A3(new_n371), .A4(new_n362), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n366), .A2(new_n368), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n374));
  AND2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT67), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(new_n363), .A3(new_n335), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n377), .A2(new_n361), .A3(new_n362), .A4(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n330), .B2(KEYINPUT23), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n379), .A2(new_n368), .A3(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n343), .B(new_n359), .C1(new_n375), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G227gat), .A2(G233gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n355), .A2(new_n358), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n382), .B1(new_n373), .B2(new_n374), .ZN(new_n387));
  AND4_X1   g186(.A1(new_n342), .A2(new_n333), .A3(new_n337), .A4(new_n340), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G15gat), .B(G43gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT71), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n394), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(KEYINPUT33), .A3(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n390), .A2(KEYINPUT32), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT32), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT33), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n393), .B1(new_n390), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT73), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT34), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n384), .B2(KEYINPUT72), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n383), .A2(new_n389), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(new_n384), .ZN(new_n407));
  AOI211_X1 g206(.A(new_n385), .B(new_n404), .C1(new_n383), .C2(new_n389), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n402), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT36), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n401), .B2(new_n398), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n398), .A2(new_n401), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n407), .A2(new_n408), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT36), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n411), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G228gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(new_n307), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G141gat), .B(G148gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  OR2_X1    g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(G155gat), .A2(G162gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(KEYINPUT2), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n426), .B(new_n425), .C1(new_n423), .C2(KEYINPUT2), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432));
  OR2_X1    g231(.A1(G197gat), .A2(G204gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(G197gat), .A2(G204gat), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT22), .ZN(new_n435));
  NAND2_X1  g234(.A1(G211gat), .A2(G218gat), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n433), .A2(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(G211gat), .A2(G218gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(G211gat), .A2(G218gat), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT74), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n435), .ZN(new_n442));
  NOR2_X1   g241(.A1(G197gat), .A2(G204gat), .ZN(new_n443));
  AND2_X1   g242(.A1(G197gat), .A2(G204gat), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT74), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n438), .A2(new_n439), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n441), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT75), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n450), .B1(new_n445), .B2(new_n447), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n437), .A2(new_n440), .A3(KEYINPUT75), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT29), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n432), .B1(new_n454), .B2(KEYINPUT80), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n441), .A2(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT80), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT29), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n431), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n456), .B1(new_n460), .B2(KEYINPUT29), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n422), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT29), .B1(new_n453), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n431), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(new_n422), .A3(new_n461), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(G22gat), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G22gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n461), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n457), .B1(new_n456), .B2(KEYINPUT29), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n453), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT29), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(KEYINPUT80), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(new_n474), .A3(new_n432), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n470), .B1(new_n475), .B2(new_n431), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n469), .B(new_n466), .C1(new_n476), .C2(new_n422), .ZN(new_n477));
  XNOR2_X1  g276(.A(G78gat), .B(G106gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT31), .B(G50gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n468), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT81), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n468), .A2(KEYINPUT81), .A3(new_n477), .A4(new_n481), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n477), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(new_n480), .ZN(new_n489));
  AOI211_X1 g288(.A(KEYINPUT82), .B(new_n481), .C1(new_n468), .C2(new_n477), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n473), .B1(new_n387), .B2(new_n388), .ZN(new_n492));
  INV_X1    g291(.A(G226gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(new_n307), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n387), .B2(new_n388), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n456), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT76), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n492), .A2(new_n499), .A3(new_n495), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n492), .B2(new_n495), .ZN(new_n501));
  INV_X1    g300(.A(new_n497), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n498), .B1(new_n503), .B2(new_n456), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n505));
  XNOR2_X1  g304(.A(G8gat), .B(G36gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(G64gat), .B(G92gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n504), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n498), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT76), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n492), .A2(new_n499), .A3(new_n495), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n497), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n511), .B1(new_n514), .B2(new_n472), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n505), .B1(new_n515), .B2(new_n508), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n504), .A2(new_n509), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G1gat), .B(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G85gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT0), .B(G57gat), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n521), .B(new_n522), .Z(new_n523));
  INV_X1    g322(.A(KEYINPUT4), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n429), .A2(new_n430), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n386), .A2(KEYINPUT77), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT77), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n355), .A2(new_n429), .A3(new_n430), .A4(new_n358), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(KEYINPUT4), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(KEYINPUT4), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G225gat), .A2(G233gat), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n432), .B1(new_n429), .B2(new_n430), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n460), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n535), .B2(new_n359), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n531), .A2(KEYINPUT78), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT78), .B1(new_n531), .B2(new_n536), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n359), .B(new_n525), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT5), .B1(new_n539), .B2(new_n532), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n386), .A2(KEYINPUT79), .A3(new_n524), .A4(new_n525), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT79), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n528), .B2(KEYINPUT4), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n544), .A3(new_n530), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT5), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n546), .A3(new_n536), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n523), .B1(new_n541), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT6), .ZN(new_n550));
  INV_X1    g349(.A(new_n538), .ZN(new_n551));
  INV_X1    g350(.A(new_n540), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n531), .A2(KEYINPUT78), .A3(new_n536), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n523), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n547), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n549), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  OAI211_X1 g356(.A(KEYINPUT6), .B(new_n523), .C1(new_n541), .C2(new_n548), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n510), .A2(new_n518), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n419), .B1(new_n491), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n472), .A2(new_n473), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT3), .B1(new_n561), .B2(new_n457), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n525), .B1(new_n562), .B2(new_n474), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n421), .B1(new_n563), .B2(new_n470), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n469), .B1(new_n564), .B2(new_n466), .ZN(new_n565));
  INV_X1    g364(.A(new_n477), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n480), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT82), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n488), .A2(new_n487), .A3(new_n480), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n568), .A2(new_n569), .B1(new_n484), .B2(new_n485), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n535), .A2(new_n359), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n545), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n533), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT83), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT83), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n575), .A3(new_n533), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT39), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n577), .B1(new_n539), .B2(new_n532), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n575), .B1(new_n572), .B2(new_n533), .ZN(new_n580));
  AOI211_X1 g379(.A(KEYINPUT83), .B(new_n532), .C1(new_n545), .C2(new_n571), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n579), .A2(new_n582), .A3(KEYINPUT40), .A4(new_n555), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n518), .A2(new_n510), .A3(new_n549), .A4(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n579), .A2(new_n582), .A3(new_n555), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT84), .B(KEYINPUT40), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n586), .A2(KEYINPUT85), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT85), .B1(new_n586), .B2(new_n587), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n570), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n557), .A2(new_n558), .A3(new_n517), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT38), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n593), .B(new_n508), .C1(new_n515), .C2(KEYINPUT37), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n496), .A2(new_n497), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n472), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n514), .B2(new_n472), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT86), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n599), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n509), .B1(new_n504), .B2(new_n598), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT86), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n593), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n508), .B1(new_n515), .B2(KEYINPUT37), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n504), .A2(new_n598), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT38), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n592), .A2(new_n600), .A3(new_n604), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n560), .B1(new_n591), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n491), .A2(new_n559), .A3(new_n410), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n568), .A2(new_n569), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n416), .B1(new_n611), .B2(new_n486), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n518), .A2(new_n510), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n557), .A2(new_n558), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n610), .A2(KEYINPUT35), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT87), .B1(new_n609), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n610), .A2(KEYINPUT35), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n612), .A2(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n613), .A2(new_n614), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n570), .A2(new_n622), .B1(new_n418), .B2(new_n411), .ZN(new_n623));
  INV_X1    g422(.A(new_n589), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n586), .A2(KEYINPUT85), .A3(new_n587), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n491), .B1(new_n626), .B2(new_n584), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n607), .A2(new_n558), .A3(new_n557), .A4(new_n517), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n604), .A2(new_n600), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n623), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT87), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n621), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n634));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G169gat), .B(G197gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT91), .ZN(new_n641));
  OR3_X1    g440(.A1(new_n277), .A2(new_n207), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n641), .B1(new_n277), .B2(new_n207), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G229gat), .A2(G233gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n279), .A2(new_n207), .A3(new_n278), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT18), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT92), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n642), .A2(new_n643), .B1(new_n277), .B2(new_n207), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n645), .B(KEYINPUT13), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n277), .A2(new_n207), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n644), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n652), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(KEYINPUT92), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n649), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n647), .A2(new_n648), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n640), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n649), .B2(KEYINPUT93), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n639), .B1(new_n657), .B2(new_n653), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT93), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n647), .A2(new_n664), .A3(new_n648), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n618), .A2(new_n633), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT94), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n618), .A2(new_n633), .A3(KEYINPUT94), .A4(new_n667), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n322), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n614), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  INV_X1    g474(.A(new_n613), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT101), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT42), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(G8gat), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n683));
  OAI211_X1 g482(.A(KEYINPUT101), .B(new_n683), .C1(new_n677), .C2(new_n679), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(G1325gat));
  AND4_X1   g484(.A1(G15gat), .A2(new_n672), .A3(new_n418), .A4(new_n411), .ZN(new_n686));
  INV_X1    g485(.A(new_n416), .ZN(new_n687));
  AOI21_X1  g486(.A(G15gat), .B1(new_n672), .B2(new_n687), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n686), .A2(new_n688), .A3(KEYINPUT102), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT102), .B1(new_n686), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1326gat));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n570), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT43), .B(G22gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(new_n298), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n618), .A2(new_n633), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT44), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n698), .B(new_n695), .C1(new_n609), .C2(new_n617), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT103), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n621), .A2(new_n631), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n698), .A4(new_n695), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n697), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n240), .A2(new_n320), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n667), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(G29gat), .B1(new_n709), .B2(new_n614), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n670), .A2(new_n671), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n240), .A2(new_n298), .A3(new_n320), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n711), .A2(new_n269), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n713), .A2(new_n714), .A3(new_n673), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n713), .B2(new_n673), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n710), .B1(new_n715), .B2(new_n716), .ZN(G1328gat));
  OAI21_X1  g516(.A(G36gat), .B1(new_n709), .B2(new_n613), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n613), .A2(G36gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n711), .A2(new_n712), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT46), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n711), .A2(new_n722), .A3(new_n712), .A4(new_n719), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n718), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n718), .A2(new_n721), .A3(new_n726), .A4(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1329gat));
  NAND4_X1  g527(.A1(new_n711), .A2(new_n259), .A3(new_n687), .A4(new_n712), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n709), .A2(new_n419), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(new_n259), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT47), .B1(new_n729), .B2(KEYINPUT105), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI221_X1 g532(.A(new_n729), .B1(KEYINPUT105), .B2(KEYINPUT47), .C1(new_n730), .C2(new_n259), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(G1330gat));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n707), .B1(new_n697), .B2(new_n704), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n261), .B1(new_n737), .B2(new_n570), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n491), .A2(G50gat), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n711), .A2(new_n712), .A3(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n736), .B(KEYINPUT48), .C1(new_n738), .C2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n711), .A2(new_n712), .A3(new_n739), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n491), .B(new_n707), .C1(new_n697), .C2(new_n704), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(new_n261), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT48), .B1(new_n745), .B2(new_n736), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n742), .A2(new_n746), .ZN(G1331gat));
  NOR2_X1   g546(.A1(new_n667), .A2(new_n321), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n701), .A2(new_n240), .A3(new_n298), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n614), .B(KEYINPUT107), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(new_n209), .ZN(G1332gat));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n613), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  AND2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n753), .B2(new_n754), .ZN(G1333gat));
  INV_X1    g556(.A(G71gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n749), .B2(new_n416), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n749), .A2(new_n758), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(new_n419), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g561(.A1(new_n749), .A2(new_n491), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT108), .B(G78gat), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1335gat));
  NOR3_X1   g564(.A1(new_n240), .A2(new_n667), .A3(new_n321), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n705), .A2(new_n766), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n767), .A2(new_n520), .A3(new_n614), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n298), .B1(new_n621), .B2(new_n631), .ZN(new_n769));
  INV_X1    g568(.A(new_n667), .ZN(new_n770));
  INV_X1    g569(.A(new_n240), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT51), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n769), .A2(new_n774), .A3(new_n770), .A4(new_n771), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n773), .A2(new_n320), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n673), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n768), .A2(new_n777), .ZN(G1336gat));
  AOI21_X1  g577(.A(G92gat), .B1(new_n776), .B2(new_n676), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n676), .A2(G92gat), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n767), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT52), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n779), .B2(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1337gat));
  XNOR2_X1  g585(.A(KEYINPUT109), .B(G99gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n776), .A2(new_n687), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n767), .A2(new_n419), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(new_n787), .ZN(G1338gat));
  NAND3_X1  g589(.A1(new_n705), .A2(new_n570), .A3(new_n766), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(G106gat), .ZN(new_n792));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n776), .A2(new_n793), .A3(new_n570), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT53), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n791), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n705), .A2(KEYINPUT111), .A3(new_n570), .A4(new_n766), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n799), .A2(G106gat), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n795), .B1(new_n797), .B2(new_n801), .ZN(G1339gat));
  NOR2_X1   g601(.A1(new_n655), .A2(new_n656), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n645), .B1(new_n644), .B2(new_n646), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n638), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n666), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n298), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n300), .A2(new_n304), .A3(new_n308), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n310), .A2(KEYINPUT54), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n308), .B1(new_n300), .B2(new_n304), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n318), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n809), .A2(KEYINPUT55), .A3(new_n812), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n319), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT112), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n815), .A2(new_n819), .A3(new_n319), .A4(new_n816), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n807), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n666), .A2(new_n320), .A3(new_n805), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n824), .B1(new_n821), .B2(new_n667), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n822), .B1(new_n825), .B2(new_n695), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n771), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n322), .A2(new_n667), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n750), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n613), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n491), .A2(new_n410), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT113), .B1(new_n832), .B2(new_n835), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n667), .A2(new_n346), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT114), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n828), .B1(new_n826), .B2(new_n771), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(new_n570), .A3(new_n416), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n676), .A2(new_n614), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n770), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT115), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n841), .A2(new_n849), .A3(new_n846), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(G1340gat));
  NAND2_X1  g650(.A1(new_n347), .A2(new_n348), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n320), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(KEYINPUT116), .Z(new_n854));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n838), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G120gat), .B1(new_n845), .B2(new_n321), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1341gat));
  NOR2_X1   g656(.A1(new_n832), .A2(new_n835), .ZN(new_n858));
  AOI21_X1  g657(.A(G127gat), .B1(new_n858), .B2(new_n240), .ZN(new_n859));
  INV_X1    g658(.A(G127gat), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n845), .A2(new_n860), .A3(new_n771), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n859), .A2(new_n861), .ZN(G1342gat));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n695), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n845), .B2(new_n298), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT56), .B1(new_n863), .B2(G134gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n830), .A2(new_n868), .A3(new_n570), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n844), .A2(new_n419), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n817), .B1(new_n661), .B2(new_n666), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n298), .B1(new_n871), .B2(new_n824), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n822), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n817), .ZN(new_n875));
  INV_X1    g674(.A(new_n666), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n660), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n695), .B1(new_n877), .B2(new_n823), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(KEYINPUT117), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n771), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n491), .B1(new_n880), .B2(new_n829), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n869), .B(new_n870), .C1(new_n881), .C2(new_n868), .ZN(new_n882));
  OAI21_X1  g681(.A(G141gat), .B1(new_n882), .B2(new_n770), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n419), .A2(new_n570), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n832), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(G141gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n886), .A3(new_n667), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT58), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n883), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1344gat));
  INV_X1    g691(.A(G148gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n885), .A2(new_n893), .A3(new_n320), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(new_n882), .B2(new_n321), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n893), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n298), .A2(new_n817), .A3(new_n806), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n771), .B1(new_n878), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n491), .B1(new_n829), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT119), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n818), .A2(new_n820), .B1(new_n661), .B2(new_n666), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n298), .B1(new_n902), .B2(new_n824), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n240), .B1(new_n903), .B2(new_n822), .ZN(new_n904));
  OAI211_X1 g703(.A(KEYINPUT57), .B(new_n570), .C1(new_n904), .C2(new_n828), .ZN(new_n905));
  INV_X1    g704(.A(new_n898), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n240), .B1(new_n872), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n570), .B1(new_n907), .B2(new_n828), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n868), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n901), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT118), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n870), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n870), .A2(new_n912), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n911), .A2(new_n320), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n895), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n894), .B1(new_n897), .B2(new_n916), .ZN(G1345gat));
  AOI21_X1  g716(.A(G155gat), .B1(new_n885), .B2(new_n240), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n882), .A2(new_n771), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g719(.A(G162gat), .B1(new_n885), .B2(new_n695), .ZN(new_n921));
  INV_X1    g720(.A(G162gat), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n882), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n923), .B2(new_n695), .ZN(G1347gat));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n842), .B2(new_n673), .ZN(new_n926));
  OAI211_X1 g725(.A(KEYINPUT120), .B(new_n614), .C1(new_n904), .C2(new_n828), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n836), .A2(new_n676), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT121), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n324), .A3(new_n667), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n831), .A2(new_n613), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n830), .A2(new_n612), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n770), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(G1348gat));
  NOR3_X1   g735(.A1(new_n934), .A2(new_n369), .A3(new_n321), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n928), .A2(new_n320), .A3(new_n930), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n939));
  OR3_X1    g738(.A1(new_n938), .A2(new_n939), .A3(G176gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n938), .B2(G176gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G1349gat));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n934), .B2(new_n771), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n843), .A2(KEYINPUT123), .A3(new_n240), .A4(new_n933), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n945), .A3(G183gat), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n928), .A2(new_n334), .A3(new_n240), .A4(new_n930), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(KEYINPUT124), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT60), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT60), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n946), .A2(KEYINPUT124), .A3(new_n950), .A4(new_n947), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n934), .B2(new_n298), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT61), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n931), .A2(new_n335), .A3(new_n695), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1351gat));
  AOI21_X1  g755(.A(new_n884), .B1(new_n926), .B2(new_n927), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(new_n676), .ZN(new_n958));
  INV_X1    g757(.A(G197gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n958), .A2(new_n959), .A3(new_n667), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n933), .A2(new_n419), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n911), .A2(new_n667), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n959), .B2(new_n962), .ZN(G1352gat));
  XNOR2_X1  g762(.A(KEYINPUT125), .B(G204gat), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n957), .A2(new_n676), .A3(new_n320), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT126), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n911), .A2(new_n320), .A3(new_n961), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(new_n964), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n966), .A2(new_n972), .A3(KEYINPUT62), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n968), .A2(new_n969), .A3(new_n971), .A4(new_n973), .ZN(G1353gat));
  INV_X1    g773(.A(G211gat), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n975), .A3(new_n240), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n911), .A2(new_n240), .A3(new_n961), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n977), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT63), .B1(new_n977), .B2(G211gat), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(G1354gat));
  INV_X1    g779(.A(G218gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n958), .A2(new_n981), .A3(new_n695), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n911), .A2(new_n983), .A3(new_n961), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n911), .B2(new_n961), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n984), .A2(new_n985), .A3(new_n298), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n982), .B1(new_n986), .B2(new_n981), .ZN(G1355gat));
endmodule


