

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X1 U325 ( .A(n471), .B(KEYINPUT119), .ZN(n472) );
  NAND2_X1 U326 ( .A1(n561), .A2(n560), .ZN(n293) );
  XNOR2_X1 U327 ( .A(n395), .B(KEYINPUT25), .ZN(n396) );
  XNOR2_X1 U328 ( .A(n397), .B(n396), .ZN(n401) );
  XNOR2_X1 U329 ( .A(n413), .B(n347), .ZN(n348) );
  XNOR2_X1 U330 ( .A(n388), .B(n348), .ZN(n349) );
  XNOR2_X1 U331 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U332 ( .A(n354), .B(n353), .ZN(n356) );
  XNOR2_X1 U333 ( .A(n333), .B(n332), .ZN(n334) );
  INV_X1 U334 ( .A(KEYINPUT55), .ZN(n471) );
  XNOR2_X1 U335 ( .A(n335), .B(n334), .ZN(n340) );
  XNOR2_X1 U336 ( .A(n351), .B(n434), .ZN(n341) );
  XNOR2_X1 U337 ( .A(n473), .B(n472), .ZN(n562) );
  XNOR2_X1 U338 ( .A(n342), .B(n341), .ZN(n577) );
  XNOR2_X1 U339 ( .A(n474), .B(G190GAT), .ZN(n475) );
  XNOR2_X1 U340 ( .A(n451), .B(G29GAT), .ZN(n452) );
  XNOR2_X1 U341 ( .A(n476), .B(n475), .ZN(G1351GAT) );
  XNOR2_X1 U342 ( .A(n453), .B(n452), .ZN(G1328GAT) );
  XOR2_X1 U343 ( .A(G127GAT), .B(KEYINPUT78), .Z(n295) );
  XNOR2_X1 U344 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n350) );
  XOR2_X1 U346 ( .A(n350), .B(KEYINPUT89), .Z(n297) );
  NAND2_X1 U347 ( .A1(G225GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U349 ( .A(G57GAT), .B(KEYINPUT87), .Z(n299) );
  XNOR2_X1 U350 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U353 ( .A(KEYINPUT86), .B(G148GAT), .Z(n303) );
  XNOR2_X1 U354 ( .A(G141GAT), .B(G120GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n305), .B(n304), .ZN(n310) );
  XOR2_X1 U357 ( .A(G85GAT), .B(G162GAT), .Z(n308) );
  XNOR2_X1 U358 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n306), .B(KEYINPUT2), .ZN(n362) );
  XNOR2_X1 U360 ( .A(G29GAT), .B(n362), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U362 ( .A(n310), .B(n309), .Z(n315) );
  XOR2_X1 U363 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n312) );
  XNOR2_X1 U364 ( .A(G1GAT), .B(KEYINPUT88), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U366 ( .A(G134GAT), .B(n313), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n543) );
  XOR2_X1 U368 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n317) );
  NAND2_X1 U369 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U371 ( .A(n318), .B(KEYINPUT30), .Z(n320) );
  XOR2_X1 U372 ( .A(G141GAT), .B(G22GAT), .Z(n366) );
  XOR2_X1 U373 ( .A(G169GAT), .B(G8GAT), .Z(n381) );
  XNOR2_X1 U374 ( .A(n366), .B(n381), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U376 ( .A(G15GAT), .B(G1GAT), .Z(n435) );
  XOR2_X1 U377 ( .A(n321), .B(n435), .Z(n323) );
  XNOR2_X1 U378 ( .A(G113GAT), .B(G197GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n328) );
  XNOR2_X1 U380 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n324), .B(G29GAT), .ZN(n325) );
  XOR2_X1 U382 ( .A(n325), .B(KEYINPUT8), .Z(n327) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(G50GAT), .ZN(n326) );
  XOR2_X1 U384 ( .A(n327), .B(n326), .Z(n420) );
  XOR2_X1 U385 ( .A(n328), .B(n420), .Z(n546) );
  XOR2_X1 U386 ( .A(n546), .B(KEYINPUT66), .Z(n557) );
  XNOR2_X1 U387 ( .A(G99GAT), .B(G85GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n329), .B(KEYINPUT67), .ZN(n410) );
  XOR2_X1 U389 ( .A(n410), .B(KEYINPUT33), .Z(n335) );
  XOR2_X1 U390 ( .A(KEYINPUT69), .B(KEYINPUT32), .Z(n331) );
  XNOR2_X1 U391 ( .A(KEYINPUT31), .B(KEYINPUT68), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n333) );
  NAND2_X1 U393 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  XOR2_X1 U394 ( .A(G78GAT), .B(G148GAT), .Z(n337) );
  XNOR2_X1 U395 ( .A(G106GAT), .B(G204GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n363) );
  XNOR2_X1 U397 ( .A(G176GAT), .B(G92GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n338), .B(G64GAT), .ZN(n384) );
  XOR2_X1 U399 ( .A(n363), .B(n384), .Z(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n342) );
  XOR2_X1 U401 ( .A(G120GAT), .B(G71GAT), .Z(n351) );
  XOR2_X1 U402 ( .A(G57GAT), .B(KEYINPUT13), .Z(n434) );
  INV_X1 U403 ( .A(n577), .ZN(n461) );
  NAND2_X1 U404 ( .A1(n557), .A2(n461), .ZN(n487) );
  XOR2_X1 U405 ( .A(KEYINPUT79), .B(KEYINPUT20), .Z(n344) );
  XNOR2_X1 U406 ( .A(G169GAT), .B(G15GAT), .ZN(n343) );
  XNOR2_X1 U407 ( .A(n344), .B(n343), .ZN(n358) );
  XOR2_X1 U408 ( .A(G183GAT), .B(KEYINPUT17), .Z(n346) );
  XNOR2_X1 U409 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n388) );
  XOR2_X1 U411 ( .A(G190GAT), .B(G134GAT), .Z(n413) );
  AND2_X1 U412 ( .A1(G227GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n349), .B(G176GAT), .ZN(n354) );
  XOR2_X1 U414 ( .A(n350), .B(KEYINPUT80), .Z(n352) );
  XOR2_X1 U415 ( .A(G43GAT), .B(G99GAT), .Z(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U417 ( .A(n358), .B(n357), .Z(n398) );
  INV_X1 U418 ( .A(n398), .ZN(n561) );
  INV_X1 U419 ( .A(n561), .ZN(n525) );
  XOR2_X1 U420 ( .A(KEYINPUT85), .B(KEYINPUT23), .Z(n360) );
  NAND2_X1 U421 ( .A1(G228GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U423 ( .A(n361), .B(KEYINPUT24), .Z(n365) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n370) );
  XOR2_X1 U426 ( .A(KEYINPUT22), .B(KEYINPUT81), .Z(n368) );
  XOR2_X1 U427 ( .A(KEYINPUT70), .B(G162GAT), .Z(n412) );
  XNOR2_X1 U428 ( .A(n366), .B(n412), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U430 ( .A(n370), .B(n369), .Z(n372) );
  XNOR2_X1 U431 ( .A(G50GAT), .B(KEYINPUT84), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n377) );
  XOR2_X1 U433 ( .A(KEYINPUT21), .B(KEYINPUT83), .Z(n374) );
  XNOR2_X1 U434 ( .A(G197GAT), .B(G211GAT), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n376) );
  XOR2_X1 U436 ( .A(G218GAT), .B(KEYINPUT82), .Z(n375) );
  XOR2_X1 U437 ( .A(n376), .B(n375), .Z(n386) );
  XOR2_X1 U438 ( .A(n377), .B(n386), .Z(n470) );
  XOR2_X1 U439 ( .A(n470), .B(KEYINPUT28), .Z(n522) );
  XOR2_X1 U440 ( .A(KEYINPUT90), .B(G204GAT), .Z(n379) );
  XNOR2_X1 U441 ( .A(G36GAT), .B(G190GAT), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U443 ( .A(n381), .B(n380), .Z(n383) );
  NAND2_X1 U444 ( .A1(G226GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U446 ( .A(n385), .B(n384), .Z(n390) );
  INV_X1 U447 ( .A(n386), .ZN(n387) );
  XOR2_X1 U448 ( .A(n388), .B(n387), .Z(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n514) );
  XNOR2_X1 U450 ( .A(n514), .B(KEYINPUT27), .ZN(n400) );
  INV_X1 U451 ( .A(n400), .ZN(n391) );
  NAND2_X1 U452 ( .A1(n522), .A2(n391), .ZN(n392) );
  NOR2_X1 U453 ( .A1(n543), .A2(n392), .ZN(n527) );
  NAND2_X1 U454 ( .A1(n525), .A2(n527), .ZN(n393) );
  XNOR2_X1 U455 ( .A(KEYINPUT91), .B(n393), .ZN(n407) );
  NOR2_X1 U456 ( .A1(n398), .A2(n514), .ZN(n394) );
  NOR2_X1 U457 ( .A1(n394), .A2(n470), .ZN(n397) );
  INV_X1 U458 ( .A(KEYINPUT92), .ZN(n395) );
  NAND2_X1 U459 ( .A1(n470), .A2(n398), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n399), .B(KEYINPUT26), .ZN(n570) );
  NOR2_X1 U461 ( .A1(n570), .A2(n400), .ZN(n545) );
  NOR2_X1 U462 ( .A1(n401), .A2(n545), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n402), .B(KEYINPUT93), .ZN(n403) );
  NAND2_X1 U464 ( .A1(n403), .A2(n543), .ZN(n405) );
  INV_X1 U465 ( .A(KEYINPUT94), .ZN(n404) );
  XNOR2_X1 U466 ( .A(n405), .B(n404), .ZN(n406) );
  NOR2_X1 U467 ( .A1(n407), .A2(n406), .ZN(n483) );
  XOR2_X1 U468 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n409) );
  XNOR2_X1 U469 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U471 ( .A(n411), .B(n410), .Z(n415) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U474 ( .A(G92GAT), .B(KEYINPUT71), .Z(n417) );
  NAND2_X1 U475 ( .A1(G232GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U477 ( .A(n419), .B(n418), .Z(n422) );
  XOR2_X1 U478 ( .A(n420), .B(G106GAT), .Z(n421) );
  XOR2_X1 U479 ( .A(n422), .B(n421), .Z(n537) );
  XNOR2_X1 U480 ( .A(n537), .B(KEYINPUT99), .ZN(n423) );
  XNOR2_X1 U481 ( .A(KEYINPUT36), .B(n423), .ZN(n586) );
  XOR2_X1 U482 ( .A(KEYINPUT77), .B(KEYINPUT73), .Z(n425) );
  XNOR2_X1 U483 ( .A(KEYINPUT76), .B(KEYINPUT74), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n445) );
  XOR2_X1 U485 ( .A(KEYINPUT75), .B(G64GAT), .Z(n427) );
  XNOR2_X1 U486 ( .A(G8GAT), .B(G155GAT), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U488 ( .A(G78GAT), .B(G211GAT), .Z(n429) );
  XNOR2_X1 U489 ( .A(G22GAT), .B(G71GAT), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n443) );
  XOR2_X1 U492 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n433) );
  XNOR2_X1 U493 ( .A(KEYINPUT12), .B(KEYINPUT72), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n439) );
  XOR2_X1 U495 ( .A(n434), .B(G183GAT), .Z(n437) );
  XNOR2_X1 U496 ( .A(n435), .B(G127GAT), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U498 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U499 ( .A1(G231GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U502 ( .A(n445), .B(n444), .Z(n552) );
  INV_X1 U503 ( .A(n552), .ZN(n580) );
  OR2_X1 U504 ( .A1(n586), .A2(n580), .ZN(n446) );
  OR2_X1 U505 ( .A1(n483), .A2(n446), .ZN(n447) );
  XOR2_X1 U506 ( .A(n447), .B(KEYINPUT37), .Z(n511) );
  NOR2_X1 U507 ( .A1(n487), .A2(n511), .ZN(n449) );
  XNOR2_X1 U508 ( .A(KEYINPUT38), .B(KEYINPUT100), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U510 ( .A(KEYINPUT101), .B(n450), .ZN(n498) );
  NOR2_X1 U511 ( .A1(n543), .A2(n498), .ZN(n453) );
  XNOR2_X1 U512 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n451) );
  INV_X1 U513 ( .A(n537), .ZN(n555) );
  XOR2_X1 U514 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n456) );
  INV_X1 U515 ( .A(n546), .ZN(n573) );
  XNOR2_X1 U516 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n454) );
  XOR2_X1 U517 ( .A(n454), .B(n577), .Z(n560) );
  NAND2_X1 U518 ( .A1(n573), .A2(n560), .ZN(n455) );
  XNOR2_X1 U519 ( .A(n456), .B(n455), .ZN(n457) );
  NOR2_X1 U520 ( .A1(n457), .A2(n580), .ZN(n458) );
  NAND2_X1 U521 ( .A1(n555), .A2(n458), .ZN(n459) );
  XNOR2_X1 U522 ( .A(n459), .B(KEYINPUT47), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n552), .A2(n586), .ZN(n460) );
  XNOR2_X1 U524 ( .A(n460), .B(KEYINPUT45), .ZN(n462) );
  NAND2_X1 U525 ( .A1(n462), .A2(n461), .ZN(n463) );
  NOR2_X1 U526 ( .A1(n557), .A2(n463), .ZN(n464) );
  NOR2_X1 U527 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT48), .ZN(n542) );
  NOR2_X1 U529 ( .A1(n514), .A2(n542), .ZN(n468) );
  XNOR2_X1 U530 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n467) );
  XNOR2_X1 U531 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U532 ( .A1(n469), .A2(n543), .ZN(n571) );
  NOR2_X1 U533 ( .A1(n470), .A2(n571), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n525), .A2(n562), .ZN(n566) );
  NAND2_X1 U535 ( .A1(n566), .A2(n537), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n474) );
  INV_X1 U537 ( .A(G43GAT), .ZN(n480) );
  NOR2_X1 U538 ( .A1(n498), .A2(n525), .ZN(n478) );
  XNOR2_X1 U539 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1330GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n482) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n482), .B(n481), .ZN(n490) );
  NOR2_X1 U545 ( .A1(n552), .A2(n537), .ZN(n484) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  NOR2_X1 U547 ( .A1(n483), .A2(n485), .ZN(n486) );
  XNOR2_X1 U548 ( .A(KEYINPUT95), .B(n486), .ZN(n500) );
  NOR2_X1 U549 ( .A1(n500), .A2(n487), .ZN(n488) );
  XOR2_X1 U550 ( .A(KEYINPUT96), .B(n488), .Z(n494) );
  NOR2_X1 U551 ( .A1(n543), .A2(n494), .ZN(n489) );
  XOR2_X1 U552 ( .A(n490), .B(n489), .Z(G1324GAT) );
  NOR2_X1 U553 ( .A1(n514), .A2(n494), .ZN(n491) );
  XOR2_X1 U554 ( .A(G8GAT), .B(n491), .Z(G1325GAT) );
  XNOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n493) );
  NOR2_X1 U556 ( .A1(n525), .A2(n494), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  NOR2_X1 U558 ( .A1(n522), .A2(n494), .ZN(n495) );
  XOR2_X1 U559 ( .A(G22GAT), .B(n495), .Z(G1327GAT) );
  NOR2_X1 U560 ( .A1(n514), .A2(n498), .ZN(n497) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(G1329GAT) );
  NOR2_X1 U563 ( .A1(n522), .A2(n498), .ZN(n499) );
  XOR2_X1 U564 ( .A(G50GAT), .B(n499), .Z(G1331GAT) );
  NAND2_X1 U565 ( .A1(n546), .A2(n560), .ZN(n510) );
  OR2_X1 U566 ( .A1(n500), .A2(n510), .ZN(n506) );
  NOR2_X1 U567 ( .A1(n543), .A2(n506), .ZN(n501) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n501), .Z(n502) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(n502), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n514), .A2(n506), .ZN(n503) );
  XOR2_X1 U571 ( .A(G64GAT), .B(n503), .Z(G1333GAT) );
  NOR2_X1 U572 ( .A1(n525), .A2(n506), .ZN(n505) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n504) );
  XNOR2_X1 U574 ( .A(n505), .B(n504), .ZN(G1334GAT) );
  NOR2_X1 U575 ( .A1(n522), .A2(n506), .ZN(n508) );
  XNOR2_X1 U576 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U577 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n509), .ZN(G1335GAT) );
  OR2_X1 U579 ( .A1(n511), .A2(n510), .ZN(n521) );
  NOR2_X1 U580 ( .A1(n543), .A2(n521), .ZN(n513) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n512) );
  XNOR2_X1 U582 ( .A(n513), .B(n512), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n514), .A2(n521), .ZN(n515) );
  XOR2_X1 U584 ( .A(KEYINPUT108), .B(n515), .Z(n516) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n516), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n525), .A2(n521), .ZN(n518) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n517) );
  XNOR2_X1 U588 ( .A(n518), .B(n517), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n520) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n519) );
  XNOR2_X1 U591 ( .A(n520), .B(n519), .ZN(n524) );
  NOR2_X1 U592 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U593 ( .A(n524), .B(n523), .Z(G1339GAT) );
  NOR2_X1 U594 ( .A1(n542), .A2(n525), .ZN(n526) );
  NAND2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U596 ( .A(KEYINPUT113), .B(n528), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n557), .A2(n538), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n529), .B(KEYINPUT114), .ZN(n530) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U601 ( .A1(n538), .A2(n560), .ZN(n531) );
  XNOR2_X1 U602 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n536) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n534) );
  NAND2_X1 U605 ( .A1(n538), .A2(n580), .ZN(n533) );
  XNOR2_X1 U606 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U607 ( .A(n536), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U609 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U610 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n541), .Z(G1343GAT) );
  NOR2_X1 U612 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U613 ( .A1(n545), .A2(n544), .ZN(n554) );
  NOR2_X1 U614 ( .A1(n546), .A2(n554), .ZN(n547) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n547), .Z(G1344GAT) );
  INV_X1 U616 ( .A(n560), .ZN(n548) );
  NOR2_X1 U617 ( .A1(n548), .A2(n554), .ZN(n550) );
  XNOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NOR2_X1 U621 ( .A1(n552), .A2(n554), .ZN(n553) );
  XOR2_X1 U622 ( .A(G155GAT), .B(n553), .Z(G1346GAT) );
  NOR2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n556), .Z(G1347GAT) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n566), .A2(n557), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n564) );
  OR2_X1 U629 ( .A1(n293), .A2(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U632 ( .A1(n580), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n569) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n575) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(n572), .B(KEYINPUT122), .Z(n587) );
  INV_X1 U639 ( .A(n587), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n581), .A2(n573), .ZN(n574) );
  XOR2_X1 U641 ( .A(n575), .B(n574), .Z(n576) );
  XNOR2_X1 U642 ( .A(KEYINPUT123), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  NAND2_X1 U644 ( .A1(n577), .A2(n581), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  XOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT125), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n585) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n589) );
  NOR2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U653 ( .A(n589), .B(n588), .Z(G1355GAT) );
endmodule

