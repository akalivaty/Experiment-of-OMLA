//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n216), .A2(G50), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G116), .ZN(new_n221));
  INV_X1    g0021(.A(G270), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT66), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(new_n223), .A2(new_n224), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G97), .A2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G58), .A2(G232), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G87), .ZN(new_n230));
  INV_X1    g0030(.A(G250), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n208), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n211), .B1(new_n214), .B2(new_n218), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n222), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n202), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G274), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT67), .B(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n220), .A2(G1698), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n257), .A2(new_n260), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G87), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G1), .A3(G13), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n255), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT71), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G232), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n268), .A2(new_n272), .A3(KEYINPUT71), .A4(G232), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n270), .A2(G190), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G200), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n279), .B1(new_n270), .B2(new_n277), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT8), .B(G58), .Z(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G20), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G1), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G13), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n212), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n284), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n286), .B1(new_n289), .B2(new_n282), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n278), .A2(new_n280), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G58), .ZN(new_n293));
  INV_X1    g0093(.A(G68), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(G20), .B1(new_n295), .B2(new_n201), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G159), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT3), .B(G33), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT7), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n301), .A2(new_n302), .A3(G20), .ZN(new_n303));
  AOI21_X1  g0103(.A(G20), .B1(new_n257), .B2(new_n262), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT70), .B1(new_n304), .B2(KEYINPUT7), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n306), .B(new_n302), .C1(new_n301), .C2(G20), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n303), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(KEYINPUT16), .B(new_n300), .C1(new_n308), .C2(new_n294), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT16), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n302), .B1(new_n301), .B2(G20), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n257), .A2(new_n262), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(KEYINPUT7), .A3(new_n283), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n294), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n310), .B1(new_n314), .B2(new_n299), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n309), .A2(new_n288), .A3(new_n315), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n292), .A2(KEYINPUT72), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT72), .B1(new_n292), .B2(new_n316), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT17), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n292), .A2(new_n316), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(KEYINPUT17), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT18), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n315), .A2(new_n288), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n291), .B1(new_n324), .B2(new_n309), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n270), .A2(new_n277), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G169), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n326), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n323), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n316), .A2(new_n290), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(new_n329), .A3(KEYINPUT18), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n319), .A2(new_n322), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G238), .A2(G1698), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n301), .B(new_n335), .C1(new_n274), .C2(G1698), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n336), .B(new_n269), .C1(G107), .C2(new_n301), .ZN(new_n337));
  INV_X1    g0137(.A(new_n255), .ZN(new_n338));
  INV_X1    g0138(.A(G244), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n273), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(G179), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(new_n340), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT15), .B(G87), .Z(new_n344));
  NOR2_X1   g0144(.A1(new_n256), .A2(G20), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n297), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n346), .B1(new_n283), .B2(new_n205), .C1(new_n282), .C2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n285), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n348), .A2(new_n288), .B1(new_n205), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n289), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n205), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n334), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G97), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G226), .A2(G1698), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n274), .B2(G1698), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n358), .B2(new_n301), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n359), .A2(new_n268), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT13), .ZN(new_n361));
  INV_X1    g0161(.A(new_n273), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G238), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n360), .A2(new_n361), .A3(new_n363), .A4(new_n338), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n363), .B(new_n338), .C1(new_n268), .C2(new_n359), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT13), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT69), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n365), .A2(KEYINPUT69), .A3(KEYINPUT13), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n328), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n364), .A2(new_n366), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(G169), .ZN(new_n373));
  AOI211_X1 g0173(.A(KEYINPUT14), .B(new_n342), .C1(new_n364), .C2(new_n366), .ZN(new_n374));
  OR3_X1    g0174(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n347), .A2(new_n202), .B1(new_n283), .B2(G68), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n256), .A2(new_n205), .A3(G20), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n288), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  XOR2_X1   g0178(.A(new_n378), .B(KEYINPUT11), .Z(new_n379));
  NOR2_X1   g0179(.A1(new_n351), .A2(new_n294), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n349), .A2(new_n294), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT12), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n381), .B(new_n382), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n379), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n375), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G190), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n368), .B2(new_n369), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n279), .B1(new_n364), .B2(new_n366), .ZN(new_n388));
  OR3_X1    g0188(.A1(new_n387), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n259), .A2(G222), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n301), .B(new_n391), .C1(new_n258), .C2(new_n259), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n392), .B(new_n269), .C1(G77), .C2(new_n301), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n362), .A2(G226), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n338), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G200), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n281), .A2(new_n345), .B1(G150), .B2(new_n297), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n204), .B2(new_n283), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n288), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n349), .A2(new_n202), .ZN(new_n400));
  OR3_X1    g0200(.A1(new_n284), .A2(KEYINPUT68), .A3(new_n202), .ZN(new_n401));
  INV_X1    g0201(.A(new_n288), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT68), .B1(new_n284), .B2(new_n202), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n285), .A4(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n399), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT9), .ZN(new_n406));
  OAI221_X1 g0206(.A(new_n396), .B1(new_n386), .B2(new_n395), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n406), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT10), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n399), .A2(new_n400), .A3(new_n404), .ZN(new_n411));
  INV_X1    g0211(.A(new_n395), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n411), .A2(KEYINPUT9), .B1(G190), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT10), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(new_n408), .A4(new_n396), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n395), .A2(new_n342), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n405), .B(new_n417), .C1(G179), .C2(new_n395), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n340), .A2(G200), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n340), .A2(new_n386), .ZN(new_n421));
  OR3_X1    g0221(.A1(new_n352), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NOR4_X1   g0223(.A1(new_n354), .A2(new_n390), .A3(new_n419), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n257), .A2(new_n262), .A3(G244), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT4), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n425), .A2(new_n426), .B1(G33), .B2(G283), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n301), .A2(KEYINPUT4), .A3(G244), .A4(new_n259), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n301), .B2(G250), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n427), .B(new_n428), .C1(new_n259), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n269), .ZN(new_n431));
  OR2_X1    g0231(.A1(KEYINPUT67), .A2(G41), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT5), .ZN(new_n433));
  NAND2_X1  g0233(.A1(KEYINPUT67), .A2(G41), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G41), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT5), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n254), .A2(G1), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n435), .A2(G274), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n269), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G257), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n431), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G200), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT73), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n297), .A2(G77), .ZN(new_n447));
  INV_X1    g0247(.A(G107), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(KEYINPUT6), .A3(G97), .ZN(new_n449));
  INV_X1    g0249(.A(G97), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(new_n448), .ZN(new_n451));
  NOR2_X1   g0251(.A1(G97), .A2(G107), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n449), .B1(new_n453), .B2(KEYINPUT6), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G20), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n311), .A2(new_n313), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n447), .B(new_n455), .C1(new_n456), .C2(new_n448), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n288), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n285), .A2(G97), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n251), .A2(G33), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n402), .A2(new_n285), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G97), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n458), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n430), .A2(new_n269), .B1(new_n441), .B2(G257), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(G190), .A3(new_n439), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n443), .A2(KEYINPUT73), .A3(G200), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n446), .A2(new_n464), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n458), .A2(new_n460), .A3(new_n463), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n443), .A2(new_n342), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n465), .A2(new_n328), .A3(new_n439), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n230), .A2(KEYINPUT79), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n474), .A2(new_n257), .A3(new_n262), .A4(new_n283), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT22), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT22), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n301), .A2(new_n477), .A3(new_n283), .A4(new_n474), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n283), .A2(G33), .A3(G116), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n283), .A2(G107), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n481), .B(KEYINPUT23), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n479), .A2(KEYINPUT80), .A3(new_n480), .A4(new_n482), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(KEYINPUT24), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n483), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n288), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n349), .A2(KEYINPUT25), .A3(new_n448), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT25), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n285), .B2(G107), .ZN(new_n493));
  AOI22_X1  g0293(.A1(G107), .A2(new_n462), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n257), .A2(new_n262), .A3(G250), .A4(new_n259), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n257), .A2(new_n262), .A3(G257), .A4(G1698), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G294), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n269), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(G264), .A3(new_n268), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n501), .A3(new_n439), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n279), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(G190), .B2(new_n502), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n490), .A2(new_n494), .A3(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(G274), .A2(new_n440), .B1(new_n498), .B2(new_n269), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n342), .B1(new_n506), .B2(new_n501), .ZN(new_n507));
  AND4_X1   g0307(.A1(G179), .A2(new_n499), .A3(new_n501), .A4(new_n439), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT81), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n502), .A2(G169), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT81), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n510), .B(new_n511), .C1(new_n328), .C2(new_n502), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n490), .A2(new_n494), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT82), .B1(new_n505), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n490), .A2(new_n494), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n509), .A2(new_n512), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT82), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n490), .A2(new_n494), .A3(new_n504), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n473), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n257), .A2(new_n262), .A3(G257), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(new_n259), .B1(G303), .B2(new_n312), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT76), .ZN(new_n524));
  AND2_X1   g0324(.A1(G264), .A2(G1698), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n257), .A2(new_n262), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT75), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT75), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n257), .A2(new_n262), .A3(new_n525), .A4(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n523), .A2(new_n524), .A3(new_n527), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n312), .A2(G303), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n257), .A2(new_n262), .A3(G257), .A4(new_n259), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n527), .A2(new_n531), .A3(new_n532), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT76), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(new_n534), .A3(new_n269), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n441), .A2(G270), .B1(G274), .B2(new_n440), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n462), .A2(G116), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n349), .A2(new_n221), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n221), .A2(G20), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n288), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT77), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT77), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n288), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(G20), .B1(G33), .B2(G283), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(G33), .B2(new_n450), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT20), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n288), .A2(new_n543), .A3(new_n540), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n543), .B1(new_n288), .B2(new_n540), .ZN(new_n550));
  OAI211_X1 g0350(.A(KEYINPUT20), .B(new_n547), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n538), .B(new_n539), .C1(new_n548), .C2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n537), .A2(new_n553), .A3(KEYINPUT21), .A4(G169), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n553), .A2(G179), .A3(new_n536), .A4(new_n535), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n537), .A2(G200), .ZN(new_n557));
  INV_X1    g0357(.A(new_n553), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n386), .C2(new_n537), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT78), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n342), .B1(new_n535), .B2(new_n536), .ZN(new_n561));
  AOI211_X1 g0361(.A(new_n560), .B(KEYINPUT21), .C1(new_n561), .C2(new_n553), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n537), .A2(G169), .A3(new_n553), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT21), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT78), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n556), .B(new_n559), .C1(new_n562), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n452), .A2(new_n230), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n567), .B(KEYINPUT19), .C1(new_n356), .C2(G20), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n257), .A2(new_n262), .A3(new_n283), .A4(G68), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT19), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n355), .B2(G20), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n288), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n462), .A2(new_n344), .ZN(new_n574));
  INV_X1    g0374(.A(new_n344), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n349), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT74), .ZN(new_n578));
  INV_X1    g0378(.A(G274), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n438), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n580), .B(new_n268), .C1(G250), .C2(new_n438), .ZN(new_n581));
  NOR2_X1   g0381(.A1(G238), .A2(G1698), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n339), .B2(G1698), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(new_n301), .B1(G33), .B2(G116), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n581), .B1(new_n584), .B2(new_n268), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G169), .ZN(new_n586));
  OAI211_X1 g0386(.A(G179), .B(new_n581), .C1(new_n584), .C2(new_n268), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n572), .A2(new_n288), .B1(new_n349), .B2(new_n575), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT74), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n590), .A3(new_n574), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n578), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n585), .A2(G200), .ZN(new_n593));
  OAI211_X1 g0393(.A(G190), .B(new_n581), .C1(new_n584), .C2(new_n268), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n462), .A2(G87), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n593), .A2(new_n589), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n566), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n424), .A2(new_n521), .A3(new_n598), .ZN(G372));
  NOR3_X1   g0399(.A1(new_n387), .A2(new_n384), .A3(new_n388), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n385), .B1(new_n600), .B2(new_n353), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n319), .A2(new_n322), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n331), .A2(new_n333), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n416), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n418), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n424), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n592), .A2(new_n596), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT26), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT26), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n472), .A2(new_n597), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n592), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n554), .A2(new_n555), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n563), .A2(new_n564), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n560), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n563), .A2(KEYINPUT78), .A3(new_n564), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n515), .B1(new_n507), .B2(new_n508), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n468), .A2(new_n519), .A3(new_n472), .A4(new_n596), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n615), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n608), .B1(new_n609), .B2(new_n625), .ZN(G369));
  INV_X1    g0426(.A(G13), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(G20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n251), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT83), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT84), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n634));
  INV_X1    g0434(.A(G213), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(G343), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n621), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n639), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n517), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n514), .A2(new_n520), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n639), .A2(new_n515), .ZN(new_n645));
  OAI211_X1 g0445(.A(KEYINPUT85), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT85), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n514), .A2(new_n520), .B1(new_n515), .B2(new_n639), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n642), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n620), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n641), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n640), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G330), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n651), .A2(new_n553), .A3(new_n639), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n620), .B(new_n559), .C1(new_n558), .C2(new_n641), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n654), .A2(new_n659), .ZN(G399));
  INV_X1    g0460(.A(new_n253), .ZN(new_n661));
  INV_X1    g0461(.A(new_n209), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n567), .A2(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n218), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n623), .B1(new_n620), .B2(new_n517), .ZN(new_n669));
  OAI211_X1 g0469(.A(KEYINPUT29), .B(new_n641), .C1(new_n669), .C2(new_n615), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT88), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT86), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n625), .B2(new_n639), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT29), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n623), .B1(new_n620), .B2(new_n621), .ZN(new_n675));
  OAI211_X1 g0475(.A(KEYINPUT86), .B(new_n641), .C1(new_n675), .C2(new_n615), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT87), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT87), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n673), .A2(new_n679), .A3(new_n674), .A4(new_n676), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n671), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n521), .A2(new_n598), .A3(new_n641), .ZN(new_n682));
  INV_X1    g0482(.A(new_n537), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n502), .A2(new_n587), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(KEYINPUT30), .A3(new_n465), .A4(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n684), .A2(new_n465), .A3(new_n536), .A4(new_n535), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n585), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n537), .A2(new_n328), .A3(new_n443), .A4(new_n502), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n685), .B(new_n688), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n639), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT31), .B1(new_n691), .B2(new_n639), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n655), .B1(new_n682), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n681), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n668), .B1(new_n696), .B2(G1), .ZN(G364));
  AOI21_X1  g0497(.A(new_n212), .B1(G20), .B2(new_n342), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n283), .A2(G179), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n386), .A3(G200), .ZN(new_n700));
  INV_X1    g0500(.A(G283), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT89), .B1(new_n283), .B2(new_n328), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT89), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(G20), .A3(G179), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n386), .A2(G200), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G322), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n699), .A2(G190), .A3(G200), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT91), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G303), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n312), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT93), .ZN(new_n721));
  INV_X1    g0521(.A(G294), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n283), .B1(new_n708), .B2(new_n328), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n720), .A2(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n713), .B(new_n724), .C1(new_n721), .C2(new_n720), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT90), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n707), .B2(new_n279), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n706), .A2(KEYINPUT90), .A3(G200), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n386), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(KEYINPUT33), .B(G317), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n727), .A2(G190), .A3(new_n728), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT92), .Z(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G326), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G190), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n699), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT94), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G329), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n725), .A2(new_n732), .A3(new_n735), .A4(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n736), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n707), .A2(new_n742), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n702), .B(new_n741), .C1(G311), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n723), .A2(new_n450), .ZN(new_n745));
  INV_X1    g0545(.A(G159), .ZN(new_n746));
  OR3_X1    g0546(.A1(new_n737), .A2(KEYINPUT32), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(KEYINPUT32), .B1(new_n737), .B2(new_n746), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n747), .B(new_n748), .C1(new_n448), .C2(new_n700), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n745), .B(new_n749), .C1(G77), .C2(new_n743), .ZN(new_n750));
  INV_X1    g0550(.A(new_n733), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G50), .A2(new_n751), .B1(new_n730), .B2(G68), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n750), .B(new_n752), .C1(new_n293), .C2(new_n711), .ZN(new_n753));
  INV_X1    g0553(.A(new_n718), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n312), .B(new_n753), .C1(G87), .C2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n698), .B1(new_n744), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n301), .A2(G355), .A3(new_n209), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n246), .A2(new_n254), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n662), .A2(new_n301), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(new_n218), .B2(G45), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n757), .B1(G116), .B2(new_n209), .C1(new_n758), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n698), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n656), .A2(new_n657), .A3(new_n764), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n628), .A2(G45), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n664), .A2(G1), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n756), .A2(new_n766), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n658), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n656), .A2(new_n655), .A3(new_n657), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n772), .A2(new_n769), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n771), .A2(new_n774), .ZN(G396));
  INV_X1    g0575(.A(new_n698), .ZN(new_n776));
  INV_X1    g0576(.A(G132), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n301), .B1(new_n738), .B2(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G143), .A2(new_n710), .B1(new_n743), .B2(G159), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G137), .A2(new_n751), .B1(new_n730), .B2(G150), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT96), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT34), .Z(new_n785));
  INV_X1    g0585(.A(new_n700), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n778), .B(new_n785), .C1(G68), .C2(new_n786), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n787), .B1(new_n202), .B2(new_n718), .C1(new_n293), .C2(new_n723), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n729), .A2(KEYINPUT95), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n729), .A2(KEYINPUT95), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n792), .A2(G283), .B1(G294), .B2(new_n710), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n786), .A2(G87), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n733), .A2(new_n719), .ZN(new_n795));
  INV_X1    g0595(.A(new_n743), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n796), .A2(new_n221), .B1(new_n718), .B2(new_n448), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n738), .A2(new_n798), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n795), .A2(new_n797), .A3(new_n745), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n793), .A2(new_n312), .A3(new_n794), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n776), .B1(new_n788), .B2(new_n801), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n698), .A2(G77), .A3(new_n762), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n353), .A2(new_n639), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n639), .A2(new_n352), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n422), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n804), .B1(new_n806), .B2(new_n353), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n763), .ZN(new_n808));
  NOR4_X1   g0608(.A1(new_n802), .A2(new_n769), .A3(new_n803), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n806), .A2(new_n353), .ZN(new_n810));
  INV_X1    g0610(.A(new_n804), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n673), .A2(new_n676), .A3(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n641), .B(new_n807), .C1(new_n675), .C2(new_n615), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(new_n695), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n816), .A2(new_n769), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n809), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G384));
  NAND2_X1  g0619(.A1(new_n639), .A2(new_n384), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n821));
  INV_X1    g0621(.A(new_n384), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n389), .B(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n384), .B(new_n639), .C1(new_n375), .C2(new_n600), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n804), .B(KEYINPUT97), .Z(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n814), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n300), .B1(new_n308), .B2(new_n294), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n829), .A2(new_n310), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n309), .A2(new_n288), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n290), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT98), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(KEYINPUT98), .B(new_n290), .C1(new_n830), .C2(new_n831), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n330), .A2(new_n637), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT72), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n309), .A2(new_n288), .A3(new_n315), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n326), .A2(G200), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n840), .B(new_n290), .C1(new_n386), .C2(new_n326), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n838), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n292), .A2(new_n316), .A3(KEYINPUT72), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n837), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n332), .A2(new_n329), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n633), .A2(new_n636), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT37), .B1(new_n848), .B2(new_n332), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n844), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT99), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n834), .A2(new_n848), .A3(new_n835), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n334), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT17), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n842), .B2(new_n843), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n604), .B1(new_n856), .B2(new_n321), .ZN(new_n857));
  INV_X1    g0657(.A(new_n853), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT99), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(KEYINPUT38), .B(new_n851), .C1(new_n854), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n852), .B1(new_n334), .B2(new_n853), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n857), .A2(KEYINPUT99), .A3(new_n858), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n864), .B2(new_n851), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n828), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT100), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n604), .A2(new_n848), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n851), .B1(new_n854), .B2(new_n859), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(KEYINPUT39), .A3(new_n860), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n847), .B1(new_n317), .B2(new_n318), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n848), .A2(new_n332), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT101), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n847), .A3(new_n320), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT101), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n844), .A2(new_n849), .A3(new_n882), .A4(new_n847), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n879), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n334), .A2(new_n876), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n872), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n860), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n385), .A2(new_n639), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n874), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n870), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n867), .B1(new_n866), .B2(new_n869), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n607), .B1(new_n681), .B2(new_n424), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n894), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n825), .A2(new_n807), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n682), .B2(new_n694), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n861), .B2(new_n865), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n887), .A2(KEYINPUT40), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n682), .A2(new_n694), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n424), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n903), .B(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n655), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n896), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n251), .B2(new_n628), .ZN(new_n909));
  OAI211_X1 g0709(.A(G20), .B(new_n213), .C1(new_n454), .C2(KEYINPUT35), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n221), .B(new_n910), .C1(KEYINPUT35), .C2(new_n454), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT36), .Z(new_n912));
  OAI21_X1  g0712(.A(G77), .B1(new_n293), .B2(new_n294), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n218), .A2(new_n913), .B1(G50), .B2(new_n294), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(G1), .A3(new_n627), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n909), .A2(new_n912), .A3(new_n915), .ZN(G367));
  NAND2_X1  g0716(.A1(new_n650), .A2(new_n653), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n468), .B(new_n472), .C1(new_n641), .C2(new_n464), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n610), .A2(new_n639), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR3_X1    g0720(.A1(new_n917), .A2(KEYINPUT42), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT42), .B1(new_n917), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n472), .B1(new_n918), .B2(new_n517), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT102), .Z(new_n924));
  OAI211_X1 g0724(.A(new_n921), .B(new_n922), .C1(new_n639), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n589), .A2(new_n595), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n639), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n927), .A2(new_n592), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n611), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n925), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n659), .ZN(new_n933));
  INV_X1    g0733(.A(new_n920), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n925), .A2(new_n935), .A3(new_n931), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n938), .B1(new_n937), .B2(new_n939), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n663), .B(KEYINPUT41), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n652), .B1(new_n646), .B2(new_n649), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n920), .B1(new_n945), .B2(new_n640), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT44), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n640), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n917), .A2(new_n949), .A3(new_n934), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT103), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT103), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n654), .A2(new_n952), .A3(new_n934), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n951), .A2(KEYINPUT45), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT45), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n952), .B1(new_n654), .B2(new_n934), .ZN(new_n956));
  NOR4_X1   g0756(.A1(new_n945), .A2(KEYINPUT103), .A3(new_n640), .A4(new_n920), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n948), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n933), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n948), .A2(new_n954), .A3(new_n958), .A4(new_n659), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n658), .A2(new_n653), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(new_n650), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n696), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n960), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n944), .B1(new_n965), .B2(new_n696), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n768), .A2(G1), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n942), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n700), .A2(new_n450), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n792), .A2(G294), .B1(new_n734), .B2(G311), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT46), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n754), .A2(G116), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n970), .B1(new_n971), .B2(new_n972), .C1(new_n448), .C2(new_n723), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT104), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n972), .B2(new_n971), .ZN(new_n975));
  AOI211_X1 g0775(.A(KEYINPUT104), .B(KEYINPUT46), .C1(new_n754), .C2(G116), .ZN(new_n976));
  OR4_X1    g0776(.A1(new_n969), .A2(new_n973), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n301), .B(new_n977), .C1(G303), .C2(new_n710), .ZN(new_n978));
  INV_X1    g0778(.A(G317), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n978), .B1(new_n701), .B2(new_n796), .C1(new_n979), .C2(new_n737), .ZN(new_n980));
  INV_X1    g0780(.A(new_n723), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n743), .A2(G50), .B1(G68), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(G137), .ZN(new_n983));
  INV_X1    g0783(.A(G150), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n982), .B1(new_n983), .B2(new_n737), .C1(new_n984), .C2(new_n711), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n301), .B1(new_n718), .B2(new_n293), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n700), .A2(new_n205), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n734), .ZN(new_n989));
  INV_X1    g0789(.A(G143), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n988), .B1(new_n746), .B2(new_n791), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n980), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n698), .ZN(new_n994));
  INV_X1    g0794(.A(new_n759), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n765), .B1(new_n209), .B2(new_n575), .C1(new_n242), .C2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n928), .A2(new_n764), .A3(new_n929), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n770), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n968), .A2(new_n998), .ZN(G387));
  NOR2_X1   g0799(.A1(new_n964), .A2(new_n664), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n696), .B2(new_n963), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n963), .A2(new_n967), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT105), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G303), .A2(new_n743), .B1(new_n710), .B2(G317), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT109), .Z(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n798), .B2(new_n791), .C1(new_n989), .C2(new_n712), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT48), .Z(new_n1007));
  OAI22_X1  g0807(.A1(new_n718), .A2(new_n722), .B1(new_n701), .B2(new_n723), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1008), .A2(KEYINPUT108), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(KEYINPUT108), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT49), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n786), .A2(G116), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n737), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(G326), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n312), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1011), .A2(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n981), .A2(new_n344), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n711), .B2(new_n202), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT106), .Z(new_n1020));
  NOR2_X1   g0820(.A1(new_n1020), .A2(new_n969), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n754), .A2(G77), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n729), .A2(new_n282), .B1(new_n294), .B2(new_n796), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT107), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n301), .B1(new_n984), .B2(new_n737), .C1(new_n733), .C2(new_n746), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1016), .A2(new_n1017), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n759), .B1(new_n239), .B2(new_n254), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n301), .A2(new_n209), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n665), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n281), .A2(new_n202), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT50), .Z(new_n1032));
  NAND2_X1  g0832(.A1(G68), .A2(G77), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1032), .A2(new_n254), .A3(new_n1033), .A4(new_n665), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(G107), .B2(new_n209), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1027), .A2(new_n698), .B1(new_n765), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n764), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1037), .B(new_n770), .C1(new_n650), .C2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1001), .A2(new_n1003), .A3(new_n1039), .ZN(G393));
  NAND2_X1  g0840(.A1(new_n960), .A2(new_n961), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n733), .A2(new_n979), .B1(new_n798), .B2(new_n711), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT111), .Z(new_n1044));
  NOR2_X1   g0844(.A1(new_n1044), .A2(KEYINPUT52), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(KEYINPUT52), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n719), .B2(new_n791), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1045), .B(new_n1047), .C1(G116), .C2(new_n981), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n301), .B1(new_n1014), .B2(G322), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n448), .B2(new_n700), .C1(new_n718), .C2(new_n701), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT112), .Z(new_n1051));
  OAI211_X1 g0851(.A(new_n1048), .B(new_n1051), .C1(new_n722), .C2(new_n796), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT113), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n733), .A2(new_n984), .B1(new_n746), .B2(new_n711), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT51), .Z(new_n1055));
  OAI211_X1 g0855(.A(new_n794), .B(new_n301), .C1(new_n990), .C2(new_n737), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n792), .A2(G50), .B1(G77), .B2(new_n981), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n282), .C2(new_n796), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G68), .B2(new_n754), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n698), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n765), .B1(new_n450), .B2(new_n209), .C1(new_n249), .C2(new_n995), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT110), .Z(new_n1063));
  AOI211_X1 g0863(.A(new_n769), .B(new_n1063), .C1(new_n920), .C2(new_n764), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1042), .A2(new_n967), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n964), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1041), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n663), .A3(new_n965), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1065), .A2(new_n1068), .ZN(G390));
  AND2_X1   g0869(.A1(new_n874), .A2(new_n889), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1070), .A2(new_n763), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G77), .A2(new_n981), .B1(new_n786), .B2(G68), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n711), .B2(new_n221), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n312), .B1(new_n796), .B2(new_n450), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n792), .B2(G107), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n230), .B2(new_n718), .C1(new_n722), .C2(new_n738), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1073), .B(new_n1076), .C1(G283), .C2(new_n751), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n792), .A2(G137), .ZN(new_n1078));
  XOR2_X1   g0878(.A(KEYINPUT54), .B(G143), .Z(new_n1079));
  NAND2_X1  g0879(.A1(new_n743), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n312), .B1(new_n981), .B2(G159), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G132), .B2(new_n710), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n751), .A2(G128), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n739), .A2(G125), .B1(G50), .B2(new_n786), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n718), .A2(new_n984), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT53), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1077), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT115), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n698), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n698), .A2(new_n762), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n282), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1071), .A2(new_n770), .A3(new_n1091), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n695), .A2(new_n807), .A3(new_n825), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n890), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n641), .B(new_n810), .C1(new_n669), .C2(new_n615), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1097), .A2(new_n811), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n887), .B(new_n1096), .C1(new_n1098), .C2(new_n826), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n828), .A2(new_n890), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1095), .B(new_n1099), .C1(new_n1070), .C2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1095), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1100), .B1(new_n889), .B2(new_n874), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1099), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1105), .A3(new_n967), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT116), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1094), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(new_n1094), .B2(new_n1106), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n904), .A2(G330), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n826), .B1(new_n1111), .B2(new_n812), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n1095), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n814), .A2(new_n827), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n1098), .A3(new_n1095), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n424), .A2(G330), .A3(new_n904), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n895), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n663), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT114), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT114), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1124), .B(new_n663), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1110), .A2(new_n1126), .ZN(G378));
  AOI21_X1  g0927(.A(new_n812), .B1(new_n823), .B2(new_n824), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n904), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n873), .B2(new_n860), .ZN(new_n1130));
  OAI211_X1 g0930(.A(G330), .B(new_n902), .C1(new_n1130), .C2(KEYINPUT40), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n637), .A2(new_n411), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n419), .A2(KEYINPUT119), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT119), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n416), .A2(new_n1135), .A3(new_n418), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1133), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1134), .A2(new_n1136), .A3(new_n1133), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1139), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1131), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n901), .A2(G330), .A3(new_n902), .A4(new_n1143), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n866), .A2(new_n869), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT100), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n891), .A3(new_n870), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT120), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n894), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(KEYINPUT121), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT121), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1152), .A2(new_n894), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1151), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1150), .A2(new_n1146), .A3(new_n1145), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT120), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1152), .A2(new_n1155), .A3(new_n894), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1155), .B1(new_n1152), .B2(new_n894), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n895), .B(new_n1118), .C1(new_n1120), .C2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1157), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT57), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1165), .A2(new_n1169), .A3(KEYINPUT57), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n663), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1157), .A2(new_n1163), .A3(new_n967), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1143), .A2(new_n762), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n661), .A2(new_n301), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1022), .A2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1177), .A2(KEYINPUT118), .B1(new_n344), .B2(new_n743), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(KEYINPUT118), .B2(new_n1177), .C1(new_n448), .C2(new_n711), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n738), .A2(new_n701), .B1(new_n294), .B2(new_n723), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n700), .A2(new_n293), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n450), .B2(new_n729), .C1(new_n221), .C2(new_n733), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT58), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G50), .B(new_n1176), .C1(new_n256), .C2(new_n436), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT117), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1186), .A2(KEYINPUT117), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n751), .A2(G125), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n743), .A2(G137), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n754), .A2(new_n1079), .B1(new_n710), .B2(G128), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n777), .B2(new_n729), .C1(new_n984), .C2(new_n723), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT59), .Z(new_n1194));
  NAND2_X1  g0994(.A1(new_n1014), .A2(G124), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G33), .B(G41), .C1(new_n786), .C2(G159), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1185), .A2(new_n1187), .A3(new_n1188), .A4(new_n1197), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n698), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1092), .A2(new_n202), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1175), .A2(new_n1200), .A3(new_n770), .A4(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1174), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1173), .A2(new_n1204), .ZN(G375));
  NAND2_X1  g1005(.A1(new_n792), .A2(new_n1079), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n754), .A2(G159), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n301), .B1(new_n711), .B2(new_n983), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n751), .B2(G132), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n796), .A2(new_n984), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1181), .B(new_n1210), .C1(G128), .C2(new_n739), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1206), .A2(new_n1207), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G50), .B2(new_n981), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n751), .A2(G294), .B1(G107), .B2(new_n743), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n791), .B2(new_n221), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT124), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n301), .B(new_n987), .C1(new_n710), .C2(G283), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1018), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G303), .B2(new_n739), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n754), .A2(G97), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1213), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1221), .A2(new_n776), .B1(new_n763), .B2(new_n825), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n769), .B1(new_n294), .B2(new_n1092), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT123), .Z(new_n1224));
  NOR2_X1   g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1117), .B2(new_n967), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n678), .A2(new_n680), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n671), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n424), .A3(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n608), .A3(new_n1118), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1230), .A2(new_n1164), .A3(KEYINPUT122), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT122), .B1(new_n1230), .B2(new_n1164), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1119), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1226), .B1(new_n1233), .B2(new_n944), .ZN(G381));
  AND4_X1   g1034(.A1(new_n968), .A2(new_n998), .A3(new_n1065), .A4(new_n1068), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(G381), .A2(G384), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(G393), .A2(G396), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT125), .Z(new_n1239));
  AND3_X1   g1039(.A1(new_n1126), .A2(new_n1106), .A3(new_n1094), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1173), .A2(new_n1204), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(G407));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n638), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G407), .A2(G213), .A3(new_n1243), .ZN(G409));
  NOR2_X1   g1044(.A1(new_n635), .A2(G343), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1119), .A2(KEYINPUT60), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1230), .A2(new_n1164), .A3(KEYINPUT60), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n663), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1226), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n818), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(G384), .A3(new_n1226), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1171), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1110), .A2(new_n1126), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1256), .A2(new_n1257), .A3(new_n1203), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1157), .A2(new_n1163), .A3(new_n943), .A4(new_n1165), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1169), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1153), .A2(new_n1158), .A3(KEYINPUT126), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n967), .A3(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1259), .A2(new_n1202), .A3(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1264), .A2(new_n1240), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1246), .B(new_n1255), .C1(new_n1258), .C2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT62), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1246), .B1(new_n1258), .B2(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1245), .A2(G2897), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1250), .A2(G384), .A3(new_n1226), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G384), .B1(new_n1250), .B2(new_n1226), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1270), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1252), .A2(new_n1253), .A3(new_n1269), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1268), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1173), .A2(G378), .A3(new_n1204), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1264), .A2(new_n1240), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT62), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n1246), .A4(new_n1255), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1267), .A2(new_n1277), .A3(new_n1278), .A4(new_n1283), .ZN(new_n1284));
  XOR2_X1   g1084(.A(G393), .B(G396), .Z(new_n1285));
  AOI22_X1  g1085(.A1(new_n968), .A2(new_n998), .B1(new_n1068), .B2(new_n1065), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1285), .B1(new_n1235), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G387), .A2(G390), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n968), .A2(new_n998), .A3(new_n1065), .A4(new_n1068), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(G393), .B(G396), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1284), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1275), .B1(new_n1281), .B2(new_n1246), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1266), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  AOI211_X1 g1096(.A(new_n1245), .B(new_n1254), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1292), .B1(new_n1297), .B2(KEYINPUT63), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1298), .A3(new_n1278), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1293), .A2(new_n1299), .ZN(G405));
  OAI21_X1  g1100(.A(new_n1240), .B1(new_n1256), .B2(new_n1203), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1301), .B1(new_n1258), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(G375), .A2(KEYINPUT127), .A3(new_n1240), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1292), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1292), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1254), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(new_n1287), .A3(new_n1291), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1292), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1255), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1307), .A2(new_n1311), .ZN(G402));
endmodule


