

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(n818), .A2(n932), .ZN(n519) );
  XNOR2_X1 U552 ( .A(KEYINPUT28), .B(KEYINPUT96), .ZN(n707) );
  XNOR2_X1 U553 ( .A(n708), .B(n707), .ZN(n731) );
  NOR2_X1 U554 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U555 ( .A1(n699), .A2(n698), .ZN(n745) );
  NAND2_X1 U556 ( .A1(G8), .A2(n745), .ZN(n788) );
  NOR2_X1 U557 ( .A1(n803), .A2(n519), .ZN(n804) );
  AND2_X1 U558 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U559 ( .A1(G651), .A2(n609), .ZN(n636) );
  AND2_X1 U560 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U561 ( .A(G132), .ZN(G219) );
  INV_X1 U562 ( .A(G120), .ZN(G236) );
  INV_X1 U563 ( .A(G69), .ZN(G235) );
  INV_X1 U564 ( .A(G108), .ZN(G238) );
  INV_X1 U565 ( .A(G2104), .ZN(n524) );
  NOR2_X1 U566 ( .A1(G2105), .A2(n524), .ZN(n885) );
  NAND2_X1 U567 ( .A1(G102), .A2(n885), .ZN(n523) );
  XNOR2_X1 U568 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n521) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XNOR2_X2 U570 ( .A(n521), .B(n520), .ZN(n883) );
  NAND2_X1 U571 ( .A1(G138), .A2(n883), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n523), .A2(n522), .ZN(n529) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n879) );
  NAND2_X1 U574 ( .A1(G114), .A2(n879), .ZN(n527) );
  NAND2_X1 U575 ( .A1(n524), .A2(G2105), .ZN(n525) );
  XNOR2_X2 U576 ( .A(n525), .B(KEYINPUT65), .ZN(n880) );
  NAND2_X1 U577 ( .A1(G126), .A2(n880), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U580 ( .A(KEYINPUT91), .B(n530), .Z(G164) );
  NOR2_X1 U581 ( .A1(G543), .A2(G651), .ZN(n639) );
  NAND2_X1 U582 ( .A1(n639), .A2(G89), .ZN(n531) );
  XNOR2_X1 U583 ( .A(n531), .B(KEYINPUT4), .ZN(n533) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n609) );
  INV_X1 U585 ( .A(G651), .ZN(n535) );
  NOR2_X1 U586 ( .A1(n609), .A2(n535), .ZN(n635) );
  NAND2_X1 U587 ( .A1(G76), .A2(n635), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U589 ( .A(KEYINPUT5), .B(n534), .ZN(n542) );
  NOR2_X1 U590 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n536), .Z(n634) );
  NAND2_X1 U592 ( .A1(n634), .A2(G63), .ZN(n537) );
  XOR2_X1 U593 ( .A(KEYINPUT77), .B(n537), .Z(n539) );
  NAND2_X1 U594 ( .A1(n636), .A2(G51), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U596 ( .A(KEYINPUT6), .B(n540), .Z(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U598 ( .A(KEYINPUT7), .B(n543), .ZN(G168) );
  XOR2_X1 U599 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U600 ( .A1(G7), .A2(G661), .ZN(n544) );
  XNOR2_X1 U601 ( .A(n544), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U602 ( .A(G223), .ZN(n822) );
  NAND2_X1 U603 ( .A1(n822), .A2(G567), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT11), .B(n545), .Z(G234) );
  NAND2_X1 U605 ( .A1(n639), .A2(G81), .ZN(n546) );
  XNOR2_X1 U606 ( .A(n546), .B(KEYINPUT12), .ZN(n548) );
  NAND2_X1 U607 ( .A1(G68), .A2(n635), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U609 ( .A(KEYINPUT13), .B(n549), .Z(n553) );
  NAND2_X1 U610 ( .A1(G56), .A2(n634), .ZN(n550) );
  XNOR2_X1 U611 ( .A(n550), .B(KEYINPUT14), .ZN(n551) );
  XNOR2_X1 U612 ( .A(n551), .B(KEYINPUT73), .ZN(n552) );
  NOR2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U614 ( .A(n554), .B(KEYINPUT74), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G43), .A2(n636), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n918) );
  INV_X1 U617 ( .A(G860), .ZN(n585) );
  OR2_X1 U618 ( .A1(n918), .A2(n585), .ZN(G153) );
  NAND2_X1 U619 ( .A1(n635), .A2(G77), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT69), .B(n557), .Z(n559) );
  NAND2_X1 U621 ( .A1(n639), .A2(G90), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U623 ( .A(KEYINPUT9), .B(n560), .ZN(n564) );
  NAND2_X1 U624 ( .A1(n636), .A2(G52), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G64), .A2(n634), .ZN(n561) );
  AND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(G301) );
  NAND2_X1 U628 ( .A1(G92), .A2(n639), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G66), .A2(n634), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G79), .A2(n635), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G54), .A2(n636), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT75), .B(n569), .Z(n570) );
  NOR2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT15), .B(n572), .ZN(n919) );
  INV_X1 U637 ( .A(G868), .ZN(n653) );
  NAND2_X1 U638 ( .A1(n919), .A2(n653), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT76), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G868), .A2(G301), .ZN(n574) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(G284) );
  NAND2_X1 U642 ( .A1(G78), .A2(n635), .ZN(n577) );
  NAND2_X1 U643 ( .A1(G91), .A2(n639), .ZN(n576) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G53), .A2(n636), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G65), .A2(n634), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U649 ( .A(KEYINPUT70), .B(n582), .Z(n924) );
  XOR2_X1 U650 ( .A(n924), .B(KEYINPUT71), .Z(G299) );
  NOR2_X1 U651 ( .A1(G299), .A2(G868), .ZN(n584) );
  NOR2_X1 U652 ( .A1(G286), .A2(n653), .ZN(n583) );
  NOR2_X1 U653 ( .A1(n584), .A2(n583), .ZN(G297) );
  NAND2_X1 U654 ( .A1(n585), .A2(G559), .ZN(n586) );
  INV_X1 U655 ( .A(n919), .ZN(n651) );
  NAND2_X1 U656 ( .A1(n586), .A2(n651), .ZN(n587) );
  XNOR2_X1 U657 ( .A(n587), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U658 ( .A1(G868), .A2(n918), .ZN(n590) );
  NAND2_X1 U659 ( .A1(G868), .A2(n651), .ZN(n588) );
  NOR2_X1 U660 ( .A1(G559), .A2(n588), .ZN(n589) );
  NOR2_X1 U661 ( .A1(n590), .A2(n589), .ZN(G282) );
  NAND2_X1 U662 ( .A1(G123), .A2(n880), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n591), .B(KEYINPUT18), .ZN(n594) );
  NAND2_X1 U664 ( .A1(G99), .A2(n885), .ZN(n592) );
  XOR2_X1 U665 ( .A(KEYINPUT79), .B(n592), .Z(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n883), .A2(G135), .ZN(n595) );
  XNOR2_X1 U668 ( .A(n595), .B(KEYINPUT78), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G111), .A2(n879), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n996) );
  XNOR2_X1 U672 ( .A(G2096), .B(n996), .ZN(n601) );
  INV_X1 U673 ( .A(G2100), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(G156) );
  NAND2_X1 U675 ( .A1(G75), .A2(n635), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G88), .A2(n639), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U678 ( .A1(G62), .A2(n634), .ZN(n604) );
  XNOR2_X1 U679 ( .A(KEYINPUT85), .B(n604), .ZN(n605) );
  NOR2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n636), .A2(G50), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(G303) );
  INV_X1 U683 ( .A(G303), .ZN(G166) );
  NAND2_X1 U684 ( .A1(G74), .A2(G651), .ZN(n614) );
  NAND2_X1 U685 ( .A1(G49), .A2(n636), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G87), .A2(n609), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n634), .A2(n612), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n615), .B(KEYINPUT82), .ZN(G288) );
  NAND2_X1 U691 ( .A1(G72), .A2(n635), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G85), .A2(n639), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G60), .A2(n634), .ZN(n618) );
  XOR2_X1 U695 ( .A(KEYINPUT68), .B(n618), .Z(n619) );
  NOR2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n636), .A2(G47), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(G290) );
  NAND2_X1 U699 ( .A1(G73), .A2(n635), .ZN(n623) );
  XOR2_X1 U700 ( .A(KEYINPUT2), .B(n623), .Z(n624) );
  XNOR2_X1 U701 ( .A(n624), .B(KEYINPUT83), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G86), .A2(n639), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G48), .A2(n636), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G61), .A2(n634), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U708 ( .A(KEYINPUT84), .B(n631), .Z(G305) );
  XOR2_X1 U709 ( .A(G299), .B(KEYINPUT86), .Z(n633) );
  XNOR2_X1 U710 ( .A(G166), .B(KEYINPUT19), .ZN(n632) );
  XNOR2_X1 U711 ( .A(n633), .B(n632), .ZN(n649) );
  NAND2_X1 U712 ( .A1(G67), .A2(n634), .ZN(n644) );
  NAND2_X1 U713 ( .A1(G80), .A2(n635), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G55), .A2(n636), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n639), .A2(G93), .ZN(n640) );
  XOR2_X1 U717 ( .A(KEYINPUT80), .B(n640), .Z(n641) );
  NOR2_X1 U718 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n645), .B(KEYINPUT81), .ZN(n833) );
  XNOR2_X1 U721 ( .A(G288), .B(n833), .ZN(n647) );
  XNOR2_X1 U722 ( .A(G290), .B(G305), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n647), .B(n646), .ZN(n648) );
  XOR2_X1 U724 ( .A(n649), .B(n648), .Z(n650) );
  XNOR2_X1 U725 ( .A(n918), .B(n650), .ZN(n896) );
  NAND2_X1 U726 ( .A1(n651), .A2(G559), .ZN(n831) );
  XNOR2_X1 U727 ( .A(n896), .B(n831), .ZN(n652) );
  NOR2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n655) );
  NOR2_X1 U729 ( .A1(n833), .A2(G868), .ZN(n654) );
  NOR2_X1 U730 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U731 ( .A(KEYINPUT87), .B(n656), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2084), .A2(G2078), .ZN(n657) );
  XOR2_X1 U733 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n658), .ZN(n660) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(KEYINPUT88), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U737 ( .A1(G2072), .A2(n661), .ZN(G158) );
  XOR2_X1 U738 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U740 ( .A1(G235), .A2(G236), .ZN(n662) );
  XOR2_X1 U741 ( .A(KEYINPUT90), .B(n662), .Z(n663) );
  NOR2_X1 U742 ( .A1(G238), .A2(n663), .ZN(n664) );
  NAND2_X1 U743 ( .A1(G57), .A2(n664), .ZN(n829) );
  NAND2_X1 U744 ( .A1(n829), .A2(G567), .ZN(n670) );
  NOR2_X1 U745 ( .A1(G220), .A2(G219), .ZN(n665) );
  XNOR2_X1 U746 ( .A(KEYINPUT22), .B(n665), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n666), .A2(G96), .ZN(n667) );
  NOR2_X1 U748 ( .A1(n667), .A2(G218), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n668), .B(KEYINPUT89), .ZN(n830) );
  NAND2_X1 U750 ( .A1(n830), .A2(G2106), .ZN(n669) );
  NAND2_X1 U751 ( .A1(n670), .A2(n669), .ZN(n835) );
  NAND2_X1 U752 ( .A1(G661), .A2(G483), .ZN(n671) );
  NOR2_X1 U753 ( .A1(n835), .A2(n671), .ZN(n826) );
  NAND2_X1 U754 ( .A1(n826), .A2(G36), .ZN(G176) );
  XOR2_X1 U755 ( .A(KEYINPUT66), .B(KEYINPUT23), .Z(n673) );
  NAND2_X1 U756 ( .A1(G101), .A2(n885), .ZN(n672) );
  XNOR2_X1 U757 ( .A(n673), .B(n672), .ZN(n675) );
  NAND2_X1 U758 ( .A1(n883), .A2(G137), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U760 ( .A1(G113), .A2(n879), .ZN(n677) );
  NAND2_X1 U761 ( .A1(G125), .A2(n880), .ZN(n676) );
  NAND2_X1 U762 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U763 ( .A1(n679), .A2(n678), .ZN(G160) );
  INV_X1 U764 ( .A(G301), .ZN(G171) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n697) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n680) );
  XNOR2_X1 U767 ( .A(n680), .B(KEYINPUT64), .ZN(n698) );
  NOR2_X1 U768 ( .A1(n697), .A2(n698), .ZN(n818) );
  NAND2_X1 U769 ( .A1(G95), .A2(n885), .ZN(n682) );
  NAND2_X1 U770 ( .A1(G131), .A2(n883), .ZN(n681) );
  NAND2_X1 U771 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U772 ( .A1(G107), .A2(n879), .ZN(n684) );
  NAND2_X1 U773 ( .A1(G119), .A2(n880), .ZN(n683) );
  NAND2_X1 U774 ( .A1(n684), .A2(n683), .ZN(n685) );
  OR2_X1 U775 ( .A1(n686), .A2(n685), .ZN(n870) );
  NAND2_X1 U776 ( .A1(G1991), .A2(n870), .ZN(n687) );
  XNOR2_X1 U777 ( .A(n687), .B(KEYINPUT92), .ZN(n696) );
  NAND2_X1 U778 ( .A1(G141), .A2(n883), .ZN(n689) );
  NAND2_X1 U779 ( .A1(G129), .A2(n880), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n689), .A2(n688), .ZN(n692) );
  NAND2_X1 U781 ( .A1(n885), .A2(G105), .ZN(n690) );
  XOR2_X1 U782 ( .A(KEYINPUT38), .B(n690), .Z(n691) );
  NOR2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n694) );
  NAND2_X1 U784 ( .A1(n879), .A2(G117), .ZN(n693) );
  NAND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n874) );
  NAND2_X1 U786 ( .A1(G1996), .A2(n874), .ZN(n695) );
  NAND2_X1 U787 ( .A1(n696), .A2(n695), .ZN(n1009) );
  AND2_X1 U788 ( .A1(n818), .A2(n1009), .ZN(n809) );
  XOR2_X1 U789 ( .A(n809), .B(KEYINPUT93), .Z(n793) );
  INV_X1 U790 ( .A(n697), .ZN(n699) );
  XNOR2_X1 U791 ( .A(n745), .B(KEYINPUT95), .ZN(n718) );
  XNOR2_X1 U792 ( .A(G2078), .B(KEYINPUT25), .ZN(n971) );
  NAND2_X1 U793 ( .A1(n718), .A2(n971), .ZN(n701) );
  INV_X1 U794 ( .A(G1961), .ZN(n945) );
  NAND2_X1 U795 ( .A1(n745), .A2(n945), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n735) );
  NAND2_X1 U797 ( .A1(n735), .A2(G171), .ZN(n734) );
  NAND2_X1 U798 ( .A1(n718), .A2(G2072), .ZN(n703) );
  INV_X1 U799 ( .A(KEYINPUT27), .ZN(n702) );
  XNOR2_X1 U800 ( .A(n703), .B(n702), .ZN(n706) );
  INV_X1 U801 ( .A(n718), .ZN(n704) );
  NAND2_X1 U802 ( .A1(G1956), .A2(n704), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U804 ( .A1(n709), .A2(n924), .ZN(n708) );
  NOR2_X1 U805 ( .A1(n709), .A2(n924), .ZN(n710) );
  XNOR2_X1 U806 ( .A(KEYINPUT99), .B(n710), .ZN(n729) );
  INV_X1 U807 ( .A(G1341), .ZN(n946) );
  XOR2_X1 U808 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n715) );
  NAND2_X1 U809 ( .A1(n946), .A2(n715), .ZN(n711) );
  NAND2_X1 U810 ( .A1(n711), .A2(n745), .ZN(n714) );
  INV_X1 U811 ( .A(G1996), .ZN(n972) );
  NOR2_X1 U812 ( .A1(n972), .A2(n745), .ZN(n712) );
  NAND2_X1 U813 ( .A1(n712), .A2(n715), .ZN(n713) );
  NAND2_X1 U814 ( .A1(n714), .A2(n713), .ZN(n724) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n715), .ZN(n716) );
  NOR2_X1 U816 ( .A1(n716), .A2(n918), .ZN(n722) );
  NAND2_X1 U817 ( .A1(G1348), .A2(n745), .ZN(n717) );
  XNOR2_X1 U818 ( .A(n717), .B(KEYINPUT98), .ZN(n720) );
  NAND2_X1 U819 ( .A1(n718), .A2(G2067), .ZN(n719) );
  NAND2_X1 U820 ( .A1(n720), .A2(n719), .ZN(n725) );
  NAND2_X1 U821 ( .A1(n919), .A2(n725), .ZN(n721) );
  NAND2_X1 U822 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U823 ( .A1(n724), .A2(n723), .ZN(n727) );
  NOR2_X1 U824 ( .A1(n725), .A2(n919), .ZN(n726) );
  NOR2_X1 U825 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U826 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U827 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U828 ( .A(n732), .B(KEYINPUT29), .Z(n733) );
  NAND2_X1 U829 ( .A1(n734), .A2(n733), .ZN(n760) );
  INV_X1 U830 ( .A(KEYINPUT100), .ZN(n744) );
  NOR2_X1 U831 ( .A1(G171), .A2(n735), .ZN(n741) );
  NOR2_X1 U832 ( .A1(G1966), .A2(n788), .ZN(n762) );
  NOR2_X1 U833 ( .A1(G2084), .A2(n745), .ZN(n758) );
  INV_X1 U834 ( .A(n758), .ZN(n736) );
  NAND2_X1 U835 ( .A1(G8), .A2(n736), .ZN(n737) );
  OR2_X1 U836 ( .A1(n762), .A2(n737), .ZN(n738) );
  XNOR2_X1 U837 ( .A(KEYINPUT30), .B(n738), .ZN(n739) );
  NOR2_X1 U838 ( .A1(n739), .A2(G168), .ZN(n740) );
  XNOR2_X1 U839 ( .A(n742), .B(KEYINPUT31), .ZN(n743) );
  XNOR2_X1 U840 ( .A(n744), .B(n743), .ZN(n759) );
  INV_X1 U841 ( .A(G8), .ZN(n750) );
  NOR2_X1 U842 ( .A1(G1971), .A2(n788), .ZN(n747) );
  NOR2_X1 U843 ( .A1(G2090), .A2(n745), .ZN(n746) );
  NOR2_X1 U844 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U845 ( .A1(n748), .A2(G303), .ZN(n749) );
  OR2_X1 U846 ( .A1(n750), .A2(n749), .ZN(n752) );
  AND2_X1 U847 ( .A1(n759), .A2(n752), .ZN(n751) );
  NAND2_X1 U848 ( .A1(n760), .A2(n751), .ZN(n755) );
  INV_X1 U849 ( .A(n752), .ZN(n753) );
  OR2_X1 U850 ( .A1(n753), .A2(G286), .ZN(n754) );
  NAND2_X1 U851 ( .A1(n755), .A2(n754), .ZN(n757) );
  XOR2_X1 U852 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n756) );
  XNOR2_X1 U853 ( .A(n757), .B(n756), .ZN(n766) );
  NAND2_X1 U854 ( .A1(G8), .A2(n758), .ZN(n764) );
  AND2_X1 U855 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U856 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U857 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n787) );
  NOR2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n773) );
  NOR2_X1 U860 ( .A1(G1971), .A2(G303), .ZN(n767) );
  NOR2_X1 U861 ( .A1(n773), .A2(n767), .ZN(n925) );
  INV_X1 U862 ( .A(KEYINPUT33), .ZN(n768) );
  AND2_X1 U863 ( .A1(n925), .A2(n768), .ZN(n769) );
  NAND2_X1 U864 ( .A1(n787), .A2(n769), .ZN(n779) );
  XOR2_X1 U865 ( .A(G305), .B(G1981), .Z(n937) );
  INV_X1 U866 ( .A(n788), .ZN(n771) );
  NAND2_X1 U867 ( .A1(G288), .A2(G1976), .ZN(n770) );
  XNOR2_X1 U868 ( .A(n770), .B(KEYINPUT102), .ZN(n926) );
  AND2_X1 U869 ( .A1(n771), .A2(n926), .ZN(n772) );
  NOR2_X1 U870 ( .A1(KEYINPUT33), .A2(n772), .ZN(n776) );
  NAND2_X1 U871 ( .A1(n773), .A2(KEYINPUT33), .ZN(n774) );
  NOR2_X1 U872 ( .A1(n788), .A2(n774), .ZN(n775) );
  NOR2_X1 U873 ( .A1(n776), .A2(n775), .ZN(n777) );
  AND2_X1 U874 ( .A1(n937), .A2(n777), .ZN(n778) );
  NAND2_X1 U875 ( .A1(n779), .A2(n778), .ZN(n784) );
  NOR2_X1 U876 ( .A1(G305), .A2(G1981), .ZN(n780) );
  XOR2_X1 U877 ( .A(n780), .B(KEYINPUT24), .Z(n781) );
  XNOR2_X1 U878 ( .A(KEYINPUT94), .B(n781), .ZN(n782) );
  OR2_X1 U879 ( .A1(n788), .A2(n782), .ZN(n783) );
  NAND2_X1 U880 ( .A1(n784), .A2(n783), .ZN(n791) );
  NOR2_X1 U881 ( .A1(G2090), .A2(G303), .ZN(n785) );
  NAND2_X1 U882 ( .A1(G8), .A2(n785), .ZN(n786) );
  NAND2_X1 U883 ( .A1(n787), .A2(n786), .ZN(n789) );
  AND2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U885 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n805) );
  XNOR2_X1 U887 ( .A(KEYINPUT37), .B(G2067), .ZN(n815) );
  NAND2_X1 U888 ( .A1(G116), .A2(n879), .ZN(n795) );
  NAND2_X1 U889 ( .A1(G128), .A2(n880), .ZN(n794) );
  NAND2_X1 U890 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U891 ( .A(n796), .B(KEYINPUT35), .ZN(n801) );
  NAND2_X1 U892 ( .A1(G104), .A2(n885), .ZN(n798) );
  NAND2_X1 U893 ( .A1(G140), .A2(n883), .ZN(n797) );
  NAND2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U895 ( .A(KEYINPUT34), .B(n799), .Z(n800) );
  NAND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U897 ( .A(n802), .B(KEYINPUT36), .Z(n893) );
  NOR2_X1 U898 ( .A1(n815), .A2(n893), .ZN(n994) );
  NAND2_X1 U899 ( .A1(n818), .A2(n994), .ZN(n812) );
  INV_X1 U900 ( .A(n812), .ZN(n803) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n932) );
  XNOR2_X1 U902 ( .A(n806), .B(KEYINPUT103), .ZN(n820) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n874), .ZN(n1005) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n870), .ZN(n995) );
  NOR2_X1 U906 ( .A1(n807), .A2(n995), .ZN(n808) );
  NOR2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U908 ( .A1(n1005), .A2(n810), .ZN(n811) );
  XNOR2_X1 U909 ( .A(n811), .B(KEYINPUT39), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U911 ( .A(n814), .B(KEYINPUT104), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n815), .A2(n893), .ZN(n1018) );
  NAND2_X1 U913 ( .A1(n816), .A2(n1018), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U916 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n822), .ZN(G217) );
  NAND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n823) );
  XOR2_X1 U919 ( .A(KEYINPUT106), .B(n823), .Z(n824) );
  NAND2_X1 U920 ( .A1(n824), .A2(G661), .ZN(n825) );
  XOR2_X1 U921 ( .A(KEYINPUT107), .B(n825), .Z(G259) );
  NAND2_X1 U922 ( .A1(G1), .A2(G3), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U924 ( .A(n828), .B(KEYINPUT108), .ZN(G188) );
  NOR2_X1 U925 ( .A1(n830), .A2(n829), .ZN(G325) );
  XNOR2_X1 U926 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U929 ( .A(n918), .B(n831), .ZN(n832) );
  NOR2_X1 U930 ( .A1(n832), .A2(G860), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(G145) );
  INV_X1 U932 ( .A(n835), .ZN(G319) );
  XOR2_X1 U933 ( .A(G2096), .B(G2678), .Z(n837) );
  XNOR2_X1 U934 ( .A(G2090), .B(KEYINPUT43), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U936 ( .A(n838), .B(KEYINPUT42), .Z(n840) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2072), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U939 ( .A(KEYINPUT110), .B(G2100), .Z(n842) );
  XNOR2_X1 U940 ( .A(G2084), .B(G2078), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1981), .B(G1961), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1991), .B(G1966), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n848) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1956), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U949 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U950 ( .A(G2474), .B(KEYINPUT111), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U952 ( .A(KEYINPUT41), .B(n853), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n854), .B(n972), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G100), .A2(n885), .ZN(n856) );
  NAND2_X1 U955 ( .A1(G112), .A2(n879), .ZN(n855) );
  NAND2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G124), .A2(n880), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n857), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U959 ( .A1(n883), .A2(G136), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U961 ( .A1(n861), .A2(n860), .ZN(G162) );
  XNOR2_X1 U962 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n872) );
  NAND2_X1 U963 ( .A1(G103), .A2(n885), .ZN(n863) );
  NAND2_X1 U964 ( .A1(G139), .A2(n883), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G115), .A2(n879), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G127), .A2(n880), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U969 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U971 ( .A(KEYINPUT113), .B(n869), .Z(n1012) );
  XNOR2_X1 U972 ( .A(n870), .B(n1012), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U974 ( .A(n996), .B(G162), .Z(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(n876), .B(n875), .Z(n878) );
  XNOR2_X1 U977 ( .A(G164), .B(G160), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n892) );
  NAND2_X1 U979 ( .A1(G118), .A2(n879), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G130), .A2(n880), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n890) );
  NAND2_X1 U982 ( .A1(n883), .A2(G142), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n884), .B(KEYINPUT112), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G106), .A2(n885), .ZN(n886) );
  NAND2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U986 ( .A(n888), .B(KEYINPUT45), .Z(n889) );
  NOR2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U988 ( .A(n892), .B(n891), .Z(n894) );
  XOR2_X1 U989 ( .A(n894), .B(n893), .Z(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U991 ( .A(n896), .B(KEYINPUT114), .ZN(n898) );
  XNOR2_X1 U992 ( .A(n919), .B(G286), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U994 ( .A(G171), .B(n899), .Z(n900) );
  NOR2_X1 U995 ( .A1(G37), .A2(n900), .ZN(n901) );
  XOR2_X1 U996 ( .A(KEYINPUT115), .B(n901), .Z(G397) );
  XOR2_X1 U997 ( .A(G2454), .B(G2435), .Z(n903) );
  XNOR2_X1 U998 ( .A(G2438), .B(G2427), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n910) );
  XOR2_X1 U1000 ( .A(KEYINPUT105), .B(G2446), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G2443), .B(G2430), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1003 ( .A(n906), .B(G2451), .Z(n908) );
  XNOR2_X1 U1004 ( .A(G1348), .B(G1341), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(n911), .A2(G14), .ZN(n917) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n917), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G57), .ZN(G237) );
  INV_X1 U1016 ( .A(n917), .ZN(G401) );
  XNOR2_X1 U1017 ( .A(KEYINPUT56), .B(G16), .ZN(n943) );
  XNOR2_X1 U1018 ( .A(n946), .B(n918), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(G301), .B(G1961), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n919), .B(G1348), .ZN(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n936) );
  XOR2_X1 U1023 ( .A(n924), .B(G1956), .Z(n931) );
  AND2_X1 U1024 ( .A1(G303), .A2(G1971), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(KEYINPUT124), .B(n929), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(KEYINPUT125), .B(n934), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n941) );
  XNOR2_X1 U1032 ( .A(G1966), .B(G168), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(n939), .B(KEYINPUT57), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(KEYINPUT126), .B(n944), .ZN(n1027) );
  XNOR2_X1 U1038 ( .A(G5), .B(n945), .ZN(n959) );
  XNOR2_X1 U1039 ( .A(G19), .B(n946), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(G1956), .B(G20), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(G1981), .B(G6), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n953) );
  XOR2_X1 U1044 ( .A(KEYINPUT59), .B(G1348), .Z(n951) );
  XNOR2_X1 U1045 ( .A(G4), .B(n951), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n955) );
  XOR2_X1 U1047 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n954) );
  XOR2_X1 U1048 ( .A(n955), .B(n954), .Z(n957) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G21), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n966) );
  XNOR2_X1 U1052 ( .A(G1971), .B(G22), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(G23), .B(G1976), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n963) );
  XOR2_X1 U1055 ( .A(G1986), .B(G24), .Z(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(KEYINPUT58), .B(n964), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT61), .B(n967), .ZN(n969) );
  INV_X1 U1060 ( .A(G16), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n970), .A2(G11), .ZN(n1025) );
  XNOR2_X1 U1063 ( .A(G2090), .B(G35), .ZN(n987) );
  XNOR2_X1 U1064 ( .A(n971), .B(G27), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n972), .B(G32), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(KEYINPUT121), .B(n975), .ZN(n977) );
  XOR2_X1 U1068 ( .A(G2072), .B(G33), .Z(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G26), .B(G2067), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(KEYINPUT122), .B(n980), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n981), .A2(G28), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(G25), .B(G1991), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(KEYINPUT120), .B(n982), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT53), .B(n985), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n990) );
  XOR2_X1 U1079 ( .A(G2084), .B(G34), .Z(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT54), .B(n988), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(KEYINPUT123), .B(n991), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(G29), .A2(n992), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n993), .B(KEYINPUT55), .ZN(n1023) );
  INV_X1 U1085 ( .A(n994), .ZN(n999) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(KEYINPUT116), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(G2084), .B(G160), .Z(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1091 ( .A(KEYINPUT117), .B(n1002), .Z(n1011) );
  XOR2_X1 U1092 ( .A(G2090), .B(G162), .Z(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT118), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n1006) );
  XNOR2_X1 U1096 ( .A(n1007), .B(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1017) );
  XOR2_X1 U1099 ( .A(G2072), .B(n1012), .Z(n1014) );
  XOR2_X1 U1100 ( .A(G164), .B(G2078), .Z(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT50), .B(n1015), .Z(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT52), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(G29), .A2(n1021), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1109 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

