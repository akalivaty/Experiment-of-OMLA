//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G125), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n459), .A2(G137), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g046(.A(new_n471), .B(KEYINPUT69), .Z(G160));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n459), .B(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(new_n465), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n465), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n476), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT71), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT72), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n465), .A2(G114), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT72), .A4(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n459), .A2(G126), .A3(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n494), .B(new_n495), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n459), .B2(new_n494), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n491), .B(new_n492), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n497), .A2(new_n496), .ZN(new_n504));
  NAND2_X1  g079(.A1(G126), .A2(G2105), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n494), .B1(new_n497), .B2(new_n496), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n506), .B1(new_n508), .B2(new_n498), .ZN(new_n509));
  AOI21_X1  g084(.A(KEYINPUT73), .B1(new_n509), .B2(new_n491), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n503), .A2(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n514), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n512), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G166));
  NAND2_X1  g103(.A1(new_n515), .A2(G51), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT74), .B(G89), .Z(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G168));
  NAND2_X1  g111(.A1(new_n515), .A2(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n522), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n526), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n542));
  OR3_X1    g117(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n539), .B2(new_n541), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(new_n515), .A2(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n522), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n526), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n515), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n519), .A2(new_n520), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n517), .A2(new_n521), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n562), .A2(G651), .B1(new_n563), .B2(G91), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n558), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  INV_X1    g141(.A(G168), .ZN(G286));
  XNOR2_X1  g142(.A(G166), .B(KEYINPUT76), .ZN(G303));
  NAND2_X1  g143(.A1(new_n515), .A2(G49), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n522), .ZN(G288));
  AOI22_X1  g147(.A1(new_n563), .A2(G86), .B1(G48), .B2(new_n515), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n519), .B2(new_n520), .ZN(new_n575));
  AND2_X1   g150(.A1(G73), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G305));
  NAND2_X1  g153(.A1(new_n515), .A2(G47), .ZN(new_n579));
  INV_X1    g154(.A(G85), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n522), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n526), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n560), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n526), .B1(new_n588), .B2(KEYINPUT77), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(KEYINPUT77), .B2(new_n588), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n515), .A2(G54), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n517), .A2(new_n521), .A3(G92), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT10), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g171(.A(new_n595), .B1(G171), .B2(G868), .ZN(G321));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G299), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G297));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G280));
  AND3_X1   g176(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n602));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(KEYINPUT78), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(KEYINPUT78), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n607), .B(new_n608), .C1(G868), .C2(new_n551), .ZN(G323));
  XNOR2_X1  g184(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n610));
  XNOR2_X1  g185(.A(G323), .B(new_n610), .ZN(G282));
  NAND2_X1  g186(.A1(new_n475), .A2(G135), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT80), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n465), .A2(G111), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n615));
  OAI221_X1 g190(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n615), .B2(new_n614), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n477), .B2(G123), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2096), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(G2096), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n459), .A2(new_n468), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(G156));
  XOR2_X1   g201(.A(G2451), .B(G2454), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n633), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n630), .B(new_n636), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(G14), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n638), .ZN(G401));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT17), .Z(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  INV_X1    g223(.A(new_n645), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(new_n643), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n647), .B(new_n648), .C1(new_n646), .C2(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n648), .A2(new_n643), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT18), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(G2100), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT82), .B(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT20), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n664), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n666), .B(new_n668), .C1(new_n661), .C2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G229));
  NOR2_X1   g251(.A1(G29), .A2(G35), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(G162), .B2(G29), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT29), .Z(new_n679));
  INV_X1    g254(.A(G2090), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT98), .Z(new_n682));
  OR2_X1    g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  INV_X1    g258(.A(G34), .ZN(new_n684));
  AOI21_X1  g259(.A(G29), .B1(new_n684), .B2(KEYINPUT24), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(KEYINPUT24), .B2(new_n684), .ZN(new_n686));
  INV_X1    g261(.A(G160), .ZN(new_n687));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G2084), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT93), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(G27), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G164), .B2(new_n688), .ZN(new_n694));
  INV_X1    g269(.A(G2078), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n475), .A2(G141), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n477), .A2(G129), .ZN(new_n699));
  NAND3_X1  g274(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT26), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n702), .A2(new_n703), .B1(G105), .B2(new_n468), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n698), .A2(new_n699), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(new_n688), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n688), .B2(G32), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT27), .B(G1996), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT94), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n708), .A2(new_n710), .B1(new_n689), .B2(new_n690), .ZN(new_n711));
  NOR2_X1   g286(.A1(G5), .A2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT96), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(G301), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT97), .B(G1961), .ZN(new_n717));
  OAI221_X1 g292(.A(new_n711), .B1(new_n716), .B2(new_n717), .C1(new_n710), .C2(new_n708), .ZN(new_n718));
  INV_X1    g293(.A(G21), .ZN(new_n719));
  AOI21_X1  g294(.A(KEYINPUT95), .B1(new_n714), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(G168), .A2(G16), .ZN(new_n721));
  MUX2_X1   g296(.A(KEYINPUT95), .B(new_n720), .S(new_n721), .Z(new_n722));
  OAI22_X1  g297(.A1(G1966), .A2(new_n722), .B1(new_n619), .B2(new_n688), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G1966), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n551), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G16), .B2(G19), .ZN(new_n726));
  INV_X1    g301(.A(G1341), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT30), .B(G28), .ZN(new_n729));
  OR2_X1    g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  NAND2_X1  g305(.A1(KEYINPUT31), .A2(G11), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n729), .A2(new_n688), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n726), .B2(new_n727), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n728), .B(new_n733), .C1(new_n716), .C2(new_n717), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT25), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n475), .B2(G139), .ZN(new_n737));
  NAND2_X1  g312(.A1(G115), .A2(G2104), .ZN(new_n738));
  INV_X1    g313(.A(G127), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n504), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n465), .B1(new_n740), .B2(KEYINPUT92), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(KEYINPUT92), .B2(new_n740), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  MUX2_X1   g318(.A(G33), .B(new_n743), .S(G29), .Z(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(G2072), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n688), .A2(G26), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT28), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n475), .A2(G140), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n477), .A2(G128), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n465), .A2(G116), .ZN(new_n750));
  OAI21_X1  g325(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n748), .B(new_n749), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n747), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2067), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n724), .A2(new_n734), .A3(new_n745), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n602), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G4), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1348), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n714), .A2(G20), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT23), .Z(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G299), .B2(G16), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1956), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n759), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n697), .A2(new_n718), .A3(new_n755), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n682), .A2(new_n683), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G166), .A2(new_n714), .ZN(new_n768));
  INV_X1    g343(.A(G1971), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n714), .A2(G22), .ZN(new_n770));
  OR3_X1    g345(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G6), .A2(G16), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n563), .A2(G86), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n515), .A2(G48), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n775), .A2(new_n577), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n774), .B1(new_n777), .B2(G16), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT32), .B(G1981), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G23), .B(G288), .S(G16), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT33), .B(G1976), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n773), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT34), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G1986), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G24), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(G290), .A2(KEYINPUT87), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT87), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n584), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n787), .B(new_n789), .C1(new_n793), .C2(new_n714), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n714), .B1(new_n790), .B2(new_n792), .ZN(new_n795));
  OAI21_X1  g370(.A(G1986), .B1(new_n795), .B2(new_n788), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n773), .A2(new_n780), .A3(new_n785), .A4(new_n783), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n688), .A2(G25), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(new_n465), .B2(G107), .ZN(new_n801));
  OR3_X1    g376(.A1(KEYINPUT86), .A2(G95), .A3(G2105), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT86), .B1(G95), .B2(G2105), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n475), .B2(G131), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n477), .A2(KEYINPUT85), .A3(G119), .ZN(new_n806));
  AOI21_X1  g381(.A(KEYINPUT85), .B1(new_n477), .B2(G119), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n800), .B1(new_n808), .B2(G29), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(KEYINPUT88), .B1(new_n799), .B2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n810), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n809), .B(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT88), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n814), .A2(new_n815), .A3(new_n798), .A4(new_n797), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n786), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT36), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT90), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n817), .A2(new_n818), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n821), .B1(new_n817), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n822), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n819), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT91), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT91), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n823), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n767), .B1(new_n829), .B2(new_n831), .ZN(G311));
  INV_X1    g407(.A(new_n767), .ZN(new_n833));
  INV_X1    g408(.A(new_n831), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n830), .B1(new_n823), .B2(new_n827), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(G150));
  NAND2_X1  g411(.A1(new_n602), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n515), .A2(G55), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n522), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n526), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n551), .B(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n838), .B(new_n845), .Z(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  INV_X1    g422(.A(G860), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n844), .A2(new_n848), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT99), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT37), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(G145));
  XNOR2_X1  g429(.A(new_n752), .B(new_n501), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(new_n706), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n706), .ZN(new_n857));
  OR3_X1    g432(.A1(new_n856), .A2(new_n857), .A3(new_n743), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n743), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n808), .B(new_n623), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n477), .A2(G130), .ZN(new_n862));
  OR2_X1    g437(.A1(G106), .A2(G2105), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n863), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(G142), .B2(new_n475), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n861), .B(new_n866), .Z(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n860), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n858), .A3(new_n859), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(G162), .A2(new_n619), .ZN(new_n872));
  NAND2_X1  g447(.A1(G162), .A2(new_n619), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT100), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n687), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(G160), .A3(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(G37), .B1(new_n871), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n870), .A2(KEYINPUT101), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n860), .B1(new_n868), .B2(KEYINPUT101), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n880), .A3(new_n879), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n602), .A2(new_n599), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n594), .A2(G299), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT41), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n893), .A3(new_n890), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n888), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT103), .B1(new_n891), .B2(KEYINPUT41), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n845), .B(KEYINPUT102), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n605), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n891), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n901), .B2(new_n899), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n584), .B(G305), .ZN(new_n903));
  XNOR2_X1  g478(.A(G166), .B(G288), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(KEYINPUT104), .B2(KEYINPUT42), .ZN(new_n906));
  NAND2_X1  g481(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT105), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n906), .B(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n902), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G868), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(G868), .B2(new_n844), .ZN(G295));
  OAI21_X1  g487(.A(new_n911), .B1(G868), .B2(new_n844), .ZN(G331));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(new_n543), .B2(new_n544), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n845), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n845), .A2(new_n916), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n543), .A2(new_n915), .A3(new_n544), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n918), .A2(new_n919), .B1(G286), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n919), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(G286), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n922), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  OAI22_X1  g499(.A1(new_n895), .A2(new_n896), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n923), .B1(new_n922), .B2(new_n917), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n901), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n905), .B1(new_n929), .B2(KEYINPUT107), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n925), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n905), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT108), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n925), .A2(new_n928), .A3(new_n936), .A4(new_n905), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n914), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n921), .A2(new_n924), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n892), .A2(new_n894), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n928), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n942), .B2(new_n934), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n938), .A2(new_n914), .A3(new_n943), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n939), .A2(new_n944), .A3(KEYINPUT44), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n938), .A2(new_n943), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n933), .A2(new_n914), .A3(new_n938), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n945), .A2(new_n950), .ZN(G397));
  AOI21_X1  g526(.A(new_n465), .B1(new_n460), .B2(new_n462), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n466), .A2(new_n469), .ZN(new_n953));
  INV_X1    g528(.A(G40), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(G1384), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n957), .B1(new_n509), .B2(new_n491), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n958), .B2(KEYINPUT45), .ZN(new_n959));
  INV_X1    g534(.A(new_n957), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n501), .A2(new_n956), .A3(KEYINPUT45), .A4(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n955), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n501), .A2(new_n502), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n509), .A2(KEYINPUT73), .A3(new_n491), .ZN(new_n965));
  AOI21_X1  g540(.A(G1384), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(KEYINPUT45), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n963), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n503), .B2(new_n510), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n464), .A2(new_n470), .A3(G40), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n960), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT111), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n976), .B2(new_n961), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT112), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n695), .B1(new_n969), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n980));
  INV_X1    g555(.A(G1961), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n509), .B2(new_n491), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n974), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n966), .B2(new_n983), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT118), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n984), .B(new_n987), .C1(new_n966), .C2(new_n983), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n979), .A2(new_n980), .B1(new_n981), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n955), .B1(new_n982), .B2(KEYINPUT45), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(KEYINPUT45), .B2(new_n966), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(KEYINPUT53), .A3(new_n695), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G171), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT125), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n470), .B(KEYINPUT124), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n980), .A2(new_n954), .A3(G2078), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n464), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n958), .A2(KEYINPUT45), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n959), .B2(new_n962), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n990), .A2(new_n996), .A3(G301), .A4(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n986), .A2(new_n981), .A3(new_n988), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n968), .B1(new_n963), .B2(new_n967), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n973), .A2(new_n977), .A3(KEYINPUT112), .ZN(new_n1006));
  AOI21_X1  g581(.A(G2078), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1004), .B(new_n1002), .C1(new_n1007), .C2(KEYINPUT53), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT125), .B1(new_n1008), .B2(G171), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n995), .A2(new_n1003), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(G171), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n979), .A2(new_n980), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1014), .A2(G301), .A3(new_n1004), .A4(new_n993), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n1015), .A3(KEYINPUT54), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1005), .A2(new_n769), .A3(new_n1006), .ZN(new_n1017));
  AOI211_X1 g592(.A(KEYINPUT50), .B(G1384), .C1(new_n964), .C2(new_n965), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n955), .B1(new_n982), .B2(new_n983), .ZN(new_n1019));
  OR3_X1    g594(.A1(new_n1018), .A2(G2090), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT117), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1017), .A2(new_n1023), .A3(new_n1020), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(G8), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G303), .A2(G8), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT55), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n966), .A2(KEYINPUT45), .ZN(new_n1033));
  INV_X1    g608(.A(new_n991), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1966), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n984), .B(new_n690), .C1(new_n966), .C2(new_n983), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(G286), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1038), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1966), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1041));
  OAI21_X1  g616(.A(G168), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1032), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(G168), .B(new_n1038), .C1(new_n992), .C2(G1966), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT51), .B1(new_n1044), .B2(G8), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1030), .B1(new_n982), .B2(new_n955), .ZN(new_n1047));
  INV_X1    g622(.A(G1981), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n775), .A2(new_n1048), .A3(new_n577), .A4(new_n776), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n573), .A2(KEYINPUT113), .A3(new_n1048), .A4(new_n577), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1051), .A2(new_n1052), .B1(G1981), .B2(G305), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1047), .B1(new_n1053), .B2(KEYINPUT49), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G305), .A2(G1981), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1055), .A2(KEYINPUT49), .A3(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1976), .ZN(new_n1059));
  OR2_X1    g634(.A1(G288), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1047), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1047), .A2(new_n1060), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1058), .A2(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n985), .A2(G2090), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1030), .B1(new_n1017), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1027), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AND4_X1   g646(.A1(new_n1016), .A2(new_n1028), .A3(new_n1046), .A4(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n986), .A2(new_n758), .A3(new_n988), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  INV_X1    g649(.A(G2067), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n982), .A2(new_n1075), .A3(new_n955), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1074), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT60), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT119), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT60), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1079), .A2(new_n1084), .A3(new_n602), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT60), .B(new_n594), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n973), .A2(new_n977), .A3(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(G299), .B(KEYINPUT57), .Z(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1088), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1089), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT123), .B1(new_n1094), .B2(KEYINPUT61), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  NOR4_X1   g672(.A1(new_n1092), .A2(new_n1093), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1086), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1097), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT122), .ZN(new_n1101));
  INV_X1    g676(.A(G1996), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n973), .A2(new_n977), .A3(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT58), .B(G1341), .Z(new_n1104));
  INV_X1    g679(.A(new_n982), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n974), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n551), .A2(KEYINPUT120), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT121), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1107), .A2(new_n1112), .A3(new_n1109), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1111), .A2(KEYINPUT59), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1116));
  AOI211_X1 g691(.A(KEYINPUT121), .B(new_n1108), .C1(new_n1103), .C2(new_n1106), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1119), .B(new_n1097), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1101), .A2(new_n1114), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1085), .A2(new_n1099), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1081), .A2(new_n602), .A3(new_n1083), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1093), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1092), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1012), .B(new_n1072), .C1(new_n1122), .C2(new_n1125), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1042), .A2(new_n1030), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT114), .B1(new_n1058), .B2(new_n1066), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT114), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1130), .A2(new_n1065), .A3(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(KEYINPUT63), .B(new_n1128), .C1(new_n1129), .C2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1127), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1017), .A2(new_n1023), .A3(new_n1020), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1023), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1030), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1071), .B(new_n1128), .C1(new_n1138), .C2(new_n1070), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1135), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1047), .B(KEYINPUT115), .Z(new_n1142));
  OR3_X1    g717(.A1(new_n1130), .A2(G1976), .A3(G288), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1055), .B(KEYINPUT116), .Z(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1127), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1071), .B1(new_n1138), .B2(new_n1070), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1040), .A2(new_n1041), .A3(G168), .ZN(new_n1149));
  AOI21_X1  g724(.A(G286), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1031), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1045), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n1152), .A3(KEYINPUT62), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n994), .A2(new_n1153), .A3(new_n1155), .A4(G171), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1147), .B1(new_n1148), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1141), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1126), .A2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n958), .A2(new_n974), .A3(KEYINPUT45), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1102), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT110), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1162), .A2(new_n706), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1160), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n752), .B(new_n1075), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n705), .A2(G1996), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n808), .B(new_n810), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1168), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n584), .B(new_n787), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1160), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1159), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT46), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1162), .B(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1165), .A2(new_n706), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1160), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT47), .ZN(new_n1179));
  NOR4_X1   g754(.A1(new_n1163), .A2(new_n1167), .A3(new_n813), .A4(new_n808), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n752), .A2(G2067), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1160), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1160), .A2(new_n787), .A3(new_n584), .ZN(new_n1183));
  XOR2_X1   g758(.A(new_n1183), .B(KEYINPUT48), .Z(new_n1184));
  OAI211_X1 g759(.A(new_n1179), .B(new_n1182), .C1(new_n1170), .C2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1173), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g763(.A(G319), .ZN(new_n1190));
  NOR4_X1   g764(.A1(G229), .A2(new_n1190), .A3(G401), .A4(G227), .ZN(new_n1191));
  OAI211_X1 g765(.A(new_n886), .B(new_n1191), .C1(new_n939), .C2(new_n944), .ZN(G225));
  INV_X1    g766(.A(G225), .ZN(G308));
endmodule


