//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n554, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1134, new_n1135;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n453), .A2(G567), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n457), .B1(new_n452), .B2(G2106), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n462), .A3(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(KEYINPUT3), .A3(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n463), .A2(new_n468), .A3(G137), .A4(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(new_n467), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G101), .A3(new_n469), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n471), .B1(new_n470), .B2(new_n473), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT67), .Z(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G125), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NOR3_X1   g055(.A1(new_n474), .A2(new_n475), .A3(new_n480), .ZN(G160));
  NAND3_X1  g056(.A1(new_n463), .A2(new_n468), .A3(new_n469), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n463), .A2(new_n468), .A3(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n463), .A2(new_n468), .A3(G138), .A4(new_n469), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n478), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n463), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  XNOR2_X1  g077(.A(KEYINPUT71), .B(G651), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n511), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT72), .A3(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n512), .A2(new_n514), .B1(KEYINPUT5), .B2(new_n507), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n509), .B1(new_n510), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(new_n503), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n519), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n517), .A2(G89), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT73), .B(G51), .Z(new_n526));
  NAND2_X1  g101(.A1(new_n508), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n515), .A2(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n525), .A2(new_n527), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(new_n508), .A2(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n536), .B2(new_n518), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n521), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n516), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(new_n503), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n544), .B(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(G43), .A2(new_n508), .B1(new_n517), .B2(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G860), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT75), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT76), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n508), .A2(G53), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(KEYINPUT77), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n558), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n516), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n517), .A2(G91), .B1(G651), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  NAND2_X1  g142(.A1(new_n517), .A2(G87), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT78), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT79), .Z(new_n571));
  NAND2_X1  g146(.A1(new_n508), .A2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(G288));
  OAI211_X1 g148(.A(G86), .B(new_n515), .C1(new_n504), .C2(new_n505), .ZN(new_n574));
  OAI211_X1 g149(.A(G48), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n515), .A2(G61), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT80), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n521), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n576), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n521), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n518), .A2(new_n584), .ZN(new_n585));
  AOI211_X1 g160(.A(new_n583), .B(new_n585), .C1(G47), .C2(new_n508), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT81), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n517), .A2(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n516), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n508), .A2(G54), .B1(G651), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n588), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n588), .B1(new_n597), .B2(G868), .ZN(G321));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G299), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n600), .B2(G168), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(new_n600), .B2(G168), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  NOR2_X1   g180(.A1(new_n596), .A2(G559), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n606), .A2(KEYINPUT82), .A3(new_n600), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT82), .B1(new_n606), .B2(new_n600), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n546), .A2(new_n547), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n607), .B(new_n608), .C1(G868), .C2(new_n609), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n472), .A2(new_n469), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n613), .A2(new_n478), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT12), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2100), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n483), .A2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n486), .A2(G123), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n469), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT83), .B(G2096), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n624), .ZN(G156));
  XOR2_X1   g200(.A(G1341), .B(G1348), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT85), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n629), .B(new_n635), .Z(new_n636));
  XOR2_X1   g211(.A(G2451), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  AOI21_X1  g223(.A(KEYINPUT18), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n646), .B2(KEYINPUT18), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n649), .B(new_n651), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT86), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1961), .B(G1966), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT87), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT20), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n657), .A2(new_n659), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n662), .A3(new_n660), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n664), .B(new_n667), .C1(new_n662), .C2(new_n666), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G229));
  NOR2_X1   g249(.A1(G4), .A2(G16), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n597), .B2(G16), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1348), .ZN(new_n677));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G20), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT23), .Z(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G299), .B2(G16), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(G1956), .Z(new_n682));
  INV_X1    g257(.A(G29), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G26), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n483), .A2(G140), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n486), .A2(G128), .ZN(new_n687));
  OR2_X1    g262(.A1(G104), .A2(G2105), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n688), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n685), .B1(new_n691), .B2(new_n683), .ZN(new_n692));
  INV_X1    g267(.A(G2067), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n683), .A2(G35), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G162), .B2(new_n683), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT29), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n694), .B1(new_n698), .B2(G2090), .ZN(new_n699));
  NOR3_X1   g274(.A1(new_n677), .A2(new_n682), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n609), .A2(new_n678), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n678), .B2(G19), .ZN(new_n702));
  INV_X1    g277(.A(G1341), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n702), .A2(new_n703), .B1(new_n698), .B2(G2090), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n700), .B(new_n704), .C1(new_n703), .C2(new_n702), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n678), .A2(G21), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G168), .B2(new_n678), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT95), .ZN(new_n708));
  INV_X1    g283(.A(G1966), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT30), .B(G28), .ZN(new_n712));
  OR2_X1    g287(.A1(KEYINPUT31), .A2(G11), .ZN(new_n713));
  NAND2_X1  g288(.A1(KEYINPUT31), .A2(G11), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n712), .A2(new_n683), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(new_n622), .B2(new_n683), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT96), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n678), .A2(G5), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G171), .B2(new_n678), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n717), .B1(new_n719), .B2(G1961), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n710), .A2(new_n711), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT97), .Z(new_n722));
  INV_X1    g297(.A(KEYINPUT24), .ZN(new_n723));
  INV_X1    g298(.A(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n723), .B2(new_n724), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G160), .B2(new_n683), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT91), .Z(new_n728));
  INV_X1    g303(.A(G2084), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n683), .A2(G33), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT25), .Z(new_n733));
  AOI22_X1  g308(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  INV_X1    g309(.A(G139), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n733), .B1(new_n734), .B2(new_n469), .C1(new_n735), .C2(new_n482), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(G29), .ZN(new_n737));
  INV_X1    g312(.A(G2072), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT93), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n683), .A2(G32), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n483), .A2(G141), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n486), .A2(G129), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT26), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n613), .A2(G105), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n743), .A2(new_n744), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n742), .B1(new_n750), .B2(G29), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n739), .B1(new_n741), .B2(new_n751), .C1(new_n719), .C2(G1961), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n741), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT94), .Z(new_n754));
  NOR2_X1   g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n728), .A2(new_n729), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n737), .A2(new_n738), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT92), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n683), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n683), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(G2078), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n760), .A2(G2078), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n758), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n755), .A2(new_n756), .A3(new_n763), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n722), .A2(new_n730), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n705), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n678), .A2(G22), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G166), .B2(new_n678), .ZN(new_n769));
  INV_X1    g344(.A(G1971), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n678), .A2(G23), .ZN(new_n772));
  INV_X1    g347(.A(G288), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n678), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT33), .B(G1976), .Z(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NOR2_X1   g352(.A1(G6), .A2(G16), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n576), .A2(new_n580), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(G16), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT32), .B(G1981), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n771), .A2(new_n776), .A3(new_n777), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(KEYINPUT34), .ZN(new_n784));
  NAND2_X1  g359(.A1(G290), .A2(G16), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n678), .A2(G24), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT88), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(KEYINPUT88), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n789), .A2(G1986), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(G1986), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n683), .A2(G25), .ZN(new_n792));
  OR2_X1    g367(.A1(G95), .A2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n794));
  INV_X1    g369(.A(G131), .ZN(new_n795));
  INV_X1    g370(.A(G119), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n794), .B1(new_n482), .B2(new_n795), .C1(new_n796), .C2(new_n485), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n792), .B1(new_n798), .B2(new_n683), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT35), .B(G1991), .Z(new_n800));
  XOR2_X1   g375(.A(new_n799), .B(new_n800), .Z(new_n801));
  NOR4_X1   g376(.A1(new_n784), .A2(new_n790), .A3(new_n791), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n783), .A2(KEYINPUT34), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT89), .B(KEYINPUT36), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n767), .B1(new_n766), .B2(new_n765), .C1(new_n805), .C2(KEYINPUT90), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(KEYINPUT90), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n802), .A2(new_n803), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(KEYINPUT36), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n809), .ZN(G311));
  INV_X1    g385(.A(G311), .ZN(G150));
  NOR2_X1   g386(.A1(new_n609), .A2(KEYINPUT100), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n521), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT99), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n508), .A2(G55), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n518), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n548), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n812), .B(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT38), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n597), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n826), .A2(new_n549), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n819), .A2(new_n549), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT37), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(G145));
  NAND2_X1  g406(.A1(new_n486), .A2(G130), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n469), .A2(G118), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G142), .B2(new_n483), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(new_n615), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n750), .B(new_n736), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT101), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n498), .A2(new_n840), .A3(new_n500), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n840), .B1(new_n498), .B2(new_n500), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n497), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n690), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n798), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n839), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(G160), .B(new_n622), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n490), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT102), .Z(new_n850));
  AOI21_X1  g425(.A(G37), .B1(new_n846), .B2(new_n848), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(G395));
  XNOR2_X1  g429(.A(G290), .B(G303), .ZN(new_n855));
  XNOR2_X1  g430(.A(G288), .B(G305), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(G299), .B(new_n596), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT41), .ZN(new_n861));
  INV_X1    g436(.A(new_n860), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n822), .B(new_n606), .Z(new_n863));
  MUX2_X1   g438(.A(new_n861), .B(new_n862), .S(new_n863), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n859), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G868), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(G868), .B2(new_n819), .ZN(G295));
  OAI21_X1  g442(.A(new_n866), .B1(G868), .B2(new_n819), .ZN(G331));
  XNOR2_X1  g443(.A(G171), .B(G286), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n822), .B(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(new_n861), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n860), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(G37), .B1(new_n876), .B2(new_n857), .ZN(new_n877));
  INV_X1    g452(.A(new_n857), .ZN(new_n878));
  INV_X1    g453(.A(new_n873), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n871), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n878), .B1(new_n874), .B2(new_n875), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT43), .B1(new_n877), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT44), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n881), .A2(KEYINPUT43), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n882), .B1(new_n877), .B2(new_n884), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n886), .B1(new_n889), .B2(KEYINPUT44), .ZN(G397));
  AOI21_X1  g465(.A(KEYINPUT106), .B1(G160), .B2(G40), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n470), .A2(new_n473), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT70), .ZN(new_n893));
  INV_X1    g468(.A(new_n480), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n893), .A2(new_n894), .A3(G40), .A4(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT45), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n492), .A2(KEYINPUT4), .B1(new_n478), .B2(new_n495), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n498), .A2(new_n500), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT101), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n498), .A2(new_n840), .A3(new_n500), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n900), .B1(new_n905), .B2(G1384), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n899), .A2(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n907), .A2(KEYINPUT107), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(KEYINPUT107), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n690), .B(new_n693), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n911), .B1(new_n750), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G1996), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(KEYINPUT46), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n910), .B2(G1996), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n919), .B(KEYINPUT47), .Z(new_n920));
  OR3_X1    g495(.A1(new_n910), .A2(G1986), .A3(G290), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n750), .B(new_n915), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n798), .A2(new_n800), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n798), .A2(new_n800), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n925), .A2(new_n912), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  AOI211_X1 g503(.A(new_n923), .B(new_n924), .C1(new_n911), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n925), .A2(new_n912), .ZN(new_n930));
  OAI22_X1  g505(.A1(new_n930), .A2(new_n927), .B1(G2067), .B2(new_n690), .ZN(new_n931));
  AOI211_X1 g506(.A(new_n920), .B(new_n929), .C1(new_n911), .C2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n905), .B2(G1384), .ZN(new_n934));
  INV_X1    g509(.A(G1384), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n843), .A2(KEYINPUT109), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT45), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT116), .B1(new_n937), .B2(new_n899), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n905), .A2(new_n933), .A3(G1384), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT109), .B1(new_n843), .B2(new_n935), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n900), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT116), .ZN(new_n942));
  NAND3_X1  g517(.A1(G160), .A2(KEYINPUT106), .A3(G40), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n896), .A2(new_n897), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n935), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT117), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n938), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n934), .A2(new_n951), .A3(new_n936), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT110), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n934), .A2(new_n954), .A3(new_n951), .A4(new_n936), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n501), .A2(new_n935), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n943), .A2(new_n944), .B1(new_n956), .B2(KEYINPUT50), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n950), .A2(new_n709), .B1(new_n958), .B2(new_n729), .ZN(new_n959));
  INV_X1    g534(.A(G8), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT123), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT123), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n941), .A2(new_n945), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n948), .B1(new_n963), .B2(KEYINPUT116), .ZN(new_n964));
  AOI21_X1  g539(.A(G1966), .B1(new_n964), .B2(new_n946), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(G2084), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n962), .B(G8), .C1(new_n965), .C2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(G168), .A2(new_n960), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(KEYINPUT51), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n961), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT124), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n961), .A2(new_n968), .A3(KEYINPUT124), .A4(new_n970), .ZN(new_n974));
  INV_X1    g549(.A(new_n959), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT51), .B(G8), .C1(new_n975), .C2(G286), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n969), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n981), .A3(new_n978), .ZN(new_n982));
  NAND2_X1  g557(.A1(G303), .A2(G8), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT55), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n843), .A2(KEYINPUT45), .A3(new_n935), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n956), .A2(new_n900), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n945), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n770), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n966), .B2(G2090), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n985), .A2(new_n990), .A3(G8), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n501), .A2(new_n951), .A3(new_n935), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n945), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT50), .B1(new_n939), .B2(new_n940), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n989), .B1(new_n995), .B2(G2090), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G8), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n984), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n991), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n773), .A2(G1976), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n934), .B(new_n936), .C1(new_n891), .C2(new_n898), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n1001), .A2(KEYINPUT111), .A3(G8), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT111), .B1(new_n1001), .B2(G8), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(G8), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1001), .A2(KEYINPUT111), .A3(G8), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(G305), .B2(G1981), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT49), .B1(new_n779), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  NAND3_X1  g589(.A1(G305), .A2(new_n1014), .A3(G1981), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1011), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1011), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1004), .A2(KEYINPUT52), .B1(new_n1009), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(G288), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1000), .B(new_n1022), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1019), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1018), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G288), .A2(new_n1021), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1023), .B(new_n1025), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT115), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n999), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n966), .A2(KEYINPUT120), .ZN(new_n1032));
  INV_X1    g607(.A(G1961), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n953), .A2(new_n1034), .A3(new_n955), .A4(new_n957), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n988), .B2(G2078), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(G2078), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n964), .A2(new_n946), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(G171), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1031), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n980), .A2(new_n982), .A3(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1009), .B(KEYINPUT113), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G288), .A2(G1976), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT114), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1047), .A2(new_n1025), .B1(new_n1012), .B2(new_n779), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n1045), .A2(new_n1048), .B1(new_n1029), .B2(new_n991), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT63), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1029), .A2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n959), .A2(new_n960), .A3(G286), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n990), .A2(G8), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n984), .ZN(new_n1054));
  AND4_X1   g629(.A1(new_n991), .A2(new_n1051), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n991), .A2(new_n998), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1020), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1029), .A2(KEYINPUT115), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1056), .B(new_n1052), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1059), .A2(KEYINPUT119), .A3(new_n1060), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1049), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n477), .A2(new_n479), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n469), .B1(new_n1067), .B2(KEYINPUT125), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(KEYINPUT125), .B2(new_n1067), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1069), .A2(G40), .A3(new_n893), .A4(new_n895), .ZN(new_n1070));
  AOI211_X1 g645(.A(new_n1037), .B(G2078), .C1(new_n1070), .C2(KEYINPUT126), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1070), .A2(KEYINPUT126), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1071), .A2(new_n986), .A3(new_n1072), .A4(new_n906), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1036), .A2(new_n1038), .A3(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(G171), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1066), .B1(new_n1042), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1066), .B1(new_n1074), .B2(G171), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(G171), .B2(new_n1041), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n1031), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n978), .B2(new_n977), .ZN(new_n1080));
  INV_X1    g655(.A(G1348), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1032), .A2(new_n1081), .A3(new_n1035), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1001), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n693), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n597), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT60), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1092), .A2(KEYINPUT122), .A3(new_n596), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1088), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(new_n1089), .A3(new_n597), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT122), .B1(new_n1092), .B2(new_n596), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1087), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1956), .B1(new_n993), .B2(new_n994), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT56), .B(G2072), .Z(new_n1099));
  NOR2_X1   g674(.A1(new_n988), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT121), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1104));
  XNOR2_X1  g679(.A(G299), .B(KEYINPUT57), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1105), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1105), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1101), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1108), .B1(new_n1112), .B2(new_n1107), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT58), .B(G1341), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1083), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n988), .A2(G1996), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n609), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(KEYINPUT59), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1110), .A2(new_n1113), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1094), .A2(new_n1097), .A3(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1107), .A2(new_n596), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1085), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1122), .A2(new_n1106), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1080), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1044), .A2(new_n1065), .A3(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(G290), .B(G1986), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n911), .B1(new_n1127), .B2(new_n928), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n1128), .B(KEYINPUT108), .Z(new_n1129));
  AND3_X1   g704(.A1(new_n1126), .A2(KEYINPUT127), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT127), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n932), .B1(new_n1130), .B2(new_n1131), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g707(.A1(new_n642), .A2(G319), .ZN(new_n1134));
  NOR3_X1   g708(.A1(G229), .A2(G227), .A3(new_n1134), .ZN(new_n1135));
  OAI211_X1 g709(.A(new_n852), .B(new_n1135), .C1(new_n887), .C2(new_n888), .ZN(G225));
  INV_X1    g710(.A(G225), .ZN(G308));
endmodule


