//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n581, new_n582, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n600, new_n601, new_n602, new_n603,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n649, new_n652, new_n654,
    new_n655, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G221), .A4(G218), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  OR2_X1    g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  NAND2_X1  g031(.A1(G113), .A2(G2104), .ZN(new_n457));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n457), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT69), .B(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n464), .A2(new_n470), .B1(new_n472), .B2(G101), .ZN(new_n473));
  INV_X1    g048(.A(new_n459), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n474), .B1(new_n471), .B2(KEYINPUT3), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G137), .A3(new_n469), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  AND2_X1   g054(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT3), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n459), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n469), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n479), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(KEYINPUT70), .A3(G124), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n483), .A2(G2105), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n487), .A2(new_n488), .B1(G136), .B2(new_n489), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n469), .C2(G112), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  AND2_X1   g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(new_n465), .B2(G114), .ZN(new_n496));
  NOR2_X1   g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n497), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT71), .A4(G2104), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n475), .A2(new_n494), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n505), .B1(new_n466), .B2(new_n468), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n504), .B1(new_n475), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n459), .B(new_n461), .C1(KEYINPUT72), .C2(new_n504), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n467), .A2(G2105), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n509), .B(G138), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n508), .B1(new_n512), .B2(new_n504), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n503), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT6), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT74), .B1(new_n517), .B2(KEYINPUT6), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(new_n525), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n522), .A2(G50), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n521), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G75), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n516), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT5), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n522), .A2(G88), .A3(new_n527), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n529), .A2(G62), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n531), .A2(new_n538), .ZN(G166));
  AND2_X1   g114(.A1(new_n532), .A2(new_n534), .ZN(new_n540));
  AND2_X1   g115(.A1(G63), .A2(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(KEYINPUT75), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n532), .A2(new_n534), .A3(new_n541), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n542), .A2(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n521), .A2(KEYINPUT6), .B1(new_n523), .B2(new_n526), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n550), .A2(G89), .A3(new_n540), .ZN(new_n551));
  INV_X1    g126(.A(G51), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(KEYINPUT76), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(KEYINPUT76), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n550), .A2(G543), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n549), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n549), .A2(new_n555), .A3(KEYINPUT77), .A4(new_n551), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(G168));
  NAND3_X1  g135(.A1(new_n522), .A2(G543), .A3(new_n527), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G52), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n540), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n521), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n522), .A2(new_n527), .A3(new_n540), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G90), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(G301));
  INV_X1    g143(.A(G301), .ZN(G171));
  NAND2_X1  g144(.A1(new_n566), .A2(G81), .ZN(new_n570));
  NAND2_X1  g145(.A1(G68), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G56), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n535), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(new_n529), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n550), .A2(G43), .A3(G543), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n570), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G860), .ZN(G153));
  AND3_X1   g153(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G36), .ZN(G176));
  NAND2_X1  g155(.A1(G1), .A2(G3), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT8), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(G188));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(G65), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(G65), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n540), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G78), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n517), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT9), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n562), .A2(KEYINPUT78), .A3(new_n590), .A4(G53), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n550), .A2(KEYINPUT78), .A3(G543), .ZN(new_n592));
  INV_X1    g167(.A(G53), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT9), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n589), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n550), .A2(G91), .A3(new_n540), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(G299));
  INV_X1    g173(.A(G168), .ZN(G286));
  NAND2_X1  g174(.A1(new_n528), .A2(new_n530), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n536), .A2(new_n537), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n540), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n603), .ZN(G303));
  NAND4_X1  g179(.A1(new_n522), .A2(G49), .A3(G543), .A4(new_n527), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n522), .A2(G87), .A3(new_n527), .A4(new_n540), .ZN(new_n606));
  OAI21_X1  g181(.A(G651), .B1(new_n540), .B2(G74), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(G288));
  INV_X1    g183(.A(G61), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT80), .B1(new_n535), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G73), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n532), .A2(new_n534), .A3(new_n612), .A4(G61), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(G86), .A2(new_n566), .B1(new_n614), .B2(new_n529), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n550), .A2(G48), .A3(G543), .ZN(new_n616));
  AOI21_X1  g191(.A(KEYINPUT81), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n529), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n550), .A2(G86), .A3(new_n540), .ZN(new_n619));
  AND4_X1   g194(.A1(KEYINPUT81), .A2(new_n618), .A3(new_n616), .A4(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n617), .A2(new_n620), .ZN(G305));
  XOR2_X1   g196(.A(KEYINPUT82), .B(G47), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n562), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n540), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(new_n521), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n566), .A2(G85), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(G290));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  OR3_X1    g203(.A1(G171), .A2(KEYINPUT83), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(KEYINPUT83), .B1(G171), .B2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n566), .A2(G92), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT10), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n566), .A2(new_n633), .A3(G92), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n561), .A2(KEYINPUT84), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n550), .A2(new_n637), .A3(G543), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n636), .A2(G54), .A3(new_n638), .ZN(new_n639));
  AOI22_X1  g214(.A1(new_n540), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(new_n517), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT85), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n639), .A2(KEYINPUT85), .A3(new_n641), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n635), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n629), .B(new_n630), .C1(new_n646), .C2(G868), .ZN(G284));
  OAI211_X1 g222(.A(new_n629), .B(new_n630), .C1(new_n646), .C2(G868), .ZN(G321));
  NAND2_X1  g223(.A1(G299), .A2(new_n628), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n628), .B2(G168), .ZN(G297));
  XNOR2_X1  g225(.A(G297), .B(KEYINPUT86), .ZN(G280));
  INV_X1    g226(.A(G559), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n646), .B1(new_n652), .B2(G860), .ZN(G148));
  NAND2_X1  g228(.A1(new_n646), .A2(new_n652), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(G868), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(G868), .B2(new_n577), .ZN(G323));
  XNOR2_X1  g231(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g232(.A1(new_n459), .A2(new_n461), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n472), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2100), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT88), .B(KEYINPUT13), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n484), .A2(G123), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n489), .A2(G135), .ZN(new_n666));
  OAI221_X1 g241(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n469), .C2(G111), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(G2096), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n669), .ZN(G156));
  XNOR2_X1  g245(.A(G2451), .B(G2454), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT16), .ZN(new_n672));
  XOR2_X1   g247(.A(G2443), .B(G2446), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1341), .B(G1348), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2427), .B(G2438), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2430), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT15), .B(G2435), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(KEYINPUT14), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n676), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G14), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G401));
  XOR2_X1   g259(.A(G2084), .B(G2090), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G2067), .B(G2678), .Z(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n687), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n689), .A2(new_n690), .A3(KEYINPUT17), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT18), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G2072), .B(G2078), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n693), .B(new_n694), .C1(new_n692), .C2(new_n688), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n694), .B2(new_n693), .ZN(new_n696));
  XNOR2_X1  g271(.A(G2096), .B(G2100), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G227));
  XOR2_X1   g273(.A(G1956), .B(G2474), .Z(new_n699));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1971), .B(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT19), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n699), .A2(new_n700), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT89), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n705), .B1(new_n708), .B2(KEYINPUT20), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n702), .A2(new_n704), .A3(new_n706), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n709), .B(new_n710), .C1(KEYINPUT20), .C2(new_n708), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1986), .B(G1996), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1981), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1991), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n713), .B(new_n716), .ZN(G229));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G26), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n484), .A2(G128), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n489), .A2(G140), .ZN(new_n721));
  OAI221_X1 g296(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n469), .C2(G116), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(new_n718), .ZN(new_n725));
  MUX2_X1   g300(.A(new_n719), .B(new_n725), .S(KEYINPUT28), .Z(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(G2067), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT31), .B(G11), .ZN(new_n729));
  INV_X1    g304(.A(G28), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT30), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT30), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n731), .A2(new_n732), .A3(new_n718), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n729), .B(new_n733), .C1(new_n668), .C2(new_n718), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n735));
  INV_X1    g310(.A(G2084), .ZN(new_n736));
  AND2_X1   g311(.A1(KEYINPUT24), .A2(G34), .ZN(new_n737));
  NOR2_X1   g312(.A1(KEYINPUT24), .A2(G34), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n737), .A2(new_n738), .A3(G29), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n477), .B2(G29), .ZN(new_n740));
  OAI22_X1  g315(.A1(new_n734), .A2(new_n735), .B1(new_n736), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G5), .A2(G16), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G171), .B2(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G1961), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT94), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(G29), .A2(G32), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n489), .A2(G141), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n484), .A2(G129), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n472), .A2(G105), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n749), .A2(new_n750), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(new_n718), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n744), .B1(new_n747), .B2(new_n755), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n741), .B(new_n756), .C1(new_n736), .C2(new_n740), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n718), .A2(G33), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n475), .A2(new_n465), .ZN(new_n759));
  INV_X1    g334(.A(G139), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n658), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n759), .A2(new_n760), .B1(new_n761), .B2(new_n469), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT25), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT93), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n758), .B1(new_n766), .B2(new_n718), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(G2072), .Z(new_n768));
  NAND2_X1  g343(.A1(G164), .A2(G29), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G27), .B2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n577), .A2(G16), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G16), .B2(G19), .ZN(new_n774));
  INV_X1    g349(.A(G1341), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n774), .A2(new_n775), .B1(new_n747), .B2(new_n755), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n771), .B2(new_n770), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n734), .A2(new_n735), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n778), .B1(new_n743), .B2(G1961), .C1(new_n774), .C2(new_n775), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n757), .A2(new_n768), .A3(new_n772), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n718), .A2(G35), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G162), .B2(new_n718), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT29), .B(G2090), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G16), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G21), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G168), .B2(new_n787), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n726), .A2(G2067), .B1(G1966), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT96), .B(KEYINPUT23), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n787), .A2(G20), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G299), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1956), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n790), .B(new_n795), .C1(G1966), .C2(new_n789), .ZN(new_n796));
  INV_X1    g371(.A(G1348), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n646), .A2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G4), .B2(G16), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n786), .B(new_n800), .C1(new_n797), .C2(new_n799), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G24), .ZN(new_n802));
  XOR2_X1   g377(.A(G290), .B(KEYINPUT92), .Z(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G16), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1986), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n484), .A2(G119), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n489), .A2(G131), .ZN(new_n807));
  NOR2_X1   g382(.A1(G95), .A2(G2105), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT91), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n809), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n806), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G29), .ZN(new_n812));
  INV_X1    g387(.A(G25), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT90), .B1(new_n813), .B2(G29), .ZN(new_n814));
  OR3_X1    g389(.A1(new_n813), .A2(KEYINPUT90), .A3(G29), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT35), .B(G1991), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(G6), .A2(G16), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G305), .B2(new_n787), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT32), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT32), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(G1981), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n787), .A2(G22), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G166), .B2(new_n787), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(G1971), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n822), .A2(G1981), .A3(new_n823), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n787), .A2(G23), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n787), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT33), .Z(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(G1976), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(G1976), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n828), .A2(G1971), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n826), .A2(new_n829), .A3(new_n830), .A4(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT34), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n805), .B(new_n819), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT36), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n839), .B(new_n840), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT36), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n846), .A2(new_n847), .A3(new_n805), .A4(new_n819), .ZN(new_n848));
  AOI211_X1 g423(.A(new_n728), .B(new_n801), .C1(new_n845), .C2(new_n848), .ZN(G311));
  AOI21_X1  g424(.A(new_n801), .B1(new_n845), .B2(new_n848), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n727), .ZN(G150));
  NAND3_X1  g426(.A1(new_n550), .A2(G93), .A3(new_n540), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  INV_X1    g428(.A(G67), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n535), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n529), .ZN(new_n856));
  INV_X1    g431(.A(G55), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n852), .B(new_n856), .C1(new_n857), .C2(new_n561), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT37), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n646), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n576), .B(new_n858), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(G860), .B1(new_n866), .B2(KEYINPUT97), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(KEYINPUT97), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n864), .A2(new_n865), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n860), .B1(new_n868), .B2(new_n869), .ZN(G145));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n668), .B(new_n477), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n492), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n811), .A2(new_n661), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n811), .A2(new_n661), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G142), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT98), .B1(new_n759), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n484), .A2(G130), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n759), .A2(KEYINPUT98), .A3(new_n877), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI221_X1 g457(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n469), .C2(G118), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n874), .A2(new_n882), .A3(new_n883), .A4(new_n875), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n885), .A2(KEYINPUT99), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT99), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n754), .B(G164), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n766), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(new_n724), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n754), .B(new_n514), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n766), .B(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n894), .A2(new_n723), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n889), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(new_n724), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n723), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n888), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n873), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n871), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI211_X1 g477(.A(KEYINPUT100), .B(new_n873), .C1(new_n896), .C2(new_n899), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n896), .A2(new_n873), .A3(new_n899), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT40), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(G395));
  NOR2_X1   g485(.A1(new_n858), .A2(G868), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n632), .A2(new_n634), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n639), .A2(KEYINPUT85), .A3(new_n641), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT85), .B1(new_n639), .B2(new_n641), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI211_X1 g490(.A(new_n596), .B(new_n589), .C1(new_n591), .C2(new_n594), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g492(.A(G299), .B(new_n912), .C1(new_n913), .C2(new_n914), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT41), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT101), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n915), .A2(new_n923), .A3(new_n916), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n863), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n654), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n919), .B2(new_n928), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(G303), .A2(new_n832), .ZN(new_n933));
  NAND2_X1  g508(.A1(G166), .A2(G288), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n933), .B(new_n934), .C1(new_n617), .C2(new_n620), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n618), .A2(new_n616), .A3(new_n619), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT81), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n615), .A2(KEYINPUT81), .A3(new_n616), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n832), .A2(new_n531), .A3(new_n538), .ZN(new_n940));
  AOI21_X1  g515(.A(G288), .B1(new_n601), .B2(new_n603), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n938), .B(new_n939), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n935), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(G290), .ZN(new_n944));
  INV_X1    g519(.A(G290), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n935), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT42), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n935), .A2(new_n942), .A3(new_n945), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n945), .B1(new_n935), .B2(new_n942), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n944), .A2(KEYINPUT102), .A3(new_n946), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n947), .B1(new_n953), .B2(KEYINPUT42), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n930), .A2(new_n931), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n932), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n954), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n930), .A2(new_n957), .A3(new_n931), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n911), .B1(new_n959), .B2(G868), .ZN(G295));
  AOI21_X1  g535(.A(new_n911), .B1(new_n959), .B2(G868), .ZN(G331));
  NAND2_X1  g536(.A1(G168), .A2(G301), .ZN(new_n962));
  NAND3_X1  g537(.A1(G171), .A2(new_n559), .A3(new_n558), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n927), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n863), .A3(new_n963), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n926), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n962), .A2(new_n863), .A3(KEYINPUT104), .A4(new_n963), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n965), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(new_n919), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT105), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n968), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT105), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n965), .A2(new_n966), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n920), .B2(new_n925), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n979), .B2(new_n973), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n980), .A3(new_n871), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT106), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n951), .A2(new_n952), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n979), .A2(new_n984), .A3(new_n973), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n919), .A2(new_n922), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n921), .A2(KEYINPUT41), .A3(new_n924), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n972), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n967), .A2(new_n919), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n953), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT107), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n988), .A2(new_n989), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n984), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n991), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n981), .A2(new_n998), .A3(KEYINPUT43), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n983), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n991), .A2(KEYINPUT43), .A3(new_n995), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n981), .A2(new_n996), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT44), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(G397));
  INV_X1    g581(.A(G1996), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n754), .B(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G2067), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n723), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n811), .A2(new_n817), .ZN(new_n1012));
  OAI22_X1  g587(.A1(new_n1011), .A2(new_n1012), .B1(G2067), .B2(new_n723), .ZN(new_n1013));
  INV_X1    g588(.A(G1384), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n514), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n473), .A2(G40), .A3(new_n476), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT125), .B(KEYINPUT46), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1019), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1021), .B1(new_n1022), .B2(G1996), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1010), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1019), .B1(new_n1024), .B2(new_n754), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1019), .B(new_n1007), .C1(KEYINPUT125), .C2(KEYINPUT46), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  XOR2_X1   g602(.A(new_n1027), .B(KEYINPUT47), .Z(new_n1028));
  NAND2_X1  g603(.A1(new_n811), .A2(new_n817), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1008), .A2(new_n1010), .A3(new_n1029), .A4(new_n1012), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n1019), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT126), .ZN(new_n1032));
  NOR2_X1   g607(.A1(G290), .A2(G1986), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1019), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT48), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1020), .B(new_n1028), .C1(new_n1032), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT63), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G303), .A2(G8), .ZN(new_n1038));
  XOR2_X1   g613(.A(new_n1038), .B(KEYINPUT55), .Z(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n512), .A2(new_n504), .ZN(new_n1041));
  INV_X1    g616(.A(new_n508), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n469), .A2(G138), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT4), .B1(new_n483), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n1046), .B2(new_n503), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n514), .A2(new_n1048), .A3(new_n1014), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1018), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OR3_X1    g627(.A1(new_n1049), .A2(new_n1052), .A3(G2090), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n514), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1017), .A2(new_n1051), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1971), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1053), .A2(new_n1054), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G8), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1054), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1040), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1018), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT108), .B1(new_n1015), .B2(KEYINPUT50), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT108), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n1065), .B(new_n1048), .C1(new_n514), .C2(new_n1014), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1063), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1058), .B1(new_n1067), .B2(G2090), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT109), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT109), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1058), .B(new_n1070), .C1(new_n1067), .C2(G2090), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(G8), .A3(new_n1039), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G8), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n832), .A2(G1976), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(KEYINPUT110), .B2(KEYINPUT52), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n832), .B2(G1976), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(KEYINPUT111), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1076), .B1(KEYINPUT110), .B2(new_n1078), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n936), .B(KEYINPUT49), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n825), .B1(new_n618), .B2(KEYINPUT112), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1081), .A2(new_n1082), .B1(new_n1085), .B2(new_n1074), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1062), .A2(new_n1072), .A3(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT115), .B(G2084), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1063), .B(new_n1088), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT116), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1065), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1015), .A2(KEYINPUT108), .A3(KEYINPUT50), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1093), .A2(new_n1094), .A3(new_n1063), .A4(new_n1088), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1055), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n514), .A2(KEYINPUT114), .A3(KEYINPUT45), .A4(new_n1014), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1097), .A2(new_n1017), .A3(new_n1051), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1966), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1090), .A2(new_n1095), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(G286), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1037), .B1(new_n1087), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1069), .A2(G8), .A3(new_n1071), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1037), .B1(new_n1107), .B2(new_n1040), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1108), .A2(new_n1072), .A3(new_n1086), .A4(new_n1104), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1107), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(new_n1039), .A3(new_n1086), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1976), .B1(new_n1085), .B2(new_n1074), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n832), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(G1981), .B2(new_n936), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1074), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1110), .A2(new_n1112), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(G168), .A2(new_n1073), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT120), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1103), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1102), .A2(new_n1119), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT51), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1103), .A2(KEYINPUT51), .A3(new_n1120), .ZN(new_n1125));
  INV_X1    g700(.A(G1961), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1067), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1017), .A2(new_n771), .A3(new_n1051), .A4(new_n1055), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1098), .A2(new_n1051), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1129), .A2(G2078), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(new_n1017), .A3(new_n1132), .A4(new_n1097), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1127), .A2(G301), .A3(new_n1130), .A4(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT124), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1067), .A2(new_n1126), .B1(new_n1129), .B2(new_n1128), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(G301), .A4(new_n1133), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1135), .A2(KEYINPUT54), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1055), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT45), .B1(new_n514), .B2(new_n1014), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1018), .A2(KEYINPUT122), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1129), .B(G2078), .C1(new_n1018), .C2(KEYINPUT122), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1052), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1145), .B(new_n1130), .C1(new_n1146), .C2(G1961), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(G171), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1124), .A2(new_n1125), .B1(new_n1139), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1133), .B(new_n1130), .C1(G1961), .C2(new_n1146), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1151), .A2(new_n1152), .A3(G171), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1152), .B1(new_n1151), .B2(G171), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1147), .A2(G171), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1150), .B1(new_n1156), .B2(KEYINPUT54), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT57), .ZN(new_n1158));
  NAND2_X1  g733(.A1(G299), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n916), .A2(KEYINPUT57), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT117), .ZN(new_n1162));
  XNOR2_X1  g737(.A(KEYINPUT56), .B(G2072), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1142), .A2(new_n1162), .A3(new_n1051), .A4(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1017), .A2(new_n1051), .A3(new_n1055), .A4(new_n1163), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT117), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(G1956), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1161), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1164), .A2(new_n1161), .A3(new_n1169), .A4(new_n1166), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1015), .A2(G2067), .A3(new_n1018), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1172), .B1(new_n1067), .B2(new_n797), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1173), .A2(new_n915), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1172), .B(new_n646), .C1(new_n1067), .C2(new_n797), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT60), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1171), .A2(KEYINPUT61), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n915), .A2(KEYINPUT60), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1171), .A2(KEYINPUT61), .B1(new_n1180), .B2(new_n1173), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1177), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(KEYINPUT118), .B(G1996), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1142), .A2(KEYINPUT119), .A3(new_n1051), .A4(new_n1183), .ZN(new_n1184));
  XOR2_X1   g759(.A(KEYINPUT58), .B(G1341), .Z(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1017), .A2(new_n1051), .A3(new_n1055), .A4(new_n1183), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT119), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1184), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT59), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1190), .A2(new_n1191), .A3(new_n577), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1191), .B1(new_n1190), .B2(new_n577), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1175), .B1(new_n1182), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT54), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1151), .A2(G171), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(KEYINPUT121), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1151), .A2(new_n1152), .A3(G171), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g775(.A(KEYINPUT123), .B(new_n1196), .C1(new_n1200), .C2(new_n1155), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1149), .A2(new_n1157), .A3(new_n1195), .A4(new_n1201), .ZN(new_n1202));
  AOI22_X1  g777(.A1(KEYINPUT51), .A2(new_n1122), .B1(new_n1103), .B2(new_n1120), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1125), .ZN(new_n1204));
  OAI21_X1  g779(.A(KEYINPUT62), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1124), .A2(new_n1206), .A3(new_n1125), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1205), .A2(new_n1200), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1202), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1087), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1117), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1030), .B1(G1986), .B2(G290), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1033), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1022), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1036), .B1(new_n1211), .B2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g790(.A(G227), .ZN(new_n1217));
  NAND3_X1  g791(.A1(new_n1217), .A2(G319), .A3(new_n683), .ZN(new_n1218));
  INV_X1    g792(.A(new_n1218), .ZN(new_n1219));
  NOR2_X1   g793(.A1(new_n1219), .A2(KEYINPUT127), .ZN(new_n1220));
  AOI21_X1  g794(.A(new_n1220), .B1(new_n904), .B2(new_n905), .ZN(new_n1221));
  AOI21_X1  g795(.A(G229), .B1(KEYINPUT127), .B2(new_n1219), .ZN(new_n1222));
  AND3_X1   g796(.A1(new_n1000), .A2(new_n1221), .A3(new_n1222), .ZN(G308));
  NAND3_X1  g797(.A1(new_n1000), .A2(new_n1221), .A3(new_n1222), .ZN(G225));
endmodule


