//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT78), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT78), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n193), .A3(new_n197), .A4(new_n194), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(G101), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT4), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n201));
  XOR2_X1   g015(.A(KEYINPUT79), .B(G101), .Z(new_n202));
  AOI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G116), .ZN(new_n206));
  INV_X1    g020(.A(G116), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n196), .A2(new_n200), .A3(G101), .A4(new_n198), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n192), .A2(G104), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n194), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n201), .A2(new_n202), .B1(G101), .B2(new_n215), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n209), .A2(new_n210), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT81), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT5), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(G113), .B1(new_n206), .B2(KEYINPUT5), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n218), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n206), .A2(KEYINPUT5), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n223), .A2(KEYINPUT81), .A3(new_n219), .A4(G113), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n216), .A2(new_n217), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n213), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT6), .ZN(new_n227));
  XNOR2_X1  g041(.A(G110), .B(G122), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n199), .A2(new_n203), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n212), .A2(new_n211), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n225), .B(new_n228), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT6), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n228), .B1(new_n213), .B2(new_n225), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n230), .B(KEYINPUT82), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n235), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT6), .A4(new_n233), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT64), .A3(G143), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(G146), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(G146), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n242), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n241), .A2(G143), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(KEYINPUT1), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G125), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n244), .A2(G146), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n249), .A2(new_n254), .A3(new_n255), .A4(G128), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n252), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n249), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n247), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n257), .B1(new_n253), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G224), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n263), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n240), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(G210), .B1(G237), .B2(G902), .ZN(new_n269));
  INV_X1    g083(.A(G902), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(KEYINPUT7), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n271), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n257), .B(new_n273), .C1(new_n253), .C2(new_n262), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n216), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n215), .A2(G101), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT79), .B(G101), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n195), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n222), .A2(new_n279), .A3(new_n217), .A4(new_n224), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n228), .B(KEYINPUT8), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n276), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n272), .A2(new_n274), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n233), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT83), .B(new_n270), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n270), .B1(new_n283), .B2(new_n284), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT83), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n268), .A2(new_n269), .A3(new_n285), .A4(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n269), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n285), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n266), .B1(new_n236), .B2(new_n239), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n188), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n264), .A2(G227), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT77), .ZN(new_n298));
  XNOR2_X1  g112(.A(G110), .B(G140), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G131), .ZN(new_n301));
  INV_X1    g115(.A(G134), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT65), .B1(new_n302), .B2(G137), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT11), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT11), .ZN(new_n305));
  OAI211_X1 g119(.A(KEYINPUT65), .B(new_n305), .C1(new_n302), .C2(G137), .ZN(new_n306));
  INV_X1    g120(.A(G137), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G134), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AND4_X1   g123(.A1(new_n301), .A2(new_n304), .A3(new_n306), .A4(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n308), .B1(new_n303), .B2(KEYINPUT11), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n301), .B1(new_n311), .B2(new_n306), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n204), .A2(new_n262), .A3(new_n212), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n252), .A2(new_n256), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(KEYINPUT10), .A3(new_n216), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n202), .A2(new_n190), .A3(new_n193), .A4(new_n194), .ZN(new_n318));
  XNOR2_X1  g132(.A(G143), .B(G146), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n256), .B1(new_n250), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n320), .A3(new_n277), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT10), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n314), .B1(new_n315), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n322), .B1(new_n252), .B2(new_n256), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n328), .A2(new_n216), .B1(new_n321), .B2(new_n322), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n204), .A2(new_n262), .A3(new_n212), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT80), .A3(new_n314), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(new_n330), .A3(new_n313), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n300), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n321), .B1(new_n316), .B2(new_n216), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n336), .A2(new_n314), .A3(KEYINPUT12), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT12), .B1(new_n336), .B2(new_n314), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n334), .ZN(new_n340));
  INV_X1    g154(.A(new_n300), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n296), .B(new_n270), .C1(new_n335), .C2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n334), .A2(new_n300), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT80), .B1(new_n331), .B2(new_n314), .ZN(new_n345));
  AOI211_X1 g159(.A(new_n326), .B(new_n313), .C1(new_n329), .C2(new_n330), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n341), .B1(new_n339), .B2(new_n340), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(G469), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n296), .A2(new_n270), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n343), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT9), .B(G234), .ZN(new_n353));
  OAI21_X1  g167(.A(G221), .B1(new_n353), .B2(G902), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n295), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT70), .ZN(new_n357));
  INV_X1    g171(.A(G140), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G125), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n253), .A2(G140), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT16), .ZN(new_n361));
  OR3_X1    g175(.A1(new_n253), .A2(KEYINPUT16), .A3(G140), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n253), .A2(KEYINPUT16), .A3(G140), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(KEYINPUT70), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n241), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n365), .ZN(new_n367));
  XNOR2_X1  g181(.A(G125), .B(G140), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n364), .B1(new_n368), .B2(KEYINPUT16), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n367), .B(G146), .C1(new_n369), .C2(new_n357), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n370), .A3(KEYINPUT71), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT71), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n372), .B(new_n241), .C1(new_n363), .C2(new_n365), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n205), .A2(G128), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n248), .A2(G119), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT24), .B(G110), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT23), .B1(new_n248), .B2(G119), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n248), .A2(G119), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n248), .A2(KEYINPUT23), .A3(G119), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n378), .B1(new_n383), .B2(G110), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n371), .A2(new_n373), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT73), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(new_n368), .B2(new_n241), .ZN(new_n387));
  AND4_X1   g201(.A1(new_n386), .A2(new_n359), .A3(new_n360), .A4(new_n241), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n363), .A2(new_n365), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n389), .B1(new_n390), .B2(G146), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT72), .ZN(new_n392));
  INV_X1    g206(.A(G110), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n381), .A2(new_n392), .A3(new_n393), .A4(new_n382), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n205), .B2(G128), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n396), .A2(new_n382), .A3(new_n393), .A4(new_n374), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n376), .A2(new_n377), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n394), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT74), .B1(new_n391), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n389), .ZN(new_n402));
  AND4_X1   g216(.A1(KEYINPUT74), .A2(new_n402), .A3(new_n400), .A4(new_n370), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n385), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT75), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT22), .B(G137), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n385), .B(new_n408), .C1(new_n401), .C2(new_n403), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT68), .B(G217), .Z(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(G234), .B2(new_n270), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT69), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G902), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n410), .A2(new_n270), .A3(new_n411), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n415), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT25), .B1(new_n418), .B2(KEYINPUT76), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n417), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n262), .B1(new_n310), .B2(new_n312), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT30), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n311), .A2(new_n301), .A3(new_n306), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n302), .A2(G137), .ZN(new_n426));
  OAI21_X1  g240(.A(G131), .B1(new_n426), .B2(new_n308), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT64), .B1(new_n241), .B2(G143), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n249), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n250), .B1(new_n242), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n256), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n425), .B(new_n427), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n423), .A2(new_n424), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n424), .B1(new_n423), .B2(new_n432), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n211), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n211), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n423), .A2(new_n436), .A3(new_n432), .ZN(new_n437));
  NOR2_X1   g251(.A1(G237), .A2(G953), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G210), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT27), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT26), .B(G101), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT66), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT66), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n437), .A2(new_n445), .A3(new_n442), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n435), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n423), .A2(new_n436), .A3(new_n432), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n436), .B1(new_n423), .B2(new_n432), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT28), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT28), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n437), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n442), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n447), .A2(KEYINPUT31), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT31), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n435), .A2(new_n444), .A3(new_n456), .A4(new_n446), .ZN(new_n457));
  AOI211_X1 g271(.A(G472), .B(G902), .C1(new_n455), .C2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n450), .A2(KEYINPUT29), .A3(new_n442), .A4(new_n452), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n270), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT67), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(KEYINPUT67), .A3(new_n270), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n450), .A2(new_n442), .A3(new_n452), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT29), .ZN(new_n465));
  INV_X1    g279(.A(new_n434), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n423), .A2(new_n424), .A3(new_n432), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n448), .B1(new_n468), .B2(new_n211), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n464), .B(new_n465), .C1(new_n469), .C2(new_n442), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n462), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n458), .A2(KEYINPUT32), .B1(G472), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n447), .A2(KEYINPUT31), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n453), .A2(new_n454), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n457), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G472), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n476), .A3(new_n270), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT32), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n422), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(G104), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n371), .A2(new_n373), .ZN(new_n484));
  INV_X1    g298(.A(G237), .ZN(new_n485));
  AND4_X1   g299(.A1(G143), .A2(new_n485), .A3(new_n264), .A4(G214), .ZN(new_n486));
  AOI21_X1  g300(.A(G143), .B1(new_n438), .B2(G214), .ZN(new_n487));
  OAI21_X1  g301(.A(G131), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n264), .A3(G214), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n244), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n438), .A2(G143), .A3(G214), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n301), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT86), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n488), .A2(new_n494), .A3(KEYINPUT86), .A4(new_n489), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n490), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n484), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n387), .ZN(new_n501));
  INV_X1    g315(.A(new_n388), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n359), .A2(new_n360), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n501), .A2(new_n502), .B1(G146), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(KEYINPUT18), .B(G131), .C1(new_n486), .C2(new_n487), .ZN(new_n505));
  NAND2_X1  g319(.A1(KEYINPUT18), .A2(G131), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n492), .A2(new_n493), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n483), .B1(new_n500), .B2(new_n510), .ZN(new_n511));
  AOI211_X1 g325(.A(new_n482), .B(new_n509), .C1(new_n484), .C2(new_n499), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n270), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT87), .B(new_n270), .C1(new_n511), .C2(new_n512), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(G475), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(G475), .A2(G902), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT19), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n368), .B(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n370), .B1(G146), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n488), .A2(new_n494), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT84), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT85), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n370), .B(new_n526), .C1(G146), .C2(new_n520), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n483), .B1(new_n528), .B2(new_n510), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n518), .B1(new_n529), .B2(new_n512), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT20), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT20), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n532), .B(new_n518), .C1(new_n529), .C2(new_n512), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n517), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n264), .A2(G952), .ZN(new_n536));
  NAND2_X1  g350(.A1(G234), .A2(G237), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(G902), .A3(G953), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT21), .B(G898), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n413), .A2(G953), .A3(new_n353), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n248), .A2(G143), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT88), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n248), .A2(G143), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n546), .B1(KEYINPUT13), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(KEYINPUT13), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT89), .ZN(new_n550));
  OAI21_X1  g364(.A(G134), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n547), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n546), .A2(new_n302), .A3(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(G116), .B(G122), .Z(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(G107), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n551), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n207), .A2(G122), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n192), .B1(new_n557), .B2(KEYINPUT14), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n558), .A2(new_n554), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n554), .ZN(new_n560));
  INV_X1    g374(.A(new_n553), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n302), .B1(new_n546), .B2(new_n552), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n559), .B(new_n560), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n544), .B1(new_n556), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n556), .A2(new_n563), .A3(new_n544), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n567), .B(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n535), .A2(new_n543), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n356), .A2(new_n480), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(new_n278), .ZN(G3));
  AND2_X1   g388(.A1(new_n352), .A2(new_n354), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n475), .A2(new_n270), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G472), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n477), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n422), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT90), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n418), .A2(KEYINPUT76), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT25), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n415), .A3(new_n419), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n577), .A2(new_n585), .A3(new_n477), .A4(new_n417), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT90), .B1(new_n355), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(KEYINPUT91), .Z(new_n589));
  INV_X1    g403(.A(new_n566), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT33), .B1(new_n590), .B2(new_n564), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n565), .A2(new_n592), .A3(new_n566), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n593), .A3(G478), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n567), .A2(new_n568), .ZN(new_n595));
  NAND2_X1  g409(.A1(G478), .A2(G902), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n517), .B2(new_n534), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n295), .A2(new_n543), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n589), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT92), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT34), .B(G104), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G6));
  AND3_X1   g417(.A1(new_n517), .A2(new_n571), .A3(new_n534), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n589), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G107), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G9));
  NOR2_X1   g421(.A1(new_n409), .A2(KEYINPUT36), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n404), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n416), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n420), .B2(new_n421), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT93), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT93), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n613), .B(new_n610), .C1(new_n420), .C2(new_n421), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n578), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n356), .A2(new_n615), .A3(new_n572), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT37), .B(G110), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G12));
  AOI22_X1  g432(.A1(new_n612), .A2(new_n614), .B1(new_n472), .B2(new_n479), .ZN(new_n619));
  INV_X1    g433(.A(new_n604), .ZN(new_n620));
  INV_X1    g434(.A(G900), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n539), .B1(new_n541), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n619), .A2(new_n356), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G128), .ZN(G30));
  XOR2_X1   g439(.A(new_n622), .B(KEYINPUT39), .Z(new_n626));
  NAND2_X1  g440(.A1(new_n575), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(KEYINPUT40), .Z(new_n628));
  NAND4_X1  g442(.A1(new_n475), .A2(KEYINPUT32), .A3(new_n476), .A4(new_n270), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n454), .B1(new_n448), .B2(new_n449), .ZN(new_n630));
  AOI21_X1  g444(.A(G902), .B1(new_n447), .B2(new_n630), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n479), .B(new_n629), .C1(new_n476), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n289), .A2(new_n293), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n635), .A2(new_n571), .A3(new_n535), .A4(new_n187), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n612), .A2(new_n614), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n628), .A2(new_n632), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G143), .ZN(G45));
  INV_X1    g454(.A(KEYINPUT95), .ZN(new_n641));
  INV_X1    g455(.A(new_n622), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n598), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n641), .B1(new_n598), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n619), .A3(new_n356), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G146), .ZN(G48));
  OAI21_X1  g461(.A(new_n334), .B1(new_n345), .B2(new_n346), .ZN(new_n648));
  INV_X1    g462(.A(new_n339), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n648), .A2(new_n341), .B1(new_n649), .B2(new_n344), .ZN(new_n650));
  OAI21_X1  g464(.A(G469), .B1(new_n650), .B2(G902), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n343), .A3(new_n652), .ZN(new_n653));
  OAI211_X1 g467(.A(KEYINPUT96), .B(G469), .C1(new_n650), .C2(G902), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n354), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT97), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n471), .A2(G472), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n479), .A2(new_n658), .A3(new_n629), .ZN(new_n659));
  INV_X1    g473(.A(new_n422), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n543), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n294), .A2(new_n662), .A3(new_n598), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT97), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n655), .A2(new_n665), .A3(new_n354), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n657), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT41), .B(G113), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G15));
  NAND3_X1  g483(.A1(new_n294), .A2(new_n604), .A3(new_n662), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n661), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n657), .A2(new_n671), .A3(new_n666), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n665), .B1(new_n655), .B2(new_n354), .ZN(new_n675));
  INV_X1    g489(.A(new_n354), .ZN(new_n676));
  AOI211_X1 g490(.A(KEYINPUT97), .B(new_n676), .C1(new_n653), .C2(new_n654), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(KEYINPUT98), .A3(new_n671), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  AND3_X1   g495(.A1(new_n655), .A2(new_n354), .A3(new_n294), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n572), .A3(new_n619), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT99), .B(G119), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G21));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n686));
  NOR2_X1   g500(.A1(G472), .A2(G902), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n457), .B1(new_n455), .B2(KEYINPUT100), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n473), .A2(KEYINPUT100), .A3(new_n474), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(G902), .B1(new_n455), .B2(new_n457), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT101), .B1(new_n691), .B2(new_n476), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n576), .A2(new_n693), .A3(G472), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n686), .B1(new_n695), .B2(new_n422), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n693), .B1(new_n576), .B2(G472), .ZN(new_n697));
  AOI211_X1 g511(.A(KEYINPUT101), .B(new_n476), .C1(new_n475), .C2(new_n270), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n699), .A2(KEYINPUT102), .A3(new_n660), .A4(new_n690), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n294), .A2(new_n571), .A3(new_n535), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n543), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n678), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  AOI21_X1  g519(.A(new_n695), .B1(new_n612), .B2(new_n614), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n682), .A2(new_n645), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G125), .ZN(G27));
  XNOR2_X1  g522(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n349), .A2(KEYINPUT103), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n347), .A2(new_n348), .A3(new_n711), .A4(G469), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n343), .A2(new_n351), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n710), .A2(new_n712), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n715), .A2(new_n716), .A3(new_n343), .A4(new_n351), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n676), .A2(new_n188), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n289), .A2(new_n293), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n480), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n597), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n535), .A2(new_n723), .A3(new_n642), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT95), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n709), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n658), .A2(new_n629), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT106), .B1(new_n477), .B2(new_n478), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n477), .A2(KEYINPUT106), .A3(new_n478), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n422), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n720), .B1(new_n714), .B2(new_n717), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n645), .A3(new_n732), .A4(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n726), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n726), .A2(new_n733), .A3(KEYINPUT107), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n301), .ZN(G33));
  NAND3_X1  g553(.A1(new_n732), .A2(new_n480), .A3(new_n623), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n347), .A2(KEYINPUT45), .A3(new_n348), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT45), .B1(new_n347), .B2(new_n348), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n296), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n350), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n742), .B(new_n343), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n750), .B(new_n350), .C1(new_n745), .C2(new_n747), .ZN(new_n752));
  INV_X1    g566(.A(new_n343), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT109), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n749), .A2(new_n750), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n751), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n354), .A3(new_n626), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n637), .A2(new_n760), .A3(new_n578), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n760), .B1(new_n637), .B2(new_n578), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n517), .A2(new_n534), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n723), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT43), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(KEYINPUT43), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n759), .B1(new_n764), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n633), .A2(new_n188), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n767), .A2(new_n768), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n772), .B(KEYINPUT44), .C1(new_n762), .C2(new_n763), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n758), .A2(new_n770), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  NAND2_X1  g589(.A1(new_n756), .A2(new_n354), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n756), .A2(new_n778), .A3(new_n354), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n771), .A2(new_n422), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n725), .A2(new_n659), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n777), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  INV_X1    g597(.A(new_n614), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n613), .B1(new_n585), .B2(new_n610), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n659), .B(new_n572), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n678), .A2(new_n664), .B1(new_n787), .B2(new_n682), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT98), .B1(new_n678), .B2(new_n671), .ZN(new_n789));
  AND4_X1   g603(.A1(KEYINPUT98), .A2(new_n657), .A3(new_n671), .A4(new_n666), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n704), .B(new_n788), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n535), .A2(new_n571), .A3(new_n622), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n721), .A2(new_n352), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n619), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n740), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n604), .A2(new_n598), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n581), .A2(new_n587), .A3(new_n599), .A4(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n572), .B(new_n356), .C1(new_n615), .C2(new_n480), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n645), .A2(new_n706), .A3(new_n732), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n795), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n791), .A2(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n726), .A2(new_n733), .A3(KEYINPUT107), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT107), .B1(new_n726), .B2(new_n733), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n356), .B(new_n619), .C1(new_n645), .C2(new_n623), .ZN(new_n805));
  INV_X1    g619(.A(new_n702), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n585), .A2(new_n354), .A3(new_n610), .A4(new_n642), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n806), .A2(new_n718), .A3(new_n632), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n805), .A2(new_n707), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n805), .A2(KEYINPUT52), .A3(new_n707), .A4(new_n809), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n801), .A2(new_n804), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n657), .A2(new_n666), .A3(new_n703), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n696), .A2(new_n700), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n667), .B(new_n683), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n799), .A2(new_n740), .A3(new_n794), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n797), .A2(new_n798), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n824), .A3(new_n680), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n734), .A2(KEYINPUT53), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n813), .A2(KEYINPUT113), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n812), .A2(KEYINPUT113), .A3(new_n813), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n817), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n801), .A2(KEYINPUT53), .A3(new_n804), .A4(new_n814), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n825), .A2(new_n738), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(KEYINPUT114), .A3(KEYINPUT53), .A4(new_n814), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n820), .B1(new_n674), .B2(new_n679), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n804), .A2(new_n838), .A3(new_n824), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n829), .A2(new_n828), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n816), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n835), .A2(new_n837), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n832), .B1(KEYINPUT54), .B2(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n819), .A2(new_n538), .A3(new_n769), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n682), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT116), .Z(new_n846));
  NAND3_X1  g660(.A1(new_n655), .A2(new_n539), .A3(new_n721), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n847), .A2(new_n422), .A3(new_n632), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n598), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n769), .A2(new_n847), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n731), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT48), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n846), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n706), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n848), .A2(new_n765), .A3(new_n597), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n635), .A2(new_n656), .A3(new_n187), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n844), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT50), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT50), .B1(new_n844), .B2(new_n857), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n777), .A2(new_n779), .B1(new_n676), .B2(new_n655), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n844), .A2(new_n771), .ZN(new_n863));
  OAI221_X1 g677(.A(new_n856), .B1(new_n860), .B2(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n864), .A2(KEYINPUT51), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(KEYINPUT51), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n853), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n843), .A2(KEYINPUT115), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n536), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT115), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n843), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(G953), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n635), .A2(new_n632), .A3(new_n766), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n660), .A2(new_n719), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT111), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n655), .B(KEYINPUT49), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT112), .Z(new_n878));
  NAND3_X1  g692(.A1(new_n869), .A2(new_n872), .A3(new_n878), .ZN(G75));
  AOI21_X1  g693(.A(new_n270), .B1(new_n817), .B2(new_n830), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n880), .B2(G210), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n240), .A2(new_n267), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n292), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT55), .Z(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n881), .A2(new_n885), .B1(G952), .B2(new_n264), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n881), .B2(new_n885), .ZN(G51));
  NOR2_X1   g701(.A1(new_n264), .A2(G952), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n817), .A2(new_n830), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT54), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n817), .A2(new_n830), .A3(new_n831), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n350), .B(KEYINPUT57), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n335), .B2(new_n342), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n880), .A2(new_n745), .A3(new_n747), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n888), .B1(new_n895), .B2(new_n896), .ZN(G54));
  NAND3_X1  g711(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n529), .A2(new_n512), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n900), .A2(new_n901), .A3(new_n888), .ZN(G60));
  INV_X1    g716(.A(KEYINPUT117), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n596), .B(KEYINPUT59), .Z(new_n904));
  NAND2_X1  g718(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n904), .B1(new_n905), .B2(new_n891), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n591), .A2(new_n593), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g723(.A(KEYINPUT117), .B(new_n907), .C1(new_n843), .C2(new_n904), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n907), .A2(new_n904), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n888), .B1(new_n892), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(G63));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT60), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n817), .B2(new_n830), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n412), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n888), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n916), .A2(KEYINPUT118), .A3(new_n609), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT118), .B1(new_n916), .B2(new_n609), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n918), .B(KEYINPUT61), .C1(new_n920), .C2(new_n919), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(G66));
  INV_X1    g739(.A(G224), .ZN(new_n926));
  OAI21_X1  g740(.A(G953), .B1(new_n542), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n791), .A2(new_n823), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(G953), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n236), .B(new_n239), .C1(G898), .C2(new_n264), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  XNOR2_X1  g745(.A(new_n520), .B(KEYINPUT119), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n468), .B(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n782), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n796), .B(KEYINPUT121), .ZN(new_n935));
  INV_X1    g749(.A(new_n627), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n935), .A2(new_n480), .A3(new_n936), .A4(new_n771), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n773), .A2(new_n354), .A3(new_n626), .A4(new_n756), .ZN(new_n938));
  INV_X1    g752(.A(new_n763), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n769), .B1(new_n939), .B2(new_n761), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n771), .B1(new_n940), .B2(KEYINPUT44), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n937), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT122), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n774), .A2(new_n944), .A3(new_n937), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n934), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n805), .A2(new_n707), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT120), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n805), .A2(new_n949), .A3(new_n707), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n639), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n951), .A2(KEYINPUT62), .A3(new_n639), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n946), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n933), .B1(new_n957), .B2(new_n264), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n774), .A2(new_n782), .A3(new_n951), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n731), .A2(new_n806), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n757), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n804), .A2(new_n740), .A3(new_n961), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n959), .A2(new_n962), .A3(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(G900), .A2(G953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n933), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n264), .B1(G227), .B2(G900), .ZN(new_n967));
  OR3_X1    g781(.A1(new_n958), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n959), .A2(new_n962), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n264), .ZN(new_n971));
  INV_X1    g785(.A(new_n965), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(KEYINPUT123), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT123), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n963), .B2(new_n965), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n969), .B(new_n967), .C1(new_n976), .C2(new_n958), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(G953), .B1(new_n946), .B2(new_n956), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n973), .B(new_n975), .C1(new_n979), .C2(new_n933), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n969), .B1(new_n980), .B2(new_n967), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n968), .B1(new_n978), .B2(new_n981), .ZN(G72));
  XNOR2_X1  g796(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n476), .A2(new_n270), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n983), .B(new_n984), .Z(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n469), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n454), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n988), .B2(new_n447), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n842), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT127), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n946), .A2(new_n928), .A3(new_n956), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n985), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(new_n442), .A3(new_n987), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n970), .A2(new_n928), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n985), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n987), .A2(new_n442), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n888), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n993), .A2(KEYINPUT126), .A3(new_n442), .A4(new_n987), .ZN(new_n1001));
  AND4_X1   g815(.A1(new_n991), .A2(new_n996), .A3(new_n1000), .A4(new_n1001), .ZN(G57));
endmodule


