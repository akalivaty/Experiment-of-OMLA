//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  AOI22_X1  g0004(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G50), .A2(G226), .ZN(new_n206));
  INV_X1    g0006(.A(G58), .ZN(new_n207));
  INV_X1    g0007(.A(G232), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  AOI21_X1  g0009(.A(new_n209), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n204), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT66), .Z(new_n220));
  INV_X1    g0020(.A(KEYINPUT0), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n204), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n220), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n207), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n231));
  INV_X1    g0031(.A(KEYINPUT65), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n232), .A2(G1), .A3(G13), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n226), .B(new_n229), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n223), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n235), .A2(KEYINPUT0), .ZN(new_n236));
  NOR4_X1   g0036(.A1(new_n224), .A2(new_n225), .A3(new_n234), .A4(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT67), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT68), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G222), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G223), .A2(G1698), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n231), .A2(new_n233), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n267), .B(new_n271), .C1(G77), .C2(new_n263), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n230), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n269), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n279), .A2(new_n274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G226), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n272), .A2(new_n277), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G190), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(G200), .ZN(new_n285));
  INV_X1    g0085(.A(G13), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G1), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n231), .A2(new_n233), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT69), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT69), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n231), .A2(new_n233), .A3(new_n293), .A4(new_n290), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n289), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G50), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n273), .B2(G20), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n295), .A2(new_n297), .B1(new_n296), .B2(new_n289), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT70), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n292), .A2(new_n294), .ZN(new_n301));
  OAI21_X1  g0101(.A(G20), .B1(new_n228), .B2(G50), .ZN(new_n302));
  INV_X1    g0102(.A(G150), .ZN(new_n303));
  NOR2_X1   g0103(.A1(G20), .A2(G33), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n226), .A2(G33), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT8), .B(G58), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n302), .B1(new_n303), .B2(new_n305), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n299), .A2(new_n300), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n300), .B1(new_n299), .B2(new_n309), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n284), .B(new_n285), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n310), .A2(new_n311), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT71), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT10), .B1(new_n285), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n282), .A2(KEYINPUT71), .A3(G200), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n316), .A2(new_n284), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n299), .A2(new_n309), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(G179), .B2(new_n282), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n282), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G238), .A2(G1698), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n263), .B(new_n327), .C1(new_n208), .C2(G1698), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(new_n271), .C1(G107), .C2(new_n263), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n276), .B1(new_n280), .B2(G244), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G200), .ZN(new_n332));
  XOR2_X1   g0132(.A(KEYINPUT15), .B(G87), .Z(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n306), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n307), .A2(new_n305), .B1(new_n226), .B2(new_n215), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n291), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n289), .A2(new_n215), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n291), .B1(new_n273), .B2(G20), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G77), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n332), .B(new_n341), .C1(new_n283), .C2(new_n331), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n320), .A2(new_n326), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n307), .B1(new_n273), .B2(G20), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n295), .A2(new_n344), .B1(new_n307), .B2(new_n289), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n256), .A2(new_n262), .A3(new_n226), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT7), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n226), .A4(new_n261), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT73), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n254), .A2(new_n255), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n352), .A2(KEYINPUT73), .A3(KEYINPUT7), .A4(new_n226), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT16), .B1(new_n355), .B2(G68), .ZN(new_n356));
  XNOR2_X1  g0156(.A(G58), .B(G68), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(G20), .B1(G159), .B2(new_n304), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT7), .B1(new_n352), .B2(new_n226), .ZN(new_n359));
  INV_X1    g0159(.A(new_n349), .ZN(new_n360));
  OAI21_X1  g0160(.A(G68), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n358), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n356), .A2(new_n358), .B1(KEYINPUT16), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n291), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n345), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT76), .B(KEYINPUT18), .ZN(new_n366));
  OAI211_X1 g0166(.A(G223), .B(new_n264), .C1(new_n254), .C2(new_n255), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT74), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n259), .A2(new_n261), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n370), .A2(KEYINPUT74), .A3(G223), .A4(new_n264), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G33), .A2(G87), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(G226), .A3(G1698), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n369), .A2(new_n371), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n271), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n279), .A2(G232), .A3(new_n274), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n375), .A2(G179), .A3(new_n277), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT75), .ZN(new_n379));
  AOI211_X1 g0179(.A(new_n276), .B(new_n376), .C1(new_n374), .C2(new_n271), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n378), .B(new_n379), .C1(new_n380), .C2(new_n323), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n375), .A2(new_n277), .A3(new_n377), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G169), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n379), .B1(new_n384), .B2(new_n378), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n365), .B(new_n366), .C1(new_n382), .C2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT76), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT18), .ZN(new_n388));
  INV_X1    g0188(.A(new_n378), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n276), .B1(new_n374), .B2(new_n271), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n323), .B1(new_n390), .B2(new_n377), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT75), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n347), .A2(new_n346), .B1(new_n351), .B2(new_n353), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n393), .B(new_n358), .C1(new_n394), .C2(new_n227), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n362), .A2(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n291), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n392), .A2(new_n381), .B1(new_n398), .B2(new_n345), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n386), .B1(new_n388), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n380), .A2(G190), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n383), .A2(G200), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n398), .A2(new_n401), .A3(new_n402), .A4(new_n345), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n364), .B1(new_n395), .B2(new_n396), .ZN(new_n406));
  INV_X1    g0206(.A(new_n345), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n408), .A2(KEYINPUT17), .A3(new_n402), .A4(new_n401), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n400), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n264), .A2(G226), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G232), .A2(G1698), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n263), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT72), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G97), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n256), .A2(new_n262), .B1(new_n413), .B2(new_n412), .ZN(new_n419));
  INV_X1    g0219(.A(new_n417), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT72), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n421), .A3(new_n271), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT13), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n276), .B1(new_n280), .B2(G238), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n423), .B1(new_n422), .B2(new_n424), .ZN(new_n426));
  OAI21_X1  g0226(.A(G169), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT14), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n425), .A2(new_n426), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G179), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT14), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(G169), .C1(new_n425), .C2(new_n426), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n227), .A2(G20), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n434), .B1(new_n306), .B2(new_n215), .C1(new_n305), .C2(new_n296), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n301), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT11), .ZN(new_n437));
  INV_X1    g0237(.A(new_n287), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(new_n434), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT12), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(G68), .B2(new_n339), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n433), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n429), .A2(G190), .ZN(new_n444));
  INV_X1    g0244(.A(new_n442), .ZN(new_n445));
  OAI21_X1  g0245(.A(G200), .B1(new_n425), .B2(new_n426), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n331), .A2(G179), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n323), .B2(new_n331), .ZN(new_n449));
  INV_X1    g0249(.A(new_n341), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n411), .A2(new_n443), .A3(new_n447), .A4(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n343), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT4), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n216), .A2(G1698), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n370), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n456), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n256), .B2(new_n262), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G283), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AND4_X1   g0262(.A1(KEYINPUT78), .A2(new_n263), .A3(G250), .A4(G1698), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n213), .B1(new_n256), .B2(new_n262), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT78), .B1(new_n464), .B2(G1698), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n270), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT5), .B(G41), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n471), .A2(new_n279), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G257), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(G274), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n468), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n454), .B(G200), .C1(new_n467), .C2(new_n477), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT68), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n260), .B1(new_n259), .B2(new_n261), .ZN(new_n480));
  OAI211_X1 g0280(.A(G250), .B(G1698), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT78), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n464), .A2(KEYINPUT78), .A3(G1698), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n460), .A3(new_n461), .A4(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n477), .B1(new_n485), .B2(new_n271), .ZN(new_n486));
  INV_X1    g0286(.A(G200), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT79), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n258), .A2(G1), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n489), .B1(new_n295), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n289), .A2(G97), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT77), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT77), .ZN(new_n495));
  INV_X1    g0295(.A(new_n493), .ZN(new_n496));
  AOI211_X1 g0296(.A(new_n490), .B(new_n289), .C1(new_n292), .C2(new_n294), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(new_n489), .ZN(new_n498));
  INV_X1    g0298(.A(G107), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(KEYINPUT6), .A3(G97), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n489), .A2(new_n499), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n500), .B1(new_n503), .B2(KEYINPUT6), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n504), .A2(G20), .B1(G77), .B2(new_n304), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n394), .B2(new_n499), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n494), .A2(new_n498), .B1(new_n291), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n486), .A2(G190), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n478), .A2(new_n488), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n494), .A2(new_n498), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n506), .A2(new_n291), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n323), .B1(new_n467), .B2(new_n477), .ZN(new_n513));
  INV_X1    g0313(.A(G179), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n486), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n512), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n226), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT80), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n212), .A2(new_n489), .A3(new_n499), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(KEYINPUT80), .A3(new_n226), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n370), .A2(new_n226), .A3(G68), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT19), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n306), .B2(new_n489), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT81), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT81), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n523), .A2(new_n529), .A3(new_n524), .A4(new_n526), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n291), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n497), .A2(new_n333), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n334), .A2(new_n289), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n216), .A2(G1698), .ZN(new_n535));
  OAI221_X1 g0335(.A(new_n535), .B1(G238), .B2(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n536));
  INV_X1    g0336(.A(G116), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n258), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n271), .ZN(new_n539));
  OAI21_X1  g0339(.A(G250), .B1(new_n469), .B2(G1), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n474), .A2(new_n540), .B1(new_n278), .B2(new_n269), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n323), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n539), .A2(new_n514), .A3(new_n542), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n534), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n487), .B1(new_n539), .B2(new_n542), .ZN(new_n547));
  AOI211_X1 g0347(.A(new_n283), .B(new_n541), .C1(new_n538), .C2(new_n271), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n497), .A2(G87), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n533), .A3(new_n531), .A4(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n509), .A2(new_n516), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT82), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT82), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n509), .A2(new_n516), .A3(new_n552), .A4(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT22), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n212), .A2(G20), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n263), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n370), .A2(new_n226), .A3(G87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT22), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n499), .A2(G20), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT23), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n226), .A2(KEYINPUT23), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT88), .B1(new_n566), .B2(new_n499), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n568), .A2(new_n499), .A3(KEYINPUT88), .A4(G20), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n563), .B(new_n565), .C1(new_n567), .C2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(KEYINPUT89), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT89), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n568), .A2(new_n499), .A3(G20), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT88), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(new_n569), .B1(KEYINPUT23), .B2(new_n564), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n573), .B1(new_n577), .B2(new_n563), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n562), .B1(new_n572), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g0379(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n571), .A2(KEYINPUT89), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(new_n573), .A3(new_n563), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n580), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n562), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(new_n291), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n497), .A2(G107), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n438), .A2(new_n564), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n589), .B(KEYINPUT25), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n213), .A2(new_n264), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n370), .B(new_n592), .C1(G257), .C2(new_n264), .ZN(new_n593));
  INV_X1    g0393(.A(G294), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n258), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n271), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n472), .A2(G264), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n476), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(G179), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n323), .B2(new_n598), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n591), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n588), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n584), .A2(new_n562), .A3(new_n585), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n585), .B1(new_n584), .B2(new_n562), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n605), .B2(new_n291), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n598), .A2(G200), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n598), .A2(new_n283), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n606), .A2(new_n590), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n537), .A2(G20), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n461), .B(new_n226), .C1(G33), .C2(new_n489), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n291), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT20), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT85), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n291), .A2(KEYINPUT20), .A3(new_n610), .A4(new_n611), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT84), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n612), .A2(KEYINPUT85), .A3(new_n613), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n616), .A2(new_n619), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n490), .A2(new_n537), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n364), .A2(new_n288), .A3(new_n623), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT83), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT83), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n287), .A2(G20), .A3(new_n537), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n622), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n256), .A2(new_n262), .A3(G303), .ZN(new_n630));
  OR2_X1    g0430(.A1(G257), .A2(G1698), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n370), .B(new_n631), .C1(G264), .C2(new_n264), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n270), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n471), .A2(G270), .A3(new_n279), .ZN(new_n634));
  INV_X1    g0434(.A(new_n476), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(new_n323), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n629), .A2(KEYINPUT21), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT21), .B1(new_n629), .B2(new_n637), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(G179), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n612), .A2(KEYINPUT85), .A3(new_n613), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT85), .B1(new_n612), .B2(new_n613), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n617), .B(KEYINPUT84), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n643), .A2(new_n644), .B1(new_n625), .B2(new_n626), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n640), .B1(new_n645), .B2(new_n628), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n638), .A2(new_n639), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n636), .A2(G190), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n648), .A2(new_n622), .A3(new_n627), .A4(new_n628), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n636), .A2(new_n487), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT86), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n629), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT86), .ZN(new_n653));
  INV_X1    g0453(.A(new_n650), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .A4(new_n648), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  AND4_X1   g0456(.A1(new_n601), .A2(new_n609), .A3(new_n647), .A4(new_n656), .ZN(new_n657));
  AND4_X1   g0457(.A1(new_n453), .A2(new_n554), .A3(new_n556), .A4(new_n657), .ZN(G372));
  NAND3_X1  g0458(.A1(new_n447), .A2(new_n450), .A3(new_n449), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n443), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT90), .ZN(new_n661));
  INV_X1    g0461(.A(new_n410), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT90), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n443), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n384), .A2(new_n378), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n406), .B2(new_n407), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT18), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n666), .B(KEYINPUT18), .C1(new_n406), .C2(new_n407), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n325), .B1(new_n672), .B2(new_n320), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n591), .A2(new_n600), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n629), .A2(new_n637), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT21), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n634), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n630), .A2(new_n632), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n678), .B(new_n476), .C1(new_n679), .C2(new_n270), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n514), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n629), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n629), .A2(KEYINPUT21), .A3(new_n637), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n677), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n674), .A2(new_n684), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n606), .A2(new_n590), .A3(new_n607), .A4(new_n608), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n685), .A2(new_n553), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n486), .A2(G169), .ZN(new_n688));
  AOI211_X1 g0488(.A(G179), .B(new_n477), .C1(new_n485), .C2(new_n271), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n688), .A2(new_n507), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT26), .B1(new_n690), .B2(new_n552), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n546), .A2(new_n551), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n516), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n546), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n453), .B1(new_n687), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n673), .A2(new_n696), .ZN(G369));
  OR3_X1    g0497(.A1(new_n438), .A2(KEYINPUT27), .A3(G20), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT27), .B1(new_n438), .B2(G20), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G343), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n652), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n684), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n647), .A2(new_n656), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(new_n704), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n591), .A2(new_n702), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n601), .B1(new_n686), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n601), .A2(new_n702), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n647), .A2(new_n702), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(new_n712), .A3(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n222), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n521), .A2(G116), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(G1), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n229), .B2(new_n723), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n728), .B(new_n703), .C1(new_n687), .C2(new_n695), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT92), .B1(new_n674), .B2(new_n684), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n509), .A2(new_n516), .A3(new_n552), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n638), .A2(new_n639), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT92), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(new_n601), .A3(new_n733), .A4(new_n682), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n730), .A2(new_n731), .A3(new_n609), .A4(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n546), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n690), .A2(KEYINPUT26), .A3(new_n552), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n692), .B1(new_n516), .B2(new_n693), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n702), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n729), .B1(new_n740), .B2(new_n728), .ZN(new_n741));
  INV_X1    g0541(.A(G330), .ZN(new_n742));
  AND4_X1   g0542(.A1(new_n539), .A2(new_n596), .A3(new_n542), .A4(new_n597), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n486), .A2(new_n681), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n486), .A2(new_n681), .A3(new_n743), .A4(KEYINPUT30), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n485), .A2(new_n271), .ZN(new_n748));
  INV_X1    g0548(.A(new_n477), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n636), .A2(G179), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n750), .A2(new_n751), .A3(new_n543), .A4(new_n598), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n746), .A2(new_n747), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT31), .B1(new_n753), .B2(new_n702), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n702), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n754), .B1(KEYINPUT91), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n702), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n757), .A2(KEYINPUT91), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n657), .A2(new_n554), .A3(new_n556), .A4(new_n703), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n742), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n741), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n727), .B1(new_n764), .B2(G1), .ZN(G364));
  OR2_X1    g0565(.A1(new_n707), .A2(G330), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n286), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n273), .B1(new_n767), .B2(G45), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n722), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n766), .A2(new_n708), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT93), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n222), .A2(G355), .A3(new_n263), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n721), .A2(new_n370), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G45), .B2(new_n229), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n252), .A2(new_n469), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n774), .B1(G116), .B2(new_n222), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n268), .B1(new_n226), .B2(G169), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT94), .Z(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n771), .B1(new_n778), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n784), .ZN(new_n787));
  INV_X1    g0587(.A(new_n263), .ZN(new_n788));
  INV_X1    g0588(.A(G303), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n487), .A2(G179), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n790), .A2(G20), .A3(G190), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n788), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT98), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n283), .A2(G20), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT96), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n797), .A2(G179), .A3(new_n487), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n797), .A2(G179), .A3(G200), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G283), .A2(new_n798), .B1(new_n799), .B2(G329), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n226), .A2(new_n514), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n801), .A2(new_n283), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  NOR4_X1   g0604(.A1(new_n226), .A2(new_n514), .A3(new_n283), .A4(new_n487), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(G326), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n792), .A2(new_n793), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n794), .A2(new_n800), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G179), .A2(G200), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n226), .B1(new_n809), .B2(G190), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n808), .B1(G294), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n801), .B(KEYINPUT95), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n813), .A2(G190), .A3(new_n487), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G322), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n813), .A2(new_n283), .A3(new_n487), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n812), .B(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT99), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n815), .A2(G58), .ZN(new_n821));
  INV_X1    g0621(.A(new_n799), .ZN(new_n822));
  INV_X1    g0622(.A(G159), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n822), .A2(KEYINPUT32), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(KEYINPUT32), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n798), .A2(G107), .ZN(new_n826));
  INV_X1    g0626(.A(new_n805), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n825), .B(new_n826), .C1(new_n296), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n818), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n824), .B(new_n828), .C1(G77), .C2(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n802), .A2(new_n227), .B1(new_n810), .B2(new_n489), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT97), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n791), .A2(new_n212), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n788), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n830), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n820), .B1(new_n821), .B2(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n786), .B1(new_n707), .B2(new_n787), .C1(new_n836), .C2(new_n780), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n773), .A2(new_n837), .ZN(G396));
  NAND2_X1  g0638(.A1(new_n647), .A2(new_n601), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n731), .A2(new_n609), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n702), .B1(new_n840), .B2(new_n739), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n342), .B1(new_n341), .B2(new_n703), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n451), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n451), .A2(new_n702), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n841), .B(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n763), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT102), .Z(new_n850));
  AOI21_X1  g0650(.A(new_n770), .B1(new_n847), .B2(new_n848), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n798), .A2(G87), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n489), .B2(new_n810), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n829), .A2(G116), .B1(G303), .B2(new_n805), .ZN(new_n855));
  INV_X1    g0655(.A(G283), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(new_n802), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT100), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n854), .B(new_n858), .C1(G311), .C2(new_n799), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n594), .B2(new_n814), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n788), .B1(new_n499), .B2(new_n791), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT101), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n810), .A2(new_n207), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n815), .A2(G143), .B1(G150), .B2(new_n803), .ZN(new_n864));
  INV_X1    g0664(.A(G137), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n864), .B1(new_n865), .B2(new_n827), .C1(new_n823), .C2(new_n818), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT34), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n791), .A2(new_n296), .ZN(new_n868));
  INV_X1    g0668(.A(new_n798), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(new_n227), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n868), .B(new_n870), .C1(G132), .C2(new_n799), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n867), .A2(new_n370), .A3(new_n871), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n860), .A2(new_n862), .B1(new_n863), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n771), .B1(new_n873), .B2(new_n781), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n781), .A2(new_n782), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n874), .B1(G77), .B2(new_n876), .C1(new_n783), .C2(new_n846), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n852), .A2(new_n877), .ZN(G384));
  INV_X1    g0678(.A(KEYINPUT107), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT106), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n755), .B1(new_n754), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n757), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(KEYINPUT106), .A3(KEYINPUT31), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n762), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n845), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n843), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n445), .A2(new_n703), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n433), .A2(KEYINPUT104), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT104), .B1(new_n433), .B2(new_n887), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n887), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n443), .A2(new_n447), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n886), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n884), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT105), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n362), .A2(new_n895), .A3(new_n393), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n361), .B(new_n358), .C1(KEYINPUT105), .C2(KEYINPUT16), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n896), .A2(new_n301), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n345), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n700), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n400), .B2(new_n410), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n666), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n403), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT37), .B1(new_n904), .B2(new_n901), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n365), .B1(new_n382), .B2(new_n385), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  INV_X1    g0707(.A(new_n700), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n406), .B2(new_n407), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n906), .A2(new_n907), .A3(new_n403), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT18), .B1(new_n365), .B2(new_n666), .ZN(new_n913));
  INV_X1    g0713(.A(new_n670), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n405), .B(new_n409), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n909), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n403), .A2(new_n667), .A3(new_n909), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n910), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT40), .B1(new_n912), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n879), .B1(new_n894), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT40), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT38), .B1(new_n902), .B2(new_n911), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n912), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n894), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT38), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n909), .B1(new_n662), .B2(new_n671), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n910), .A2(new_n919), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n911), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n924), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n933), .A2(KEYINPUT107), .A3(new_n884), .A4(new_n893), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n923), .A2(new_n927), .A3(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n453), .A2(new_n884), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(G330), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n912), .B2(new_n921), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n902), .A2(new_n911), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n928), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(KEYINPUT39), .A3(new_n932), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n443), .A2(new_n702), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n433), .A2(new_n887), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT104), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n433), .A2(KEYINPUT104), .A3(new_n887), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n892), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n703), .B(new_n846), .C1(new_n687), .C2(new_n695), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n885), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n942), .A2(new_n932), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n671), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n700), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n945), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n741), .A2(new_n453), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n673), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n957), .B(new_n959), .Z(new_n960));
  XNOR2_X1  g0760(.A(new_n938), .B(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n273), .B2(new_n767), .ZN(new_n962));
  OAI211_X1 g0762(.A(G20), .B(new_n268), .C1(new_n504), .C2(KEYINPUT35), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n537), .B(new_n963), .C1(KEYINPUT35), .C2(new_n504), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT36), .Z(new_n965));
  OAI21_X1  g0765(.A(G77), .B1(new_n207), .B2(new_n227), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n229), .A2(new_n966), .B1(G50), .B2(new_n227), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(G1), .A3(new_n286), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT103), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n962), .A2(new_n965), .A3(new_n969), .ZN(G367));
  OAI211_X1 g0770(.A(new_n509), .B(new_n516), .C1(new_n507), .C2(new_n703), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n516), .B2(new_n703), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(KEYINPUT109), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(KEYINPUT109), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n714), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT108), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n531), .A2(new_n533), .A3(new_n550), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n702), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n552), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n546), .A2(new_n980), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n978), .B(new_n984), .Z(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n976), .A2(new_n718), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT42), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n976), .A2(new_n674), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n702), .B1(new_n989), .B2(new_n516), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n986), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n985), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n985), .A2(new_n991), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n722), .B(KEYINPUT41), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n719), .A2(new_n712), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n975), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT44), .Z(new_n998));
  NOR2_X1   g0798(.A1(new_n996), .A2(new_n975), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n714), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n998), .A2(new_n715), .A3(new_n1000), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n713), .B(new_n716), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(new_n708), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n764), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n995), .B1(new_n1006), .B2(new_n764), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n992), .B(new_n993), .C1(new_n1007), .C2(new_n769), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n352), .B1(new_n814), .B2(new_n789), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n791), .ZN(new_n1010));
  AOI21_X1  g0810(.A(KEYINPUT46), .B1(new_n1010), .B2(G116), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G294), .B2(new_n803), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n798), .A2(G97), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1010), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1009), .B(new_n1015), .C1(G107), .C2(new_n811), .ZN(new_n1016));
  INV_X1    g0816(.A(G317), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n817), .B2(new_n827), .C1(new_n1017), .C2(new_n822), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n818), .A2(new_n856), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n815), .A2(G150), .B1(G143), .B2(new_n805), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n227), .B2(new_n810), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n818), .A2(new_n296), .B1(new_n823), .B2(new_n802), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT111), .Z(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1010), .A2(G58), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n215), .A2(new_n869), .B1(new_n822), .B2(new_n865), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1027), .A2(new_n788), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1018), .A2(new_n1019), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n1031));
  XNOR2_X1  g0831(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n781), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n981), .A2(new_n784), .A3(new_n982), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n775), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n785), .B1(new_n222), .B2(new_n334), .C1(new_n245), .C2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n770), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1008), .A2(new_n1037), .ZN(G387));
  OAI221_X1 g0838(.A(new_n1013), .B1(new_n215), .B2(new_n791), .C1(new_n296), .C2(new_n814), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n307), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n352), .B(new_n1039), .C1(new_n1040), .C2(new_n803), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n811), .A2(new_n333), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n805), .A2(G159), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n829), .A2(G68), .B1(G150), .B2(new_n799), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n815), .A2(G317), .B1(G311), .B2(new_n803), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n805), .A2(G322), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n789), .C2(new_n818), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT115), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT48), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n856), .B2(new_n810), .C1(new_n594), .C2(new_n791), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT49), .Z(new_n1052));
  AOI21_X1  g0852(.A(new_n370), .B1(new_n799), .B2(G326), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n537), .B2(new_n869), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1045), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n771), .B1(new_n1055), .B2(new_n781), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n713), .A2(new_n784), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n785), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n307), .A2(G50), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT113), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT50), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(KEYINPUT50), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1061), .A2(new_n1062), .A3(new_n469), .A4(new_n724), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n227), .A2(new_n215), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n775), .B1(new_n469), .B2(new_n241), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n222), .A2(new_n263), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1065), .B1(G107), .B2(new_n222), .C1(new_n724), .C2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT114), .Z(new_n1068));
  OAI211_X1 g0868(.A(new_n1056), .B(new_n1057), .C1(new_n1058), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1005), .A2(new_n769), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1005), .A2(new_n764), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1005), .A2(new_n764), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1071), .A2(new_n722), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1069), .A2(new_n1070), .A3(new_n1073), .ZN(G393));
  NAND2_X1  g0874(.A1(new_n975), .A2(new_n784), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT116), .Z(new_n1076));
  OAI21_X1  g0876(.A(new_n788), .B1(new_n818), .B2(new_n594), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n814), .A2(new_n817), .B1(new_n1017), .B2(new_n827), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT52), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n799), .A2(G322), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n826), .A3(new_n1080), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1077), .B(new_n1081), .C1(G283), .C2(new_n1010), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n537), .B2(new_n810), .C1(new_n789), .C2(new_n802), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n810), .A2(new_n215), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n814), .A2(new_n823), .B1(new_n303), .B2(new_n827), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n853), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1084), .B(new_n1087), .C1(G143), .C2(new_n799), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n803), .A2(G50), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1010), .A2(G68), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n352), .B1(new_n829), .B2(new_n1040), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n780), .B1(new_n1083), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n785), .B1(new_n489), .B2(new_n222), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n249), .B2(new_n775), .ZN(new_n1095));
  OR4_X1    g0895(.A1(new_n771), .A2(new_n1076), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n768), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n723), .B1(new_n1097), .B2(new_n1072), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1006), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(G390));
  AOI21_X1  g0901(.A(new_n944), .B1(new_n931), .B2(new_n932), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n845), .B1(new_n740), .B2(new_n843), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n950), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n755), .A2(KEYINPUT91), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(KEYINPUT31), .B2(new_n882), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n762), .A2(new_n1106), .A3(new_n759), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n890), .A2(new_n892), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1107), .A2(G330), .A3(new_n846), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n912), .A2(new_n925), .A3(new_n939), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT39), .B1(new_n931), .B2(new_n932), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n951), .A2(new_n885), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n944), .B1(new_n1114), .B2(new_n1108), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1104), .B(new_n1110), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n845), .B1(new_n841), .B2(new_n846), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1117), .A2(new_n950), .B1(new_n443), .B2(new_n702), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n940), .A2(new_n943), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n702), .B(new_n844), .C1(new_n735), .C2(new_n739), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1108), .B1(new_n1120), .B2(new_n845), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1118), .A2(new_n1119), .B1(new_n1121), .B2(new_n1102), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n884), .A2(G330), .A3(new_n893), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n453), .A2(new_n884), .A3(G330), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n673), .A2(new_n958), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1108), .B1(new_n763), .B2(new_n846), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1114), .B1(new_n1127), .B2(new_n1123), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n884), .A2(G330), .A3(new_n846), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1103), .B(new_n1109), .C1(new_n1129), .C2(new_n1108), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1126), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1124), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n723), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(G132), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n263), .B1(new_n814), .B2(new_n1136), .C1(new_n869), .C2(new_n296), .ZN(new_n1137));
  XOR2_X1   g0937(.A(KEYINPUT54), .B(G143), .Z(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n818), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(G125), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n822), .A2(new_n1141), .B1(new_n823), .B2(new_n810), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1010), .A2(G150), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT53), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1137), .A2(new_n1140), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(G128), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n827), .C1(new_n865), .C2(new_n802), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n833), .B(new_n870), .C1(G294), .C2(new_n799), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n818), .A2(new_n489), .B1(new_n499), .B2(new_n802), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT117), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n815), .A2(G116), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1084), .B(new_n263), .C1(G283), .C2(new_n805), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1148), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n780), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n771), .B(new_n1154), .C1(new_n307), .C2(new_n875), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n1113), .B2(new_n783), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1124), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n768), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1135), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(G378));
  AND4_X1   g0960(.A1(G330), .A2(new_n923), .A3(new_n927), .A4(new_n934), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n952), .A2(new_n953), .B1(new_n955), .B2(new_n700), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1163));
  AOI22_X1  g0963(.A1(KEYINPUT10), .A2(new_n312), .B1(new_n314), .B2(new_n318), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n325), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1163), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n320), .A2(new_n326), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n321), .A2(new_n908), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1165), .A2(new_n1167), .A3(new_n321), .A4(new_n908), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1162), .A2(new_n945), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1172), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n957), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1161), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n923), .A2(new_n927), .A3(G330), .A4(new_n934), .ZN(new_n1177));
  AND4_X1   g0977(.A1(new_n945), .A2(new_n954), .A3(new_n1172), .A4(new_n956), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1172), .B1(new_n1162), .B2(new_n945), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1126), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT57), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT120), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT57), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1188), .A2(new_n722), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1183), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1186), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1176), .A2(new_n1180), .A3(new_n769), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT119), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n296), .B1(new_n254), .B2(G41), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n869), .A2(new_n207), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G41), .B1(new_n803), .B2(G97), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n352), .B(new_n1196), .C1(new_n818), .C2(new_n334), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n810), .A2(new_n227), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n814), .A2(new_n499), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n799), .A2(G283), .B1(G77), .B2(new_n1010), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n537), .C2(new_n827), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT58), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n802), .A2(new_n1136), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n827), .A2(new_n1141), .B1(new_n810), .B2(new_n303), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT118), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n1010), .C2(new_n1138), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n1146), .B2(new_n814), .C1(new_n865), .C2(new_n818), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n798), .A2(G159), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G41), .B1(new_n799), .B2(G124), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1209), .A2(new_n258), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1194), .B(new_n1203), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n771), .B1(new_n1214), .B2(new_n781), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(G50), .B2(new_n876), .C1(new_n1174), .C2(new_n783), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1192), .A2(new_n1193), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1193), .B1(new_n1192), .B2(new_n1216), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1191), .A2(new_n1220), .ZN(G375));
  NAND2_X1  g1021(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n950), .A2(new_n782), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n876), .A2(G68), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n799), .A2(G128), .B1(G159), .B2(new_n1010), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT123), .Z(new_n1226));
  NAND2_X1  g1026(.A1(new_n805), .A2(G132), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1195), .B1(G150), .B2(new_n829), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1139), .A2(new_n802), .B1(new_n296), .B2(new_n810), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n352), .B(new_n1229), .C1(new_n815), .C2(G137), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1042), .B1(new_n814), .B2(new_n856), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT122), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n822), .A2(new_n789), .B1(new_n537), .B2(new_n802), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G97), .B2(new_n1010), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n263), .B1(new_n798), .B2(G77), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT121), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n805), .A2(G294), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1233), .A2(new_n1235), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n818), .A2(new_n499), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1231), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n771), .B(new_n1224), .C1(new_n1241), .C2(new_n781), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1222), .A2(new_n769), .B1(new_n1223), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1128), .A2(new_n1130), .A3(new_n1126), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n994), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1245), .B2(new_n1131), .ZN(G381));
  NOR2_X1   g1046(.A1(G375), .A2(G378), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1008), .A2(new_n1037), .A3(new_n1100), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT124), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G381), .A2(new_n1248), .A3(new_n1249), .A4(new_n1251), .ZN(G407));
  OAI211_X1 g1052(.A(G407), .B(G213), .C1(G343), .C2(new_n1248), .ZN(G409));
  INV_X1    g1053(.A(new_n1131), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT60), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1254), .B(new_n722), .C1(new_n1255), .C2(new_n1244), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1244), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(KEYINPUT60), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1243), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT125), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(G375), .A2(G378), .B1(G213), .B2(new_n701), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1183), .A2(new_n994), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1159), .A2(new_n1192), .A3(new_n1216), .A4(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1264), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT120), .B1(new_n1183), .B2(KEYINPUT57), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1188), .A2(new_n722), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(new_n1181), .A2(new_n1182), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(G378), .B1(new_n1272), .B2(new_n1219), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n701), .A2(G213), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n1264), .A3(new_n1274), .A4(new_n1267), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(KEYINPUT63), .B(new_n1263), .C1(new_n1268), .C2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1273), .A2(new_n1263), .A3(new_n1274), .A4(new_n1267), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1219), .B1(new_n1279), .B2(new_n1189), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1274), .B(new_n1267), .C1(new_n1280), .C2(new_n1159), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n701), .A2(G213), .A3(G2897), .ZN(new_n1282));
  OR3_X1    g1082(.A1(new_n1261), .A2(new_n1262), .A3(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1282), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1278), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  XOR2_X1   g1089(.A(G393), .B(G396), .Z(new_n1290));
  INV_X1    g1090(.A(new_n1249), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1100), .B1(new_n1008), .B2(new_n1037), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1290), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1292), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1290), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1295), .A3(new_n1249), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1277), .A2(new_n1288), .A3(new_n1289), .A4(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1281), .A2(KEYINPUT125), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n1285), .A3(new_n1275), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1289), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1278), .A2(KEYINPUT126), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT126), .B1(new_n1278), .B2(new_n1302), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(KEYINPUT62), .B(new_n1263), .C1(new_n1268), .C2(new_n1276), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1301), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1298), .B1(new_n1307), .B2(new_n1297), .ZN(G405));
  NAND2_X1  g1108(.A1(new_n1248), .A2(new_n1273), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1263), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1309), .B(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT127), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1293), .A2(new_n1296), .A3(KEYINPUT127), .ZN(new_n1314));
  OR2_X1    g1114(.A1(new_n1314), .A2(new_n1312), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1315), .B2(new_n1311), .ZN(G402));
endmodule


