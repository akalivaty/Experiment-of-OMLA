//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n202));
  INV_X1    g001(.A(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT24), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G169gat), .B2(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT23), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n211), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(KEYINPUT24), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n206), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n203), .A2(new_n204), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n210), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT65), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(G169gat), .B2(G176gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT23), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n213), .A2(KEYINPUT25), .A3(new_n214), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n229), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT27), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G183gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n203), .A2(KEYINPUT27), .ZN(new_n240));
  AND4_X1   g039(.A1(KEYINPUT28), .A2(new_n239), .A3(new_n240), .A4(new_n204), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(new_n203), .B2(KEYINPUT27), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT27), .B(G183gat), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n204), .B(new_n243), .C1(new_n244), .C2(new_n242), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT28), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n241), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT26), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n232), .A3(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n250), .A2(new_n214), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n206), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n247), .A2(KEYINPUT68), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n242), .B1(new_n239), .B2(new_n240), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n243), .A2(new_n204), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n246), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n241), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n249), .A2(new_n251), .B1(G183gat), .B2(G190gat), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n237), .B1(new_n254), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(G113gat), .B(G120gat), .Z(new_n264));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G127gat), .B(G134gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(KEYINPUT69), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n270), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n263), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G227gat), .ZN(new_n276));
  INV_X1    g075(.A(G233gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT68), .B1(new_n247), .B2(new_n253), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n260), .A2(new_n255), .A3(new_n261), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n281), .A2(new_n273), .A3(new_n237), .A4(new_n272), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n275), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT70), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n275), .A2(new_n285), .A3(new_n278), .A4(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT33), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT33), .B1(new_n284), .B2(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT71), .ZN(new_n293));
  XNOR2_X1  g092(.A(G15gat), .B(G43gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT72), .ZN(new_n295));
  XNOR2_X1  g094(.A(G71gat), .B(G99gat), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(new_n287), .B2(KEYINPUT32), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n291), .A2(new_n293), .A3(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n287), .B(KEYINPUT32), .C1(new_n288), .C2(new_n297), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n275), .A2(new_n282), .ZN(new_n301));
  INV_X1    g100(.A(new_n278), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n303), .A2(KEYINPUT34), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(KEYINPUT34), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT73), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n299), .A2(new_n300), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n307), .B1(new_n299), .B2(new_n300), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT36), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(KEYINPUT29), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n260), .A2(new_n261), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n237), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n234), .B1(new_n225), .B2(new_n228), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n233), .A2(new_n316), .B1(new_n219), .B2(new_n220), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n279), .B2(new_n280), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n315), .B1(new_n318), .B2(new_n311), .ZN(new_n319));
  XNOR2_X1  g118(.A(G197gat), .B(G204gat), .ZN(new_n320));
  INV_X1    g119(.A(G211gat), .ZN(new_n321));
  INV_X1    g120(.A(G218gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n320), .B1(KEYINPUT22), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G211gat), .B(G218gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT75), .B1(new_n319), .B2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n237), .B(new_n311), .C1(new_n254), .C2(new_n262), .ZN(new_n328));
  INV_X1    g127(.A(new_n315), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n331));
  INV_X1    g130(.A(new_n326), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n237), .A2(new_n314), .A3(new_n311), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n326), .B(new_n335), .C1(new_n318), .C2(new_n313), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT74), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n263), .A2(new_n312), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n326), .A4(new_n335), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(G8gat), .B(G36gat), .Z(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT76), .ZN(new_n343));
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n334), .A2(new_n341), .A3(KEYINPUT30), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT77), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n327), .A2(new_n333), .B1(new_n337), .B2(new_n340), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT30), .A4(new_n346), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n341), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n345), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n334), .A2(new_n341), .A3(new_n346), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT30), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n356), .A2(new_n355), .A3(new_n357), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n352), .B(new_n354), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G1gat), .B(G29gat), .Z(new_n361));
  XNOR2_X1  g160(.A(G57gat), .B(G85gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G141gat), .B(G148gat), .Z(new_n366));
  INV_X1    g165(.A(G155gat), .ZN(new_n367));
  INV_X1    g166(.A(G162gat), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT2), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G155gat), .B(G162gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n366), .A2(new_n371), .A3(new_n369), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n269), .A2(new_n373), .A3(new_n270), .A4(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT4), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n374), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT3), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(new_n379), .A3(new_n374), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n272), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT79), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT39), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n272), .A2(new_n377), .ZN(new_n387));
  INV_X1    g186(.A(new_n375), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n384), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n365), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(KEYINPUT39), .B2(new_n385), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT86), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT40), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n393), .B2(new_n394), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n388), .A2(KEYINPUT4), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n375), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n401), .A2(new_n381), .A3(new_n390), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n376), .A2(new_n390), .A3(new_n381), .A4(new_n399), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n365), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n396), .A2(new_n397), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n360), .A2(new_n410), .ZN(new_n411));
  AND2_X1   g210(.A1(G228gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n380), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n326), .B1(new_n413), .B2(KEYINPUT29), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT84), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n379), .B1(new_n326), .B2(KEYINPUT29), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n377), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n414), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G22gat), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n418), .B(new_n414), .C1(new_n415), .C2(new_n412), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n420), .A2(new_n422), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(G22gat), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n420), .A2(KEYINPUT85), .A3(new_n421), .A4(new_n422), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(G50gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT83), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n426), .B2(G22gat), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n429), .A2(new_n434), .B1(new_n435), .B2(new_n423), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n334), .A2(new_n341), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n338), .A2(new_n332), .A3(new_n335), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n439), .B(KEYINPUT37), .C1(new_n332), .C2(new_n319), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n345), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT38), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n353), .A2(KEYINPUT37), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n444), .A2(KEYINPUT38), .A3(new_n345), .A4(new_n438), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT6), .B1(new_n407), .B2(new_n408), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(new_n408), .B2(new_n407), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n405), .A2(KEYINPUT6), .A3(new_n365), .A4(new_n406), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n448), .A2(new_n449), .A3(new_n356), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n436), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n411), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n287), .A2(KEYINPUT32), .ZN(new_n453));
  INV_X1    g252(.A(new_n297), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n453), .B(new_n454), .C1(KEYINPUT71), .C2(new_n292), .ZN(new_n455));
  INV_X1    g254(.A(new_n293), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n300), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n306), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT36), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n304), .A2(new_n305), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n299), .A2(new_n300), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n447), .B(new_n409), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n436), .B1(new_n360), .B2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n310), .A2(new_n452), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT35), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n308), .A2(new_n309), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n360), .A2(new_n463), .A3(new_n436), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n436), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n458), .A2(new_n470), .A3(new_n461), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n354), .B1(new_n359), .B2(new_n358), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n348), .A2(new_n351), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n463), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n466), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n465), .B1(new_n469), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G15gat), .B(G22gat), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT16), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(G1gat), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n481), .B(KEYINPUT90), .C1(G1gat), .C2(new_n479), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n482), .A2(G8gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(G8gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(G71gat), .A2(G78gat), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n486), .B(KEYINPUT92), .Z(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(KEYINPUT9), .ZN(new_n488));
  XNOR2_X1  g287(.A(G57gat), .B(G64gat), .ZN(new_n489));
  OAI221_X1 g288(.A(new_n487), .B1(G71gat), .B2(G78gat), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G57gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(G64gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT9), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n494), .A2(G71gat), .A3(G78gat), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n485), .B1(KEYINPUT21), .B2(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n498), .B(KEYINPUT95), .Z(new_n499));
  NAND2_X1  g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT94), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n499), .B(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n497), .A2(KEYINPUT21), .ZN(new_n505));
  XNOR2_X1  g304(.A(G127gat), .B(G155gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G183gat), .B(G211gat), .Z(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n504), .A2(new_n509), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  INV_X1    g314(.A(G99gat), .ZN(new_n516));
  INV_X1    g315(.A(G106gat), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT8), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT98), .B(G92gat), .Z(new_n519));
  OAI211_X1 g318(.A(new_n515), .B(new_n518), .C1(G85gat), .C2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G99gat), .B(G106gat), .Z(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT99), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(KEYINPUT99), .A3(new_n521), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n520), .A2(new_n521), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n527), .A2(KEYINPUT100), .ZN(new_n528));
  INV_X1    g327(.A(G29gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT14), .ZN(new_n530));
  INV_X1    g329(.A(G36gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G43gat), .B(G50gat), .Z(new_n533));
  INV_X1    g332(.A(KEYINPUT15), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n529), .A2(KEYINPUT14), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n533), .A2(new_n534), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT89), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n542), .A2(KEYINPUT89), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n539), .A2(KEYINPUT89), .A3(new_n542), .A4(new_n540), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n527), .A2(KEYINPUT100), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n528), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n527), .A2(new_n541), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT101), .ZN(new_n551));
  NAND3_X1  g350(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n556), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n549), .B(new_n558), .C1(new_n553), .C2(new_n554), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G190gat), .B(G218gat), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT102), .ZN(new_n562));
  XOR2_X1   g361(.A(G134gat), .B(G162gat), .Z(new_n563));
  AOI21_X1  g362(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n562), .B(new_n565), .Z(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OR3_X1    g366(.A1(new_n557), .A2(new_n560), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n557), .B2(new_n560), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n513), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G113gat), .B(G141gat), .Z(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT88), .B(G197gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT11), .B(G169gat), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT12), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n485), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n547), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n485), .A2(new_n541), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT18), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n485), .B(new_n541), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n582), .B(KEYINPUT13), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(new_n584), .B2(new_n585), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n579), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n586), .A2(KEYINPUT91), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT91), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n584), .A2(new_n594), .A3(new_n585), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n590), .B(new_n578), .C1(new_n584), .C2(new_n585), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n592), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n527), .A2(KEYINPUT10), .A3(new_n497), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT103), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n497), .A2(new_n522), .A3(new_n526), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(new_n527), .B2(new_n497), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(KEYINPUT10), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n600), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n600), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n606), .A2(new_n608), .A3(new_n612), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n572), .A2(new_n599), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n478), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n463), .B(KEYINPUT104), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g421(.A(KEYINPUT16), .B(G8gat), .Z(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(new_n360), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT42), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(G8gat), .B1(new_n618), .B2(new_n474), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n625), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n626), .A2(KEYINPUT105), .A3(new_n627), .A4(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(G1325gat));
  AND3_X1   g432(.A1(new_n299), .A2(new_n300), .A3(new_n460), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n460), .B1(new_n299), .B2(new_n300), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n634), .A2(new_n635), .A3(KEYINPUT36), .ZN(new_n636));
  INV_X1    g435(.A(new_n307), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n457), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n299), .A2(new_n307), .A3(new_n300), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n459), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(G15gat), .B1(new_n618), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n634), .A2(new_n635), .ZN(new_n643));
  INV_X1    g442(.A(G15gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n642), .B1(new_n618), .B2(new_n645), .ZN(G1326gat));
  NOR2_X1   g445(.A1(new_n618), .A2(new_n470), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT43), .B(G22gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1327gat));
  NAND2_X1  g448(.A1(new_n638), .A2(new_n639), .ZN(new_n650));
  INV_X1    g449(.A(new_n358), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n356), .A2(new_n355), .A3(new_n357), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n651), .A2(new_n652), .B1(new_n353), .B2(new_n345), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n653), .A2(new_n475), .A3(new_n352), .A4(new_n470), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT35), .B1(new_n650), .B2(new_n654), .ZN(new_n655));
  NOR4_X1   g454(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT35), .A4(new_n463), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n656), .A2(new_n470), .A3(new_n461), .A4(new_n458), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n571), .B1(new_n658), .B2(new_n465), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n513), .A2(new_n599), .A3(new_n616), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n529), .A3(new_n620), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT45), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n653), .A2(new_n475), .A3(new_n352), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n665), .A2(new_n436), .B1(new_n411), .B2(new_n451), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n641), .A2(new_n666), .B1(new_n655), .B2(new_n657), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n664), .B1(new_n667), .B2(new_n571), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n478), .A2(KEYINPUT44), .A3(new_n570), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n670), .A2(new_n620), .A3(new_n660), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n663), .B1(new_n529), .B2(new_n671), .ZN(G1328gat));
  NAND4_X1  g471(.A1(new_n668), .A2(new_n360), .A3(new_n669), .A4(new_n660), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(G36gat), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n659), .A2(new_n531), .A3(new_n360), .A4(new_n660), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT46), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n675), .A2(KEYINPUT46), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT106), .ZN(G1329gat));
  INV_X1    g478(.A(G43gat), .ZN(new_n680));
  INV_X1    g479(.A(new_n641), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n668), .A2(new_n681), .A3(new_n669), .A4(new_n660), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n683), .B2(new_n682), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n661), .A2(new_n680), .A3(new_n643), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(KEYINPUT47), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n682), .A2(G43gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n686), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n691), .ZN(G1330gat));
  NAND4_X1  g491(.A1(new_n668), .A2(new_n436), .A3(new_n669), .A4(new_n660), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G50gat), .ZN(new_n694));
  INV_X1    g493(.A(G50gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n661), .A2(new_n695), .A3(new_n436), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g497(.A(new_n616), .ZN(new_n699));
  NOR4_X1   g498(.A1(new_n667), .A2(new_n598), .A3(new_n572), .A4(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n620), .B(KEYINPUT109), .Z(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n360), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT49), .B(G64gat), .Z(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n704), .B2(new_n706), .ZN(G1333gat));
  NAND2_X1  g506(.A1(new_n700), .A2(new_n681), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n634), .A2(new_n635), .A3(G71gat), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n708), .A2(G71gat), .B1(new_n700), .B2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1334gat));
  NAND2_X1  g511(.A1(new_n700), .A2(new_n436), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g513(.A1(new_n513), .A2(new_n598), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n616), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT111), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n668), .A2(new_n620), .A3(new_n669), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G85gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n478), .A2(new_n570), .A3(new_n715), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT51), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT51), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n659), .A2(new_n722), .A3(new_n715), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(G85gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n620), .A2(new_n725), .A3(new_n616), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n719), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1336gat));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n668), .A2(new_n360), .A3(new_n669), .A4(new_n717), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n731), .A2(new_n519), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n474), .A2(G92gat), .A3(new_n699), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n721), .A2(new_n723), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n731), .A2(new_n519), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n722), .A2(KEYINPUT113), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n659), .B2(new_n715), .ZN(new_n740));
  AND4_X1   g539(.A1(new_n478), .A2(new_n570), .A3(new_n715), .A4(new_n739), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n733), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n735), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n730), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n738), .A2(new_n735), .A3(new_n734), .ZN(new_n745));
  INV_X1    g544(.A(new_n739), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n720), .B(new_n746), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n747), .A2(new_n733), .B1(new_n519), .B2(new_n731), .ZN(new_n748));
  OAI211_X1 g547(.A(KEYINPUT114), .B(new_n745), .C1(new_n748), .C2(new_n735), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n744), .A2(new_n749), .ZN(G1337gat));
  AND3_X1   g549(.A1(new_n670), .A2(new_n681), .A3(new_n717), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n643), .A2(new_n516), .A3(new_n616), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n751), .A2(new_n516), .B1(new_n724), .B2(new_n752), .ZN(G1338gat));
  NOR3_X1   g552(.A1(new_n699), .A2(G106gat), .A3(new_n470), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n721), .A2(new_n723), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT116), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n668), .A2(new_n436), .A3(new_n669), .A4(new_n717), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G106gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n754), .B(KEYINPUT115), .Z(new_n761));
  AOI22_X1  g560(.A1(new_n747), .A2(new_n761), .B1(G106gat), .B2(new_n757), .ZN(new_n762));
  OAI22_X1  g561(.A1(new_n756), .A2(new_n760), .B1(new_n759), .B2(new_n762), .ZN(G1339gat));
  NAND4_X1  g562(.A1(new_n513), .A2(new_n599), .A3(new_n571), .A4(new_n699), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n601), .B(new_n766), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n604), .A2(KEYINPUT10), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n607), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n612), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(new_n768), .A3(new_n607), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n606), .A2(new_n772), .A3(KEYINPUT54), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n771), .A2(KEYINPUT55), .A3(new_n773), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n776), .A2(new_n598), .A3(new_n777), .A4(new_n615), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n582), .B1(new_n581), .B2(new_n583), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n588), .A2(new_n589), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n577), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n616), .B(new_n781), .C1(new_n597), .C2(new_n596), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n571), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n781), .B1(new_n596), .B2(new_n597), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(KEYINPUT117), .B(new_n781), .C1(new_n596), .C2(new_n597), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n570), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n776), .A2(new_n615), .A3(new_n777), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n784), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n765), .B1(new_n792), .B2(new_n512), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n471), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n620), .A2(new_n474), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(G113gat), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n797), .A2(new_n798), .A3(new_n599), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n570), .B1(new_n778), .B2(new_n782), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n789), .A2(new_n790), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n512), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n764), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n803), .A2(new_n701), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n650), .A2(new_n436), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n474), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n598), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n799), .B1(new_n809), .B2(new_n798), .ZN(G1340gat));
  INV_X1    g609(.A(G120gat), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n797), .A2(new_n811), .A3(new_n699), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n616), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n813), .B2(new_n811), .ZN(G1341gat));
  OAI21_X1  g613(.A(G127gat), .B1(new_n797), .B2(new_n512), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n512), .A2(G127gat), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n815), .B(KEYINPUT118), .C1(new_n807), .C2(new_n816), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(G1342gat));
  NAND2_X1  g620(.A1(new_n474), .A2(new_n570), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(G134gat), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n824), .A2(KEYINPUT56), .ZN(new_n825));
  OAI21_X1  g624(.A(G134gat), .B1(new_n797), .B2(new_n571), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(KEYINPUT56), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(G1343gat));
  NOR2_X1   g627(.A1(new_n681), .A2(new_n795), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n793), .B2(new_n470), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n803), .A2(KEYINPUT57), .A3(new_n436), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(G141gat), .A3(new_n598), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n681), .A2(new_n470), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n804), .A2(new_n474), .A3(new_n598), .A4(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(G141gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n835), .A2(KEYINPUT58), .A3(new_n839), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1344gat));
  AND2_X1   g643(.A1(new_n804), .A2(new_n836), .ZN(new_n845));
  INV_X1    g644(.A(G148gat), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n845), .A2(new_n846), .A3(new_n474), .A4(new_n616), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT57), .B1(new_n803), .B2(new_n436), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n831), .B(new_n470), .C1(new_n802), .C2(new_n764), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n616), .B(new_n829), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n846), .A2(KEYINPUT59), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g654(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n803), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n436), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n832), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n849), .A2(KEYINPUT121), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n616), .B(new_n829), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n856), .B1(new_n860), .B2(G148gat), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n847), .B1(new_n855), .B2(new_n861), .ZN(G1345gat));
  AOI21_X1  g661(.A(new_n367), .B1(new_n834), .B2(new_n513), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n512), .A2(G155gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n845), .A2(new_n474), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n867), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT122), .B1(new_n869), .B2(new_n863), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1346gat));
  NOR2_X1   g670(.A1(new_n822), .A2(G162gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n845), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT123), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n834), .A2(new_n570), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G162gat), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n620), .A2(new_n474), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n803), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n805), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n216), .B1(new_n880), .B2(new_n599), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n701), .A2(new_n474), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n794), .A2(G169gat), .A3(new_n598), .A4(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n881), .A2(new_n883), .ZN(G1348gat));
  NAND3_X1  g683(.A1(new_n794), .A2(new_n616), .A3(new_n882), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G176gat), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n616), .A2(new_n217), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n880), .B2(new_n887), .ZN(G1349gat));
  NAND2_X1  g687(.A1(new_n513), .A2(new_n244), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n879), .A2(new_n805), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892));
  INV_X1    g691(.A(new_n471), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n803), .A2(new_n882), .A3(new_n893), .A4(new_n513), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G183gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n892), .B1(new_n891), .B2(new_n895), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n891), .A2(new_n895), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT125), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n902), .A2(new_n896), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n900), .A2(new_n903), .ZN(G1350gat));
  NOR2_X1   g703(.A1(new_n571), .A2(G190gat), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n803), .A2(new_n805), .A3(new_n878), .A4(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT126), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n803), .A2(new_n882), .A3(new_n893), .A4(new_n570), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G190gat), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n907), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT127), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(G1351gat));
  NOR3_X1   g714(.A1(new_n681), .A2(new_n701), .A3(new_n474), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n858), .B2(new_n859), .ZN(new_n917));
  OAI21_X1  g716(.A(G197gat), .B1(new_n917), .B2(new_n599), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n879), .A2(new_n836), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n599), .A2(G197gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G1352gat));
  NOR3_X1   g720(.A1(new_n919), .A2(G204gat), .A3(new_n699), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT62), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n616), .B(new_n916), .C1(new_n858), .C2(new_n859), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G204gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1353gat));
  NAND4_X1  g725(.A1(new_n879), .A2(new_n321), .A3(new_n513), .A4(new_n836), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n513), .B(new_n916), .C1(new_n858), .C2(new_n859), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT63), .B1(new_n928), .B2(G211gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1354gat));
  OAI21_X1  g730(.A(G218gat), .B1(new_n917), .B2(new_n571), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n570), .A2(new_n322), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n919), .B2(new_n933), .ZN(G1355gat));
endmodule


