

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591;

  XNOR2_X1 U321 ( .A(n367), .B(n366), .ZN(n465) );
  XOR2_X1 U322 ( .A(n360), .B(n359), .Z(n367) );
  NOR2_X1 U323 ( .A1(n419), .A2(n540), .ZN(n420) );
  NOR2_X1 U324 ( .A1(n390), .A2(n573), .ZN(n391) );
  XNOR2_X1 U325 ( .A(n289), .B(n291), .ZN(n356) );
  XNOR2_X1 U326 ( .A(n354), .B(n371), .ZN(n289) );
  XOR2_X1 U327 ( .A(G120GAT), .B(G71GAT), .Z(n430) );
  NOR2_X1 U328 ( .A1(n476), .A2(n512), .ZN(n541) );
  XNOR2_X2 U329 ( .A(n398), .B(KEYINPUT48), .ZN(n539) );
  XOR2_X1 U330 ( .A(n386), .B(n385), .Z(n584) );
  XNOR2_X1 U331 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U332 ( .A(n357), .B(n356), .Z(n290) );
  XOR2_X1 U333 ( .A(G120GAT), .B(G71GAT), .Z(n291) );
  NAND2_X1 U334 ( .A1(n574), .A2(n573), .ZN(n292) );
  XOR2_X1 U335 ( .A(G8GAT), .B(G183GAT), .Z(n399) );
  XNOR2_X1 U336 ( .A(n416), .B(KEYINPUT121), .ZN(n417) );
  XNOR2_X1 U337 ( .A(n377), .B(n376), .ZN(n378) );
  INV_X1 U338 ( .A(KEYINPUT104), .ZN(n496) );
  XNOR2_X1 U339 ( .A(n379), .B(n378), .ZN(n381) );
  XNOR2_X1 U340 ( .A(n497), .B(n496), .ZN(n498) );
  OR2_X1 U341 ( .A1(n472), .A2(n476), .ZN(n553) );
  XNOR2_X1 U342 ( .A(n455), .B(KEYINPUT124), .ZN(n587) );
  XOR2_X1 U343 ( .A(KEYINPUT38), .B(n501), .Z(n513) );
  XNOR2_X1 U344 ( .A(n456), .B(G204GAT), .ZN(n457) );
  XNOR2_X1 U345 ( .A(n458), .B(n457), .ZN(G1353GAT) );
  XOR2_X1 U346 ( .A(G134GAT), .B(KEYINPUT77), .Z(n326) );
  XOR2_X1 U347 ( .A(KEYINPUT92), .B(G85GAT), .Z(n294) );
  XNOR2_X1 U348 ( .A(G29GAT), .B(G162GAT), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U350 ( .A(n326), .B(n295), .Z(n297) );
  NAND2_X1 U351 ( .A1(G225GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n299) );
  XNOR2_X1 U353 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n298), .B(KEYINPUT2), .ZN(n450) );
  XOR2_X1 U355 ( .A(n299), .B(n450), .Z(n301) );
  XNOR2_X1 U356 ( .A(G120GAT), .B(G57GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U358 ( .A(KEYINPUT4), .B(G148GAT), .Z(n303) );
  XNOR2_X1 U359 ( .A(KEYINPUT91), .B(KEYINPUT5), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U361 ( .A(n305), .B(n304), .Z(n313) );
  XOR2_X1 U362 ( .A(KEYINPUT83), .B(KEYINPUT0), .Z(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT82), .B(G127GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U365 ( .A(G113GAT), .B(n308), .Z(n434) );
  XOR2_X1 U366 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n310) );
  XNOR2_X1 U367 ( .A(G1GAT), .B(G141GAT), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n434), .B(n311), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n540) );
  XOR2_X1 U371 ( .A(G29GAT), .B(G43GAT), .Z(n315) );
  XNOR2_X1 U372 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n315), .B(n314), .ZN(n343) );
  XNOR2_X1 U374 ( .A(G99GAT), .B(G85GAT), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n316), .B(KEYINPUT74), .ZN(n359) );
  XNOR2_X1 U376 ( .A(n343), .B(n359), .ZN(n330) );
  XOR2_X1 U377 ( .A(G36GAT), .B(G190GAT), .Z(n402) );
  XOR2_X1 U378 ( .A(G50GAT), .B(G162GAT), .Z(n441) );
  XOR2_X1 U379 ( .A(n402), .B(n441), .Z(n318) );
  NAND2_X1 U380 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U382 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n320) );
  XNOR2_X1 U383 ( .A(G92GAT), .B(G106GAT), .ZN(n319) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U385 ( .A(n322), .B(n321), .Z(n328) );
  XOR2_X1 U386 ( .A(KEYINPUT65), .B(KEYINPUT78), .Z(n324) );
  XNOR2_X1 U387 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n323) );
  XNOR2_X1 U388 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n573) );
  INV_X1 U392 ( .A(KEYINPUT112), .ZN(n389) );
  XOR2_X1 U393 ( .A(G141GAT), .B(G22GAT), .Z(n440) );
  XOR2_X1 U394 ( .A(G113GAT), .B(G36GAT), .Z(n332) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(G50GAT), .ZN(n331) );
  XNOR2_X1 U396 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U397 ( .A(n440), .B(n333), .Z(n335) );
  NAND2_X1 U398 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n347) );
  XOR2_X1 U400 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n337) );
  XNOR2_X1 U401 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U403 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n339) );
  XNOR2_X1 U404 ( .A(G197GAT), .B(G8GAT), .ZN(n338) );
  XNOR2_X1 U405 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U406 ( .A(n341), .B(n340), .Z(n345) );
  XNOR2_X1 U407 ( .A(G1GAT), .B(KEYINPUT70), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n342), .B(G15GAT), .ZN(n382) );
  XNOR2_X1 U409 ( .A(n343), .B(n382), .ZN(n344) );
  XNOR2_X1 U410 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U411 ( .A(n347), .B(n346), .Z(n579) );
  XOR2_X1 U412 ( .A(KEYINPUT76), .B(KEYINPUT32), .Z(n349) );
  XNOR2_X1 U413 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n349), .B(n348), .ZN(n357) );
  INV_X1 U415 ( .A(KEYINPUT13), .ZN(n350) );
  NAND2_X1 U416 ( .A1(G57GAT), .A2(n350), .ZN(n353) );
  INV_X1 U417 ( .A(G57GAT), .ZN(n351) );
  NAND2_X1 U418 ( .A1(n351), .A2(KEYINPUT13), .ZN(n352) );
  NAND2_X1 U419 ( .A1(n353), .A2(n352), .ZN(n371) );
  XOR2_X1 U420 ( .A(KEYINPUT71), .B(KEYINPUT75), .Z(n354) );
  NAND2_X1 U421 ( .A1(G230GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n290), .B(n358), .ZN(n360) );
  XNOR2_X1 U423 ( .A(G176GAT), .B(G92GAT), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n361), .B(G64GAT), .ZN(n405) );
  XNOR2_X1 U425 ( .A(G204GAT), .B(KEYINPUT73), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n362), .B(G78GAT), .ZN(n363) );
  XOR2_X1 U427 ( .A(n363), .B(G106GAT), .Z(n365) );
  XNOR2_X1 U428 ( .A(G148GAT), .B(KEYINPUT72), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n447) );
  XNOR2_X1 U430 ( .A(n405), .B(n447), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n465), .B(KEYINPUT41), .ZN(n461) );
  NOR2_X1 U432 ( .A1(n579), .A2(n461), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n368), .B(KEYINPUT46), .ZN(n387) );
  XOR2_X1 U434 ( .A(KEYINPUT12), .B(G64GAT), .Z(n370) );
  XNOR2_X1 U435 ( .A(G22GAT), .B(G211GAT), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n386) );
  XOR2_X1 U437 ( .A(n371), .B(n399), .Z(n373) );
  XNOR2_X1 U438 ( .A(G127GAT), .B(G155GAT), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n379) );
  XOR2_X1 U440 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n375) );
  XNOR2_X1 U441 ( .A(G71GAT), .B(KEYINPUT80), .ZN(n374) );
  XOR2_X1 U442 ( .A(n375), .B(n374), .Z(n377) );
  NAND2_X1 U443 ( .A1(G231GAT), .A2(G233GAT), .ZN(n376) );
  INV_X1 U444 ( .A(KEYINPUT14), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n382), .B(G78GAT), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n385) );
  NOR2_X1 U448 ( .A1(n387), .A2(n584), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(KEYINPUT47), .ZN(n397) );
  INV_X1 U451 ( .A(n573), .ZN(n466) );
  XNOR2_X1 U452 ( .A(KEYINPUT36), .B(n466), .ZN(n588) );
  INV_X1 U453 ( .A(n584), .ZN(n392) );
  NOR2_X1 U454 ( .A1(n588), .A2(n392), .ZN(n393) );
  XOR2_X1 U455 ( .A(KEYINPUT45), .B(n393), .Z(n394) );
  NOR2_X1 U456 ( .A1(n465), .A2(n394), .ZN(n395) );
  NAND2_X1 U457 ( .A1(n395), .A2(n579), .ZN(n396) );
  NAND2_X1 U458 ( .A1(n397), .A2(n396), .ZN(n398) );
  XNOR2_X1 U459 ( .A(KEYINPUT93), .B(G204GAT), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U461 ( .A(n402), .B(n401), .Z(n404) );
  NAND2_X1 U462 ( .A1(G226GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n406) );
  XOR2_X1 U464 ( .A(n406), .B(n405), .Z(n415) );
  XOR2_X1 U465 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n408) );
  XNOR2_X1 U466 ( .A(G169GAT), .B(KEYINPUT85), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n410) );
  XOR2_X1 U468 ( .A(KEYINPUT86), .B(KEYINPUT18), .Z(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n435) );
  INV_X1 U470 ( .A(n435), .ZN(n413) );
  XOR2_X1 U471 ( .A(G211GAT), .B(KEYINPUT21), .Z(n412) );
  XNOR2_X1 U472 ( .A(G197GAT), .B(G218GAT), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n449) );
  XNOR2_X1 U474 ( .A(n413), .B(n449), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n506) );
  NAND2_X1 U476 ( .A1(n539), .A2(n506), .ZN(n418) );
  XOR2_X1 U477 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n416) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U479 ( .A(n420), .B(KEYINPUT64), .Z(n459) );
  XOR2_X1 U480 ( .A(G99GAT), .B(G190GAT), .Z(n422) );
  XNOR2_X1 U481 ( .A(G43GAT), .B(G134GAT), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U483 ( .A(KEYINPUT87), .B(G183GAT), .Z(n424) );
  XNOR2_X1 U484 ( .A(G15GAT), .B(G176GAT), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U486 ( .A(n426), .B(n425), .Z(n432) );
  XOR2_X1 U487 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n428) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U493 ( .A(n436), .B(n435), .Z(n574) );
  INV_X1 U494 ( .A(n574), .ZN(n533) );
  XOR2_X1 U495 ( .A(KEYINPUT90), .B(KEYINPUT22), .Z(n438) );
  XNOR2_X1 U496 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n444) );
  XOR2_X1 U498 ( .A(KEYINPUT88), .B(KEYINPUT24), .Z(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U501 ( .A(n444), .B(n443), .Z(n446) );
  NAND2_X1 U502 ( .A1(G228GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n448) );
  XOR2_X1 U504 ( .A(n448), .B(n447), .Z(n452) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n475) );
  NAND2_X1 U507 ( .A1(n533), .A2(n475), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n453), .B(KEYINPUT26), .ZN(n454) );
  XNOR2_X1 U509 ( .A(KEYINPUT96), .B(n454), .ZN(n472) );
  OR2_X1 U510 ( .A1(n459), .A2(n472), .ZN(n455) );
  INV_X1 U511 ( .A(n587), .ZN(n585) );
  NAND2_X1 U512 ( .A1(n585), .A2(n465), .ZN(n458) );
  XOR2_X1 U513 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n456) );
  NOR2_X1 U514 ( .A1(n459), .A2(n475), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT55), .ZN(n575) );
  NOR2_X2 U516 ( .A1(n575), .A2(n533), .ZN(n570) );
  INV_X1 U517 ( .A(n461), .ZN(n555) );
  NAND2_X1 U518 ( .A1(n570), .A2(n555), .ZN(n464) );
  XOR2_X1 U519 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(G176GAT), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n464), .B(n463), .ZN(G1349GAT) );
  INV_X1 U522 ( .A(n540), .ZN(n529) );
  NOR2_X1 U523 ( .A1(n579), .A2(n465), .ZN(n500) );
  XOR2_X1 U524 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n468) );
  NAND2_X1 U525 ( .A1(n584), .A2(n466), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n468), .B(n467), .ZN(n482) );
  INV_X1 U527 ( .A(n506), .ZN(n531) );
  NOR2_X1 U528 ( .A1(n531), .A2(n533), .ZN(n469) );
  NOR2_X1 U529 ( .A1(n475), .A2(n469), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n470), .B(KEYINPUT25), .ZN(n473) );
  XOR2_X1 U531 ( .A(n506), .B(KEYINPUT94), .Z(n471) );
  XNOR2_X1 U532 ( .A(KEYINPUT27), .B(n471), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n473), .A2(n553), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n474), .A2(n529), .ZN(n480) );
  XNOR2_X1 U535 ( .A(n475), .B(KEYINPUT28), .ZN(n512) );
  NAND2_X1 U536 ( .A1(n541), .A2(n533), .ZN(n477) );
  NOR2_X1 U537 ( .A1(n529), .A2(n477), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(KEYINPUT95), .ZN(n479) );
  NAND2_X1 U539 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U540 ( .A(KEYINPUT97), .B(n481), .ZN(n495) );
  NOR2_X1 U541 ( .A1(n482), .A2(n495), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n483), .B(KEYINPUT98), .ZN(n516) );
  NAND2_X1 U543 ( .A1(n500), .A2(n516), .ZN(n492) );
  NOR2_X1 U544 ( .A1(n529), .A2(n492), .ZN(n484) );
  XOR2_X1 U545 ( .A(KEYINPUT34), .B(n484), .Z(n485) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NOR2_X1 U547 ( .A1(n531), .A2(n492), .ZN(n486) );
  XOR2_X1 U548 ( .A(G8GAT), .B(n486), .Z(G1325GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n488) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U551 ( .A(n488), .B(n487), .ZN(n490) );
  NOR2_X1 U552 ( .A1(n533), .A2(n492), .ZN(n489) );
  XOR2_X1 U553 ( .A(n490), .B(n489), .Z(n491) );
  XNOR2_X1 U554 ( .A(KEYINPUT99), .B(n491), .ZN(G1326GAT) );
  INV_X1 U555 ( .A(n512), .ZN(n536) );
  NOR2_X1 U556 ( .A1(n536), .A2(n492), .ZN(n493) );
  XOR2_X1 U557 ( .A(KEYINPUT102), .B(n493), .Z(n494) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(n494), .ZN(G1327GAT) );
  NOR2_X1 U559 ( .A1(n495), .A2(n584), .ZN(n497) );
  NOR2_X1 U560 ( .A1(n588), .A2(n498), .ZN(n499) );
  XOR2_X1 U561 ( .A(KEYINPUT37), .B(n499), .Z(n528) );
  NAND2_X1 U562 ( .A1(n528), .A2(n500), .ZN(n501) );
  NAND2_X1 U563 ( .A1(n513), .A2(n540), .ZN(n505) );
  XOR2_X1 U564 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n503) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NAND2_X1 U568 ( .A1(n513), .A2(n506), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(KEYINPUT106), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(n508), .ZN(G1329GAT) );
  NAND2_X1 U571 ( .A1(n574), .A2(n513), .ZN(n510) );
  XOR2_X1 U572 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n509) );
  XNOR2_X1 U573 ( .A(G43GAT), .B(n511), .ZN(G1330GAT) );
  NAND2_X1 U574 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n514), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U576 ( .A(G50GAT), .B(n515), .ZN(G1331GAT) );
  INV_X1 U577 ( .A(n579), .ZN(n568) );
  NOR2_X1 U578 ( .A1(n568), .A2(n461), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n527), .A2(n516), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n529), .A2(n523), .ZN(n518) );
  XNOR2_X1 U581 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NOR2_X1 U584 ( .A1(n531), .A2(n523), .ZN(n520) );
  XOR2_X1 U585 ( .A(G64GAT), .B(n520), .Z(G1333GAT) );
  NOR2_X1 U586 ( .A1(n533), .A2(n523), .ZN(n521) );
  XOR2_X1 U587 ( .A(KEYINPUT110), .B(n521), .Z(n522) );
  XNOR2_X1 U588 ( .A(G71GAT), .B(n522), .ZN(G1334GAT) );
  NOR2_X1 U589 ( .A1(n536), .A2(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U592 ( .A(G78GAT), .B(n526), .Z(G1335GAT) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n535) );
  NOR2_X1 U594 ( .A1(n529), .A2(n535), .ZN(n530) );
  XOR2_X1 U595 ( .A(G85GAT), .B(n530), .Z(G1336GAT) );
  NOR2_X1 U596 ( .A1(n531), .A2(n535), .ZN(n532) );
  XOR2_X1 U597 ( .A(G92GAT), .B(n532), .Z(G1337GAT) );
  NOR2_X1 U598 ( .A1(n533), .A2(n535), .ZN(n534) );
  XOR2_X1 U599 ( .A(G99GAT), .B(n534), .Z(G1338GAT) );
  NOR2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U601 ( .A(KEYINPUT44), .B(n537), .Z(n538) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n552) );
  NAND2_X1 U604 ( .A1(n574), .A2(n541), .ZN(n542) );
  NOR2_X1 U605 ( .A1(n552), .A2(n542), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n549), .A2(n568), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U609 ( .A1(n549), .A2(n555), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n547) );
  NAND2_X1 U612 ( .A1(n549), .A2(n584), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U616 ( .A1(n549), .A2(n573), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NOR2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n564) );
  NAND2_X1 U619 ( .A1(n564), .A2(n568), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  NAND2_X1 U621 ( .A1(n564), .A2(n555), .ZN(n561) );
  XOR2_X1 U622 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT114), .Z(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  XOR2_X1 U628 ( .A(G155GAT), .B(KEYINPUT117), .Z(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n584), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1346GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n566) );
  NAND2_X1 U632 ( .A1(n564), .A2(n573), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  NAND2_X1 U635 ( .A1(n568), .A2(n570), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U637 ( .A1(n570), .A2(n584), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT122), .ZN(n572) );
  XNOR2_X1 U639 ( .A(G183GAT), .B(n572), .ZN(G1350GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n577) );
  OR2_X1 U641 ( .A1(n575), .A2(n292), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G190GAT), .B(n578), .ZN(G1351GAT) );
  NOR2_X1 U644 ( .A1(n587), .A2(n579), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n588), .A2(n587), .ZN(n590) );
  INV_X1 U652 ( .A(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U654 ( .A(n591), .B(G218GAT), .ZN(G1355GAT) );
endmodule

