//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT86), .ZN(new_n203));
  OR2_X1    g002(.A1(KEYINPUT70), .A2(G134gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT70), .A2(G134gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(G127gat), .A3(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G127gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G134gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT71), .ZN(new_n210));
  XNOR2_X1  g009(.A(G113gat), .B(G120gat), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT71), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n206), .A2(new_n213), .A3(new_n208), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n211), .A2(KEYINPUT72), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(KEYINPUT72), .ZN(new_n217));
  XNOR2_X1  g016(.A(G127gat), .B(G134gat), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT73), .B(KEYINPUT1), .Z(new_n219));
  NAND4_X1  g018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT74), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT24), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G169gat), .ZN(new_n232));
  INV_X1    g031(.A(G176gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(KEYINPUT65), .B2(KEYINPUT23), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n234), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n233), .A2(KEYINPUT23), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(new_n232), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n231), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(new_n235), .A3(new_n237), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT64), .B(G169gat), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n245), .A2(new_n234), .B1(new_n246), .B2(new_n241), .ZN(new_n247));
  OR2_X1    g046(.A1(G183gat), .A2(G190gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n248), .ZN(new_n249));
  AOI211_X1 g048(.A(KEYINPUT66), .B(KEYINPUT25), .C1(new_n247), .C2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n241), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n239), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n251), .B1(new_n253), .B2(new_n240), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n243), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(KEYINPUT68), .B(new_n243), .C1(new_n250), .C2(new_n254), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT27), .B(G183gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n223), .A2(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n261), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT26), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n226), .B1(new_n234), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT26), .B1(new_n232), .B2(new_n233), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n235), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n263), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n222), .B1(new_n259), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G227gat), .ZN(new_n273));
  INV_X1    g072(.A(G233gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT74), .B1(new_n215), .B2(new_n220), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n253), .A2(new_n240), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n253), .A2(new_n251), .A3(new_n240), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT68), .B1(new_n282), .B2(new_n243), .ZN(new_n283));
  INV_X1    g082(.A(new_n258), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n270), .B(new_n278), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n272), .A2(new_n276), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n270), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n257), .B2(new_n258), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n285), .B(new_n276), .C1(new_n289), .C2(new_n222), .ZN(new_n290));
  INV_X1    g089(.A(new_n286), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI211_X1 g093(.A(new_n288), .B(new_n277), .C1(new_n257), .C2(new_n258), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n275), .B1(new_n271), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT32), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT33), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G15gat), .B(G43gat), .Z(new_n300));
  XNOR2_X1  g099(.A(G71gat), .B(G99gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n302), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n296), .B(KEYINPUT32), .C1(new_n298), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n294), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI211_X1 g107(.A(KEYINPUT76), .B(new_n293), .C1(new_n303), .C2(new_n305), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT36), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT36), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n303), .A3(new_n305), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n294), .B1(new_n303), .B2(new_n305), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G141gat), .B(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G155gat), .ZN(new_n318));
  INV_X1    g117(.A(G162gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(KEYINPUT2), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n321), .B(new_n320), .C1(new_n316), .C2(KEYINPUT2), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n221), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n324), .A2(new_n325), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n215), .A2(new_n328), .A3(new_n220), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n326), .B2(KEYINPUT3), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT79), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n326), .A2(KEYINPUT3), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n221), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n329), .A2(new_n341), .A3(KEYINPUT4), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n342), .A3(new_n331), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n329), .A2(KEYINPUT4), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n215), .A2(new_n328), .A3(new_n345), .A4(new_n220), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n344), .A2(KEYINPUT80), .A3(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(KEYINPUT5), .B(new_n333), .C1(new_n343), .C2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n344), .A2(KEYINPUT81), .A3(new_n346), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT81), .B1(new_n344), .B2(new_n346), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n340), .B(new_n349), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G1gat), .B(G29gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT0), .ZN(new_n355));
  XNOR2_X1  g154(.A(G57gat), .B(G85gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n348), .A2(new_n352), .A3(new_n357), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n357), .B1(new_n348), .B2(new_n352), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT6), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G211gat), .A2(G218gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT22), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(G197gat), .A2(G204gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G211gat), .B(G218gat), .Z(new_n377));
  OR2_X1    g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n377), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n270), .B1(new_n283), .B2(new_n284), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n289), .A2(KEYINPUT78), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT77), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n255), .A2(new_n270), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(new_n389), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n380), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n380), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n289), .A2(KEYINPUT78), .ZN(new_n397));
  AOI211_X1 g196(.A(new_n382), .B(new_n288), .C1(new_n257), .C2(new_n258), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n388), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n392), .A2(KEYINPUT29), .A3(new_n388), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n396), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n370), .B1(new_n395), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n389), .B1(new_n383), .B2(new_n385), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n380), .B1(new_n404), .B2(new_n400), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n393), .B1(new_n386), .B2(new_n389), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n405), .B(new_n369), .C1(new_n406), .C2(new_n380), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(KEYINPUT30), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n394), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n402), .B1(new_n409), .B2(new_n396), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n369), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n366), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT31), .B(G50gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n418), .B(KEYINPUT82), .Z(new_n419));
  AOI21_X1  g218(.A(KEYINPUT29), .B1(new_n335), .B2(new_n337), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(new_n380), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n378), .A2(KEYINPUT83), .A3(new_n379), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n422), .B(new_n384), .C1(KEYINPUT83), .C2(new_n379), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n328), .B1(new_n423), .B2(new_n336), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n419), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n336), .B1(new_n396), .B2(KEYINPUT29), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n418), .B1(new_n426), .B2(new_n326), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n380), .B2(new_n420), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(G22gat), .ZN(new_n430));
  INV_X1    g229(.A(G22gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n425), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n417), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n416), .B1(new_n429), .B2(G22gat), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT84), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n425), .A2(new_n428), .A3(new_n435), .A4(new_n431), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(KEYINPUT84), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT85), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n434), .A2(new_n437), .A3(KEYINPUT85), .A4(new_n436), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n433), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n310), .B(new_n315), .C1(new_n413), .C2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT38), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n369), .B1(new_n410), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n405), .B1(new_n406), .B2(new_n380), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT37), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n445), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT88), .B1(new_n363), .B2(KEYINPUT6), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n365), .B2(KEYINPUT88), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n370), .B1(new_n448), .B2(KEYINPUT37), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n396), .B1(new_n404), .B2(new_n400), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT37), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n396), .B1(new_n390), .B2(new_n394), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n445), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n452), .B(new_n407), .C1(new_n453), .C2(new_n457), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n450), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n340), .B1(new_n350), .B2(new_n351), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT39), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n332), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n357), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT39), .B1(new_n330), .B2(new_n332), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n460), .B2(new_n332), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n359), .B1(new_n466), .B2(KEYINPUT40), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n462), .A2(new_n357), .ZN(new_n468));
  INV_X1    g267(.A(new_n465), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT40), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT87), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(new_n472), .A3(KEYINPUT40), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n467), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n408), .A2(new_n474), .A3(new_n412), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n475), .A2(new_n443), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n203), .A2(new_n444), .B1(new_n459), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n408), .A2(new_n412), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n365), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n442), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n306), .A2(new_n293), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT36), .B1(new_n481), .B2(new_n312), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n306), .A2(new_n307), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n293), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n306), .A2(new_n307), .A3(new_n294), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n482), .B1(new_n486), .B2(KEYINPUT36), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n480), .A2(KEYINPUT86), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT35), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n308), .A2(new_n309), .A3(new_n442), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(new_n413), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n442), .B1(new_n481), .B2(new_n312), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n477), .A2(new_n488), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n499), .A2(KEYINPUT95), .ZN(new_n500));
  XOR2_X1   g299(.A(G57gat), .B(G64gat), .Z(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(KEYINPUT95), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G71gat), .B(G78gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n500), .A2(new_n501), .A3(new_n504), .A4(new_n502), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G231gat), .A2(G233gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G127gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(G183gat), .B(G211gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(new_n318), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(G1gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n522), .B(new_n523), .C1(G1gat), .C2(new_n520), .ZN(new_n524));
  NOR2_X1   g323(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n524), .B(new_n525), .Z(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n508), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT21), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n513), .A2(new_n514), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n514), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n517), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n519), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n530), .B1(new_n519), .B2(new_n533), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n498), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n533), .ZN(new_n538));
  INV_X1    g337(.A(new_n530), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n497), .A3(new_n534), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT91), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  OR3_X1    g344(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n547), .A2(KEYINPUT92), .B1(G29gat), .B2(G36gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(KEYINPUT92), .B2(new_n547), .ZN(new_n549));
  XOR2_X1   g348(.A(G43gat), .B(G50gat), .Z(new_n550));
  OR2_X1    g349(.A1(new_n550), .A2(KEYINPUT90), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(KEYINPUT90), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(KEYINPUT15), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n546), .A2(new_n543), .ZN(new_n556));
  XOR2_X1   g355(.A(KEYINPUT93), .B(KEYINPUT15), .Z(new_n557));
  AOI22_X1  g356(.A1(new_n550), .A2(new_n557), .B1(G29gat), .B2(G36gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n553), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n561), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT99), .B(KEYINPUT7), .ZN(new_n565));
  NAND2_X1  g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(G85gat), .ZN(new_n570));
  INV_X1    g369(.A(G92gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(KEYINPUT8), .A2(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G99gat), .B(G106gat), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n563), .A2(new_n564), .A3(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G190gat), .B(G218gat), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n575), .ZN(new_n579));
  AND2_X1   g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n560), .A2(new_n579), .B1(KEYINPUT41), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n576), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n580), .A2(KEYINPUT41), .ZN(new_n583));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n578), .B1(new_n576), .B2(new_n581), .ZN(new_n587));
  OR3_X1    g386(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n582), .B2(new_n587), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n573), .A2(new_n574), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n573), .A2(new_n574), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n528), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  OR3_X1    g395(.A1(new_n595), .A2(KEYINPUT100), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n575), .A2(new_n508), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n598), .A2(new_n596), .A3(new_n595), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT100), .B1(new_n595), .B2(new_n596), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n592), .B(new_n597), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n595), .ZN(new_n604));
  INV_X1    g403(.A(new_n592), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n579), .A2(KEYINPUT10), .A3(new_n528), .ZN(new_n607));
  OAI211_X1 g406(.A(KEYINPUT100), .B(new_n607), .C1(new_n604), .C2(KEYINPUT10), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n608), .A2(KEYINPUT101), .A3(new_n592), .A4(new_n597), .ZN(new_n609));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  NAND4_X1  g411(.A1(new_n603), .A2(new_n606), .A3(new_n609), .A4(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n601), .A2(new_n606), .ZN(new_n615));
  INV_X1    g414(.A(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n614), .B1(new_n613), .B2(new_n617), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n542), .A2(new_n591), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G229gat), .A2(G233gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n560), .A2(new_n526), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n564), .A2(new_n527), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n562), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT18), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n563), .A2(new_n527), .A3(new_n564), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n629), .A2(KEYINPUT18), .A3(new_n623), .A4(new_n624), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n555), .A2(new_n559), .A3(new_n527), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n623), .B(KEYINPUT13), .Z(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n628), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G113gat), .B(G141gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G197gat), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT11), .B(G169gat), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT89), .B(KEYINPUT12), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n628), .A2(new_n630), .A3(new_n643), .A4(new_n634), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n622), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n202), .B1(new_n496), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n443), .B1(new_n478), .B2(new_n365), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n310), .A2(new_n315), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n203), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n459), .A2(new_n476), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n488), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n492), .A2(new_n495), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n646), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(KEYINPUT103), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n647), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n366), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  INV_X1    g458(.A(new_n478), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT16), .B(G8gat), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT103), .B1(new_n654), .B2(new_n655), .ZN(new_n663));
  AOI211_X1 g462(.A(new_n202), .B(new_n646), .C1(new_n652), .C2(new_n653), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n660), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(G8gat), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n657), .B2(new_n660), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670));
  AOI211_X1 g469(.A(new_n478), .B(new_n661), .C1(new_n647), .C2(new_n656), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n670), .B1(new_n671), .B2(KEYINPUT42), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n665), .A2(KEYINPUT104), .A3(new_n668), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(G1325gat));
  NOR2_X1   g473(.A1(new_n663), .A2(new_n664), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n313), .A2(new_n314), .ZN(new_n676));
  OR3_X1    g475(.A1(new_n675), .A2(G15gat), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G15gat), .B1(new_n675), .B2(new_n487), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1326gat));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n657), .B2(new_n442), .ZN(new_n683));
  AOI211_X1 g482(.A(KEYINPUT105), .B(new_n443), .C1(new_n647), .C2(new_n656), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT105), .B1(new_n675), .B2(new_n443), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n657), .A2(new_n682), .A3(new_n442), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n687), .A3(new_n680), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n688), .ZN(G1327gat));
  AOI21_X1  g488(.A(new_n590), .B1(new_n652), .B2(new_n653), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n537), .A2(new_n541), .ZN(new_n691));
  INV_X1    g490(.A(new_n644), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n626), .A2(new_n627), .B1(new_n632), .B2(new_n633), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n643), .B1(new_n693), .B2(new_n630), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n691), .A2(new_n695), .A3(new_n621), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(G29gat), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n698), .A3(new_n366), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n450), .A2(new_n458), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n475), .A2(new_n443), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n495), .ZN(new_n704));
  OAI22_X1  g503(.A1(new_n703), .A2(new_n444), .B1(new_n491), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT44), .B1(new_n705), .B2(new_n591), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n690), .B2(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n696), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n365), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n700), .A2(new_n709), .ZN(G1328gat));
  INV_X1    g509(.A(G36gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n697), .A2(new_n711), .A3(new_n660), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n712), .A2(KEYINPUT46), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n708), .B2(new_n478), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(KEYINPUT46), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(G1329gat));
  NAND3_X1  g515(.A1(new_n654), .A2(KEYINPUT44), .A3(new_n591), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n705), .A2(new_n591), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n717), .A2(new_n649), .A3(new_n696), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n723), .A3(new_n649), .A4(new_n696), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n724), .A3(G43gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n690), .A2(new_n696), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n726), .A2(G43gat), .A3(new_n676), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n721), .A2(G43gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n728), .B1(new_n731), .B2(new_n727), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(G1330gat));
  INV_X1    g532(.A(G50gat), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n443), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n707), .A2(new_n696), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n726), .B2(new_n443), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g538(.A(new_n621), .ZN(new_n740));
  NOR4_X1   g539(.A1(new_n542), .A2(new_n645), .A3(new_n740), .A4(new_n591), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n705), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n366), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT107), .B(G57gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1332gat));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n660), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n747));
  XOR2_X1   g546(.A(KEYINPUT49), .B(G64gat), .Z(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n746), .B2(new_n748), .ZN(G1333gat));
  NAND4_X1  g548(.A1(new_n705), .A2(G71gat), .A3(new_n649), .A4(new_n741), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT108), .Z(new_n751));
  INV_X1    g550(.A(G71gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n705), .A2(new_n741), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n676), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT50), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n751), .A2(new_n757), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1334gat));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n442), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g560(.A1(new_n691), .A2(new_n645), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n705), .A2(new_n591), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n705), .A2(KEYINPUT51), .A3(new_n591), .A4(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n767), .A2(new_n570), .A3(new_n366), .A4(new_n621), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n691), .A2(new_n645), .A3(new_n740), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n707), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(new_n366), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n771), .B2(new_n570), .ZN(G1336gat));
  NAND4_X1  g571(.A1(new_n717), .A2(new_n660), .A3(new_n720), .A4(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G92gat), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n767), .A2(new_n571), .A3(new_n660), .A4(new_n621), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT52), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n774), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1337gat));
  NAND2_X1  g579(.A1(new_n770), .A2(new_n649), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G99gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n676), .A2(new_n740), .A3(G99gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1338gat));
  NAND4_X1  g584(.A1(new_n717), .A2(new_n442), .A3(new_n720), .A4(new_n769), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n740), .A2(G106gat), .A3(new_n443), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n767), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n791));
  XNOR2_X1  g590(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n767), .B2(new_n788), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n787), .A2(new_n793), .A3(KEYINPUT110), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT110), .B1(new_n787), .B2(new_n793), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(G1339gat));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n605), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(new_n603), .A3(new_n609), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n608), .A2(new_n797), .A3(new_n592), .A4(new_n597), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n616), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n613), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(KEYINPUT111), .A3(new_n613), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n800), .A2(new_n802), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n806), .A2(new_n645), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n633), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n624), .A2(new_n631), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n623), .B1(new_n629), .B2(new_n624), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n639), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n644), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n621), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n591), .B1(new_n811), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n588), .A3(new_n589), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT111), .B1(new_n803), .B2(new_n613), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n810), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n542), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n691), .A2(new_n695), .A3(new_n590), .A4(new_n740), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n365), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n827), .A2(new_n478), .A3(new_n490), .ZN(new_n828));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n645), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n826), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(new_n493), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n366), .A3(new_n478), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n645), .A2(G113gat), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n829), .B1(new_n835), .B2(new_n836), .ZN(G1340gat));
  AOI21_X1  g636(.A(G120gat), .B1(new_n828), .B2(new_n621), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n621), .A2(G120gat), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n835), .B2(new_n839), .ZN(G1341gat));
  OAI21_X1  g639(.A(G127gat), .B1(new_n834), .B2(new_n542), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n828), .A2(new_n207), .A3(new_n691), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1342gat));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n204), .A3(new_n205), .A4(new_n591), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT56), .Z(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n834), .B2(new_n590), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1343gat));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n848), .A3(new_n442), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n649), .A2(new_n365), .A3(new_n660), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT55), .B1(new_n800), .B2(new_n802), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n804), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n810), .A2(KEYINPUT114), .A3(new_n613), .A4(new_n803), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n645), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n591), .B1(new_n855), .B2(new_n819), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n542), .B1(new_n856), .B2(new_n824), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n443), .B1(new_n857), .B2(new_n826), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n849), .B(new_n850), .C1(new_n848), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n645), .A2(G141gat), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n487), .A2(new_n442), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n660), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n827), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n695), .ZN(new_n864));
  OAI22_X1  g663(.A1(new_n859), .A2(new_n860), .B1(new_n864), .B2(G141gat), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT58), .ZN(G1344gat));
  OR3_X1    g667(.A1(new_n859), .A2(KEYINPUT59), .A3(new_n740), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  INV_X1    g669(.A(new_n863), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n621), .ZN(new_n872));
  NOR4_X1   g671(.A1(new_n542), .A2(new_n645), .A3(new_n591), .A4(new_n621), .ZN(new_n873));
  INV_X1    g672(.A(new_n824), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n817), .A2(new_n644), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n619), .A3(new_n620), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n804), .A2(new_n852), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n695), .B1(new_n877), .B2(KEYINPUT114), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n878), .B2(new_n853), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n874), .B1(new_n879), .B2(new_n591), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n873), .B1(new_n880), .B2(new_n542), .ZN(new_n881));
  OAI211_X1 g680(.A(KEYINPUT116), .B(new_n848), .C1(new_n881), .C2(new_n443), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n858), .B2(KEYINPUT57), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n830), .A2(KEYINPUT57), .A3(new_n442), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n886), .A2(new_n621), .A3(new_n850), .ZN(new_n887));
  NAND2_X1  g686(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n888));
  OAI221_X1 g687(.A(new_n869), .B1(G148gat), .B2(new_n872), .C1(new_n887), .C2(new_n888), .ZN(G1345gat));
  AOI21_X1  g688(.A(G155gat), .B1(new_n871), .B2(new_n691), .ZN(new_n890));
  INV_X1    g689(.A(new_n859), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n691), .A2(G155gat), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT117), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(G1346gat));
  OAI21_X1  g693(.A(G162gat), .B1(new_n859), .B2(new_n590), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n871), .A2(new_n319), .A3(new_n591), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT118), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n478), .A2(new_n366), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT120), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n831), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n695), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n366), .B1(new_n825), .B2(new_n826), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n660), .A2(new_n490), .A3(KEYINPUT119), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  INV_X1    g704(.A(new_n490), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(new_n478), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n246), .A3(new_n645), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n902), .A2(new_n909), .ZN(G1348gat));
  OAI21_X1  g709(.A(G176gat), .B1(new_n901), .B2(new_n740), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(new_n233), .A3(new_n621), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1349gat));
  OAI21_X1  g712(.A(G183gat), .B1(new_n901), .B2(new_n542), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n908), .A2(new_n260), .A3(new_n691), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(KEYINPUT121), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n919), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n914), .A2(new_n921), .A3(new_n915), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n920), .B(new_n922), .C1(new_n917), .C2(new_n918), .ZN(G1350gat));
  NAND3_X1  g722(.A1(new_n831), .A2(new_n591), .A3(new_n900), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G190gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT61), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(KEYINPUT123), .A3(KEYINPUT61), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n925), .B2(KEYINPUT61), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n924), .A2(KEYINPUT124), .A3(new_n932), .A4(G190gat), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n928), .A2(new_n929), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n908), .A2(new_n223), .A3(new_n591), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1351gat));
  NOR2_X1   g735(.A1(new_n861), .A2(new_n478), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n903), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(G197gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n645), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT125), .Z(new_n941));
  AND2_X1   g740(.A1(new_n900), .A2(new_n487), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n886), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(G197gat), .B1(new_n943), .B2(new_n695), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n941), .A2(new_n944), .ZN(G1352gat));
  INV_X1    g744(.A(G204gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n938), .A2(new_n946), .A3(new_n621), .ZN(new_n947));
  OR3_X1    g746(.A1(new_n947), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT127), .B1(new_n947), .B2(KEYINPUT62), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(G204gat), .B1(new_n943), .B2(new_n740), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(KEYINPUT126), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n952), .A2(KEYINPUT126), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n950), .B(new_n951), .C1(new_n953), .C2(new_n954), .ZN(G1353gat));
  INV_X1    g754(.A(G211gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n938), .A2(new_n956), .A3(new_n691), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n886), .A2(new_n691), .A3(new_n942), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  OAI21_X1  g760(.A(G218gat), .B1(new_n943), .B2(new_n590), .ZN(new_n962));
  INV_X1    g761(.A(G218gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n938), .A2(new_n963), .A3(new_n591), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1355gat));
endmodule


