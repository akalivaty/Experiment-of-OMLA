//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1209;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT65), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n460), .B1(new_n465), .B2(G2105), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n458), .C1(new_n461), .C2(new_n462), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n470), .A2(KEYINPUT66), .A3(G137), .A4(new_n458), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n470), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n470), .A2(new_n458), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  AND2_X1   g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n461), .B2(new_n462), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT67), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT67), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(new_n488), .C1(new_n461), .C2(new_n462), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT69), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(new_n458), .C1(new_n462), .C2(new_n461), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n470), .A2(new_n499), .A3(new_n458), .A4(new_n496), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n493), .A2(new_n494), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n487), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n491), .B1(new_n470), .B2(new_n488), .ZN(new_n503));
  INV_X1    g078(.A(new_n492), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT68), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n515), .A2(new_n516), .B1(new_n509), .B2(new_n510), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n518), .A2(new_n524), .ZN(G166));
  NOR2_X1   g100(.A1(new_n509), .A2(new_n510), .ZN(new_n526));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n528), .A2(G51), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n521), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  INV_X1    g113(.A(new_n517), .ZN(new_n539));
  AOI22_X1  g114(.A1(G90), .A2(new_n539), .B1(new_n528), .B2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n516), .A2(new_n515), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n539), .A2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n528), .A2(G43), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n548), .B(new_n549), .C1(new_n523), .C2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT70), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n542), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(G651), .A2(new_n561), .B1(new_n539), .B2(G91), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n528), .B2(G53), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n562), .B1(new_n564), .B2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G52), .ZN(new_n568));
  INV_X1    g143(.A(G90), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n512), .A2(new_n568), .B1(new_n569), .B2(new_n517), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n544), .A2(G651), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT71), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT71), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n540), .A2(new_n573), .A3(new_n545), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G301));
  INV_X1    g151(.A(G166), .ZN(G303));
  OAI21_X1  g152(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  INV_X1    g154(.A(G49), .ZN(new_n580));
  OAI221_X1 g155(.A(new_n578), .B1(new_n579), .B2(new_n517), .C1(new_n512), .C2(new_n580), .ZN(G288));
  OAI211_X1 g156(.A(G48), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n517), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(G61), .B1(new_n516), .B2(new_n515), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n523), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT72), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT72), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(new_n584), .B2(new_n587), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n589), .A2(new_n591), .ZN(G305));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n512), .A2(new_n593), .B1(new_n594), .B2(new_n517), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n523), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT73), .B(KEYINPUT10), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n517), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n542), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT74), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n528), .A2(G54), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n517), .B2(new_n600), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n602), .A2(new_n608), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT75), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  MUX2_X1   g192(.A(G301), .B(new_n616), .S(new_n617), .Z(G284));
  MUX2_X1   g193(.A(G301), .B(new_n616), .S(new_n617), .Z(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(new_n616), .ZN(new_n624));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND3_X1  g201(.A1(new_n613), .A2(new_n625), .A3(new_n615), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n479), .A2(G135), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT77), .Z(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(G111), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G2105), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n476), .B2(G123), .ZN(new_n636));
  AND2_X1   g211(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n470), .A2(new_n459), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n643), .A2(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n638), .A2(G2096), .ZN(new_n646));
  NAND4_X1  g221(.A1(new_n639), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(G156));
  XOR2_X1   g222(.A(KEYINPUT15), .B(G2435), .Z(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT81), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT80), .B(KEYINPUT14), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1341), .B(G1348), .Z(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT79), .ZN(new_n661));
  XOR2_X1   g236(.A(G2451), .B(G2454), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2067), .B(G2678), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT82), .ZN(new_n669));
  NOR2_X1   g244(.A1(G2072), .A2(G2078), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n442), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2084), .B(G2090), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n671), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n671), .B(KEYINPUT17), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n672), .C1(new_n669), .C2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n672), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n669), .A2(new_n678), .A3(new_n676), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n674), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2096), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(KEYINPUT84), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  OR3_X1    g264(.A1(new_n683), .A2(new_n684), .A3(KEYINPUT84), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n683), .A2(new_n684), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n685), .A2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(new_n695), .B(new_n694), .S(new_n689), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1991), .B(G1996), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n700), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n699), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n702), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n703), .A2(new_n707), .ZN(G229));
  NOR2_X1   g283(.A1(G6), .A2(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n589), .A2(new_n591), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G16), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT32), .B(G1981), .Z(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(KEYINPUT88), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1971), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n716), .A2(G23), .ZN(new_n720));
  INV_X1    g295(.A(G288), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n716), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT33), .B(G1976), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR3_X1   g299(.A1(new_n715), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT87), .B(KEYINPUT34), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n714), .A2(KEYINPUT88), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G16), .A2(G24), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n598), .B(KEYINPUT86), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1986), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n476), .A2(G119), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n479), .A2(G131), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n458), .A2(G107), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n733), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  MUX2_X1   g312(.A(G25), .B(new_n737), .S(G29), .Z(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n738), .B(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n732), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n728), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n743), .B2(new_n744), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT94), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G29), .B2(G32), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n479), .A2(G141), .B1(G105), .B2(new_n459), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n476), .A2(G129), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT26), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G29), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  MUX2_X1   g334(.A(new_n752), .B(new_n751), .S(new_n759), .Z(new_n760));
  XOR2_X1   g335(.A(KEYINPUT27), .B(G1996), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G4), .A2(G16), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT90), .Z(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n616), .B2(new_n716), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT91), .B(G1348), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT97), .B(KEYINPUT23), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT98), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n716), .A2(G20), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n769), .B(new_n770), .Z(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n621), .B2(new_n716), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G1956), .Z(new_n773));
  NOR2_X1   g348(.A1(G5), .A2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT95), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G171), .B2(G16), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G1961), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT96), .Z(new_n778));
  NAND4_X1  g353(.A1(new_n762), .A2(new_n767), .A3(new_n773), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n758), .A2(G35), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G162), .B2(new_n758), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT29), .B(G2090), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(G11), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(G11), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(G28), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n758), .B1(new_n787), .B2(G28), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n785), .B(new_n786), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n637), .B2(G29), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n758), .A2(G33), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT25), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n470), .A2(G127), .ZN(new_n795));
  NAND2_X1  g370(.A1(G115), .A2(G2104), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n458), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n794), .B(new_n797), .C1(G139), .C2(new_n479), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n792), .B1(new_n798), .B2(new_n758), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n783), .B(new_n791), .C1(G2072), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n716), .A2(G21), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G168), .B2(new_n716), .ZN(new_n802));
  INV_X1    g377(.A(G1966), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n799), .A2(G2072), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n804), .B(new_n805), .C1(G1961), .C2(new_n776), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n800), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(G16), .A2(G19), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n552), .B2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT92), .B(G1341), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n758), .A2(G26), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT28), .ZN(new_n813));
  OR2_X1    g388(.A1(G104), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n815));
  INV_X1    g390(.A(G140), .ZN(new_n816));
  INV_X1    g391(.A(G128), .ZN(new_n817));
  OAI221_X1 g392(.A(new_n815), .B1(new_n478), .B2(new_n816), .C1(new_n817), .C2(new_n475), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(new_n758), .ZN(new_n820));
  INV_X1    g395(.A(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G34), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(KEYINPUT24), .ZN(new_n824));
  AOI21_X1  g399(.A(G29), .B1(new_n823), .B2(KEYINPUT24), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(KEYINPUT93), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(KEYINPUT93), .B2(new_n825), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n473), .B2(new_n758), .ZN(new_n828));
  INV_X1    g403(.A(G2084), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n811), .A2(new_n822), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n758), .A2(G27), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G164), .B2(new_n758), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G2078), .ZN(new_n835));
  NOR4_X1   g410(.A1(new_n779), .A2(new_n807), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n747), .A2(new_n750), .A3(new_n836), .ZN(G150));
  INV_X1    g412(.A(G150), .ZN(G311));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT101), .B(G93), .Z(new_n840));
  OAI22_X1  g415(.A1(new_n512), .A2(new_n839), .B1(new_n517), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n521), .A2(G67), .ZN(new_n842));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n523), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G860), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n624), .A2(G559), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n552), .A2(new_n845), .A3(KEYINPUT102), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n841), .B2(new_n844), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n842), .A2(new_n843), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G651), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n517), .A2(new_n840), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n528), .A2(G55), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT102), .A4(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n855), .A2(new_n860), .A3(new_n551), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n852), .A2(new_n862), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n852), .A2(new_n862), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n866), .B1(new_n869), .B2(new_n863), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n849), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n846), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n868), .A2(new_n870), .A3(new_n849), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n848), .B1(new_n872), .B2(new_n873), .ZN(G145));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n875));
  OR2_X1    g450(.A1(G106), .A2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(G2104), .C1(G118), .C2(new_n458), .ZN(new_n877));
  INV_X1    g452(.A(G130), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n475), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(G142), .B2(new_n479), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n641), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n737), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n498), .A2(new_n500), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n493), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n818), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n757), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n798), .B(KEYINPUT103), .Z(new_n889));
  OR2_X1    g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n798), .A2(KEYINPUT103), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n884), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n882), .A2(new_n883), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(G160), .B(new_n483), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n637), .B(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n884), .A2(new_n890), .A3(new_n894), .A4(new_n892), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n898), .B1(new_n896), .B2(new_n899), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n875), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n905), .A2(KEYINPUT40), .A3(new_n901), .A4(new_n900), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n904), .A2(new_n906), .ZN(G395));
  XOR2_X1   g482(.A(new_n627), .B(new_n862), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n605), .B(KEYINPUT74), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n603), .B2(new_n542), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n910), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n602), .A2(new_n610), .ZN(new_n912));
  NAND3_X1  g487(.A1(G299), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n565), .B(KEYINPUT9), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n611), .A2(new_n914), .A3(KEYINPUT105), .A4(new_n562), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT105), .B1(new_n621), .B2(new_n611), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT106), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n612), .B2(G299), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n920), .A2(new_n921), .A3(new_n913), .A4(new_n915), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n908), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n913), .A2(new_n915), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(KEYINPUT41), .A3(new_n920), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n916), .B2(new_n917), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n908), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n925), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  NAND2_X1  g509(.A1(G305), .A2(G290), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n598), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n721), .B(G166), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n935), .A3(new_n936), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(KEYINPUT107), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT108), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n925), .A2(new_n945), .A3(new_n932), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n934), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n944), .B1(new_n934), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(G868), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n617), .B1(new_n841), .B2(new_n844), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(G295));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n950), .ZN(G331));
  NAND2_X1  g527(.A1(new_n940), .A2(new_n941), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n927), .A2(new_n929), .A3(KEYINPUT109), .ZN(new_n954));
  AOI21_X1  g529(.A(G286), .B1(new_n572), .B2(new_n574), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n540), .A2(new_n545), .B1(new_n532), .B2(new_n536), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n853), .B(new_n861), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n575), .B2(G168), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n862), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n957), .B(new_n959), .C1(new_n927), .C2(KEYINPUT109), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n918), .A2(new_n922), .B1(new_n959), .B2(new_n957), .ZN(new_n961));
  OAI22_X1  g536(.A1(new_n954), .A2(new_n960), .B1(new_n961), .B2(KEYINPUT110), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n957), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n923), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n953), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n963), .B1(new_n929), .B2(new_n927), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n959), .A2(new_n957), .B1(new_n920), .B2(new_n926), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n970), .B2(new_n942), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n953), .B1(new_n968), .B2(new_n969), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n963), .B1(new_n917), .B2(new_n916), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n976), .B(new_n942), .C1(new_n930), .C2(new_n963), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n901), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT43), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n973), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n927), .A2(new_n929), .A3(KEYINPUT109), .ZN(new_n983));
  NOR4_X1   g558(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT109), .A4(new_n928), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(new_n963), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n983), .A2(new_n985), .B1(new_n964), .B2(new_n965), .ZN(new_n986));
  INV_X1    g561(.A(new_n966), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n942), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT43), .B1(new_n988), .B2(new_n978), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n974), .A2(new_n977), .A3(new_n972), .A4(new_n901), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT44), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT111), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n972), .B1(new_n967), .B2(new_n971), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n994), .A2(new_n991), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n982), .B1(new_n993), .B2(new_n996), .ZN(G397));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n886), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n466), .A2(G40), .A3(new_n472), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1986), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n598), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(G1986), .A3(G290), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n1007), .B(KEYINPUT113), .Z(new_n1008));
  XNOR2_X1  g583(.A(new_n818), .B(G2067), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT114), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n757), .B(G1996), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1011), .B1(new_n1003), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n737), .A2(new_n740), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n737), .A2(new_n740), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1003), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1008), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT115), .ZN(new_n1018));
  INV_X1    g593(.A(G2078), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1384), .B1(new_n493), .B2(new_n885), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1002), .B1(new_n1020), .B2(KEYINPUT45), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n501), .B2(new_n506), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1000), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1019), .B(new_n1021), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1002), .B1(new_n1020), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1029));
  INV_X1    g604(.A(G1961), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT125), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT53), .B1(new_n1032), .B2(G2078), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n1032), .B2(G2078), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1021), .A2(new_n1001), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1026), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT126), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1026), .A2(new_n1031), .A3(KEYINPUT126), .A4(new_n1035), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(G171), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT127), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT127), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1038), .A2(new_n1042), .A3(G171), .A4(new_n1039), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1002), .B1(new_n999), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n885), .B1(new_n505), .B2(KEYINPUT68), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n493), .A2(new_n494), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n998), .B(new_n1023), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n1048), .A3(new_n1019), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT124), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1045), .A2(new_n1048), .A3(KEYINPUT124), .A4(new_n1019), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(KEYINPUT53), .A3(new_n1052), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1024), .A2(new_n1025), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(G301), .A3(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1055), .A2(KEYINPUT54), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1041), .A2(new_n1043), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n1058));
  AOI21_X1  g633(.A(G301), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1036), .A2(new_n575), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT121), .B(G1956), .ZN(new_n1062));
  AOI211_X1 g637(.A(KEYINPUT50), .B(G1384), .C1(new_n501), .C2(new_n506), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n466), .A2(G40), .A3(new_n472), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n1020), .B2(new_n1027), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1062), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(G299), .B(KEYINPUT57), .Z(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1021), .B(new_n1068), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1348), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1064), .A2(new_n1020), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1029), .A2(new_n1071), .B1(new_n821), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(new_n611), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1067), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1070), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT61), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(new_n1076), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1067), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(KEYINPUT61), .A3(new_n1070), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(G1341), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1072), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(G1996), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n552), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1029), .A2(new_n1071), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1073), .A2(new_n821), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n611), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n611), .A2(new_n1096), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT123), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1090), .A2(KEYINPUT59), .A3(new_n552), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1074), .A2(new_n1100), .A3(new_n1097), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1093), .A2(new_n1102), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1077), .B1(new_n1085), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G8), .ZN(new_n1107));
  NOR2_X1   g682(.A1(G166), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(G166), .B2(new_n1107), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1065), .B1(new_n1027), .B2(new_n1022), .ZN(new_n1115));
  INV_X1    g690(.A(G2090), .ZN(new_n1116));
  INV_X1    g691(.A(G1971), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1115), .A2(new_n1116), .B1(new_n1089), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1114), .B1(new_n1118), .B2(new_n1107), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1089), .A2(new_n1117), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1116), .B(new_n1028), .C1(new_n1022), .C2(new_n1027), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1107), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1113), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1107), .B1(new_n1064), .B2(new_n1020), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n721), .A2(G1976), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT52), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT117), .B(G1976), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT52), .B1(G288), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1124), .A2(new_n1125), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n1132));
  OAI21_X1  g707(.A(G1981), .B1(new_n584), .B2(new_n587), .ZN(new_n1133));
  INV_X1    g708(.A(G61), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n519), .B2(new_n520), .ZN(new_n1135));
  INV_X1    g710(.A(new_n586), .ZN(new_n1136));
  OAI21_X1  g711(.A(G651), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n511), .A2(G86), .A3(new_n521), .ZN(new_n1138));
  INV_X1    g713(.A(G1981), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .A4(new_n582), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1133), .A2(new_n1140), .A3(KEYINPUT49), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1141), .B(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1133), .A2(new_n1140), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT49), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1124), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1132), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1141), .B(KEYINPUT118), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1149), .A2(KEYINPUT119), .A3(new_n1124), .A4(new_n1146), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1131), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1119), .A2(new_n1123), .A3(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT120), .B(G2084), .Z(new_n1153));
  OAI211_X1 g728(.A(new_n1028), .B(new_n1153), .C1(new_n1022), .C2(new_n1027), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1064), .B1(new_n1020), .B2(KEYINPUT45), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(new_n1023), .B2(new_n1022), .ZN(new_n1156));
  OAI211_X1 g731(.A(G168), .B(new_n1154), .C1(new_n1156), .C2(G1966), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(G8), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n803), .ZN(new_n1160));
  AOI21_X1  g735(.A(G168), .B1(new_n1160), .B2(new_n1154), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT51), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT51), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1157), .A2(new_n1163), .A3(G8), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1152), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  AND4_X1   g740(.A1(new_n1057), .A2(new_n1061), .A3(new_n1106), .A4(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT62), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1162), .A2(new_n1169), .A3(new_n1164), .ZN(new_n1170));
  AND4_X1   g745(.A1(new_n1059), .A2(new_n1119), .A3(new_n1123), .A4(new_n1151), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1131), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1173), .A2(new_n1122), .A3(new_n1174), .A4(new_n1113), .ZN(new_n1175));
  NOR2_X1   g750(.A1(G288), .A2(G1976), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1173), .A2(new_n1176), .B1(new_n1139), .B2(new_n588), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1124), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1175), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(G168), .A2(G8), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1180), .B1(new_n1160), .B2(new_n1154), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1119), .A2(new_n1123), .A3(new_n1151), .A4(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1122), .A2(new_n1113), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1181), .A2(KEYINPUT63), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1185), .A2(new_n1186), .A3(new_n1123), .A4(new_n1151), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1179), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1172), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1018), .B1(new_n1166), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1003), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n819), .A2(new_n821), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1195));
  XOR2_X1   g770(.A(new_n1005), .B(KEYINPUT48), .Z(new_n1196));
  NOR2_X1   g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OR3_X1    g772(.A1(new_n1191), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1198));
  OAI21_X1  g773(.A(KEYINPUT46), .B1(new_n1191), .B2(G1996), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1009), .A2(new_n757), .ZN(new_n1200));
  AOI22_X1  g775(.A1(new_n1198), .A2(new_n1199), .B1(new_n1200), .B2(new_n1003), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT47), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n1194), .A2(new_n1197), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1190), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g779(.A(G319), .ZN(new_n1206));
  NOR2_X1   g780(.A1(G227), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n1207), .A2(new_n666), .ZN(new_n1208));
  AOI21_X1  g782(.A(new_n1208), .B1(new_n703), .B2(new_n707), .ZN(new_n1209));
  OAI211_X1 g783(.A(new_n980), .B(new_n1209), .C1(new_n903), .C2(new_n902), .ZN(G225));
  INV_X1    g784(.A(G225), .ZN(G308));
endmodule


