//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G141gat), .B(G148gat), .Z(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT2), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G155gat), .B(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n208), .A2(new_n213), .A3(new_n211), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT70), .ZN(new_n221));
  INV_X1    g020(.A(G113gat), .ZN(new_n222));
  INV_X1    g021(.A(G120gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT1), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G113gat), .A2(G120gat), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n220), .A2(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(G127gat), .B(G134gat), .Z(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT70), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n226), .B(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(new_n215), .B2(new_n216), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n219), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n215), .A2(new_n216), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n233), .A3(KEYINPUT4), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT5), .ZN(new_n237));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT4), .B1(new_n229), .B2(new_n233), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n236), .A2(new_n237), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n242));
  INV_X1    g041(.A(new_n229), .ZN(new_n243));
  INV_X1    g042(.A(new_n231), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n243), .B(new_n244), .C1(new_n217), .C2(new_n218), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n245), .A2(new_n240), .A3(new_n238), .A4(new_n234), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n229), .B(new_n233), .ZN(new_n247));
  INV_X1    g046(.A(new_n238), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n237), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n241), .A2(new_n242), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n246), .A3(new_n242), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n207), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT6), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n242), .B1(new_n246), .B2(KEYINPUT5), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n249), .A2(new_n246), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(new_n206), .A3(new_n251), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(KEYINPUT6), .B(new_n207), .C1(new_n250), .C2(new_n252), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT73), .ZN(new_n261));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT22), .ZN(new_n263));
  INV_X1    g062(.A(G211gat), .ZN(new_n264));
  INV_X1    g063(.A(G218gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n262), .A3(new_n266), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n272), .A2(new_n273), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n261), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n270), .A2(new_n271), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT72), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(new_n274), .A3(KEYINPUT73), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT74), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT23), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n288), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT25), .B1(new_n291), .B2(KEYINPUT66), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n289), .A2(new_n290), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n295));
  OR2_X1    g094(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(G190gat), .A3(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n293), .A2(new_n287), .A3(new_n295), .A4(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n292), .A2(new_n299), .ZN(new_n301));
  INV_X1    g100(.A(G183gat), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT27), .B1(new_n302), .B2(KEYINPUT67), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT27), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G183gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n303), .B(new_n294), .C1(KEYINPUT67), .C2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n302), .A2(KEYINPUT27), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n309), .A2(new_n305), .A3(KEYINPUT28), .A4(new_n294), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT69), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n308), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G169gat), .ZN(new_n315));
  INV_X1    g114(.A(G176gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT26), .ZN(new_n318));
  OAI22_X1  g117(.A1(new_n317), .A2(new_n318), .B1(new_n302), .B2(new_n294), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT26), .B1(new_n315), .B2(new_n316), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(new_n290), .B2(new_n320), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n300), .A2(new_n301), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n285), .B1(new_n322), .B2(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT75), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n300), .A2(new_n301), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n314), .A2(new_n321), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n284), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT75), .B1(new_n323), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n282), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n284), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n322), .A2(new_n285), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n275), .A2(new_n276), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G64gat), .B(G92gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  NAND3_X1  g139(.A1(new_n331), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n259), .A2(new_n260), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT82), .ZN(new_n343));
  INV_X1    g142(.A(new_n340), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n333), .B2(new_n334), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n281), .B1(new_n346), .B2(new_n324), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(new_n336), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT37), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n343), .B(new_n344), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n349), .B1(new_n331), .B2(new_n337), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT82), .B1(new_n351), .B2(new_n340), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT38), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n348), .B2(new_n349), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n331), .A2(new_n337), .A3(new_n349), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n344), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n346), .A2(new_n324), .A3(new_n281), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n335), .B1(new_n333), .B2(new_n334), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n349), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n353), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n342), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n332), .B1(new_n217), .B2(new_n218), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT29), .B1(new_n270), .B2(new_n271), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n217), .B1(new_n365), .B2(new_n218), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n335), .A2(new_n363), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n366), .A2(new_n364), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G22gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n277), .A2(new_n280), .A3(new_n363), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n230), .B1(new_n278), .B2(KEYINPUT29), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n370), .B1(new_n374), .B2(new_n217), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n367), .A2(new_n368), .B1(G228gat), .B2(G233gat), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n373), .A2(new_n375), .ZN(new_n379));
  OAI21_X1  g178(.A(G22gat), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT31), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(G50gat), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n381), .A2(KEYINPUT80), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n377), .A2(new_n380), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n384), .B1(new_n381), .B2(KEYINPUT80), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n344), .B1(new_n347), .B2(new_n336), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(KEYINPUT30), .A3(new_n341), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT30), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n348), .A2(new_n392), .A3(new_n340), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n236), .A2(new_n240), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n248), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n397), .B(KEYINPUT39), .C1(new_n247), .C2(new_n248), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT39), .B1(new_n247), .B2(new_n248), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT81), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n238), .B1(new_n236), .B2(new_n240), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT39), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n207), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n401), .A2(new_n404), .A3(KEYINPUT40), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT40), .B1(new_n401), .B2(new_n404), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n253), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n389), .B1(new_n394), .B2(new_n408), .ZN(new_n409));
  OR2_X1    g208(.A1(new_n362), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n411), .B(KEYINPUT64), .Z(new_n412));
  NAND2_X1  g211(.A1(new_n328), .A2(new_n229), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n322), .A2(new_n243), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT34), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n413), .A2(new_n414), .A3(new_n412), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419));
  XOR2_X1   g218(.A(G15gat), .B(G43gat), .Z(new_n420));
  XNOR2_X1  g219(.A(G71gat), .B(G99gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n418), .B(KEYINPUT32), .C1(new_n419), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n418), .A2(KEYINPUT32), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n418), .A2(new_n419), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n422), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n417), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT71), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n417), .A2(KEYINPUT71), .B1(new_n427), .B2(new_n424), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT36), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n417), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n427), .A2(new_n424), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n428), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n432), .B1(new_n436), .B2(KEYINPUT36), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n259), .A2(new_n260), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n394), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n388), .A2(new_n387), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n381), .A2(KEYINPUT80), .A3(new_n384), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n440), .B(new_n441), .C1(new_n430), .C2(new_n431), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT35), .B1(new_n445), .B2(new_n439), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT35), .B1(new_n259), .B2(new_n260), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n389), .A2(new_n447), .A3(new_n394), .A4(new_n436), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n410), .A2(new_n444), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT15), .ZN(new_n450));
  INV_X1    g249(.A(G43gat), .ZN(new_n451));
  INV_X1    g250(.A(G50gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G43gat), .A2(G50gat), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AND2_X1   g254(.A1(G43gat), .A2(G50gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n450), .A2(KEYINPUT83), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT15), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n456), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n451), .A2(KEYINPUT84), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(G43gat), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n463), .A3(new_n452), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(G29gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n467));
  INV_X1    g266(.A(G36gat), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n466), .B2(KEYINPUT14), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT14), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(G29gat), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n467), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n455), .B1(new_n465), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n455), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT85), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n466), .A2(KEYINPUT14), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n470), .A2(G29gat), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n468), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n464), .A2(new_n460), .B1(new_n480), .B2(new_n467), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n477), .B(new_n474), .C1(new_n481), .C2(new_n455), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n483));
  NAND3_X1  g282(.A1(new_n476), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n372), .A2(G15gat), .ZN(new_n485));
  INV_X1    g284(.A(G15gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G22gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G1gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(KEYINPUT16), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(new_n491), .B2(G1gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(G8gat), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G8gat), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n490), .B(new_n493), .C1(new_n495), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT17), .B1(new_n473), .B2(new_n475), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n484), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n476), .A2(new_n500), .A3(new_n482), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n503), .A2(KEYINPUT18), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n476), .A2(new_n482), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n501), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n505), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n504), .B(KEYINPUT13), .Z(new_n511));
  AOI21_X1  g310(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n476), .A2(new_n500), .A3(new_n482), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n500), .B1(new_n476), .B2(new_n482), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n507), .B(new_n511), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n506), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G113gat), .B(G141gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G197gat), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT11), .B(G169gat), .Z(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT12), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n520), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT91), .B1(new_n517), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT90), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n515), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n526), .B1(new_n518), .B2(new_n519), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n506), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n518), .A2(KEYINPUT89), .A3(new_n519), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n538), .A2(new_n506), .A3(new_n532), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n526), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(KEYINPUT41), .ZN(new_n545));
  XNOR2_X1  g344(.A(G134gat), .B(G162gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT97), .ZN(new_n549));
  INV_X1    g348(.A(G92gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT95), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT95), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G92gat), .ZN(new_n553));
  INV_X1    g352(.A(G85gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT7), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT7), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(G85gat), .A3(G92gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G99gat), .A2(G106gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT8), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G99gat), .B(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n555), .A2(new_n560), .A3(new_n564), .A4(new_n562), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n566), .A2(KEYINPUT96), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT96), .B1(new_n566), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n549), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT95), .B(G92gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n572), .A2(new_n554), .B1(KEYINPUT8), .B2(new_n561), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n564), .B1(new_n573), .B2(new_n560), .ZN(new_n574));
  INV_X1    g373(.A(new_n567), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n571), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n566), .A2(KEYINPUT96), .A3(new_n567), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(KEYINPUT97), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n570), .A2(new_n578), .A3(new_n484), .A4(new_n502), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT98), .ZN(new_n580));
  XOR2_X1   g379(.A(G190gat), .B(G218gat), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n508), .A2(new_n568), .A3(new_n569), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n583), .B1(KEYINPUT41), .B2(new_n544), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n582), .B1(new_n580), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n548), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n580), .A2(new_n584), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n581), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(new_n547), .A3(new_n585), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G57gat), .B(G64gat), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G57gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G64gat), .ZN(new_n600));
  INV_X1    g399(.A(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G57gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G71gat), .B(G78gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n597), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n608));
  AND2_X1   g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT20), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n610), .B(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n500), .B1(KEYINPUT21), .B2(new_n607), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n613), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n617), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n592), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n598), .A2(new_n606), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n576), .A2(new_n577), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n607), .B1(new_n574), .B2(new_n575), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n566), .A2(new_n624), .A3(new_n567), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT10), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n623), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n623), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n628), .A2(new_n632), .A3(new_n629), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n636), .B1(new_n631), .B2(new_n633), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OR4_X1    g440(.A1(new_n449), .A2(new_n543), .A3(new_n622), .A4(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n438), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n489), .ZN(G1324gat));
  OAI21_X1  g443(.A(G8gat), .B1(new_n642), .B2(new_n394), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n645), .A2(KEYINPUT42), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n642), .A2(new_n394), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT16), .B(G8gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n651));
  MUX2_X1   g450(.A(KEYINPUT100), .B(new_n651), .S(new_n649), .Z(new_n652));
  AOI22_X1  g451(.A1(new_n646), .A2(new_n650), .B1(new_n647), .B2(new_n652), .ZN(G1325gat));
  XNOR2_X1  g452(.A(new_n437), .B(KEYINPUT101), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(G15gat), .B1(new_n642), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n436), .A2(new_n486), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n642), .B2(new_n657), .ZN(G1326gat));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n389), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT43), .B(G22gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n543), .A2(new_n621), .A3(new_n641), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n449), .A2(new_n592), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n438), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n466), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT45), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n446), .A2(new_n448), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n391), .A2(new_n393), .B1(new_n259), .B2(new_n260), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n672), .B2(new_n389), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n439), .A2(KEYINPUT102), .A3(new_n442), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n674), .A3(new_n437), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n362), .A2(new_n409), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n670), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n670), .B(KEYINPUT103), .C1(new_n675), .C2(new_n676), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n592), .A2(KEYINPUT44), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT44), .B1(new_n449), .B2(new_n592), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n664), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n466), .B1(new_n684), .B2(new_n666), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n662), .B1(new_n669), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n685), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n667), .B(KEYINPUT45), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n688), .A3(KEYINPUT104), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(G1328gat));
  INV_X1    g489(.A(new_n394), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n665), .A2(new_n468), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT46), .Z(new_n693));
  INV_X1    g492(.A(new_n684), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT105), .B1(new_n694), .B2(new_n394), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G36gat), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n694), .A2(KEYINPUT105), .A3(new_n394), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n693), .B1(new_n696), .B2(new_n697), .ZN(G1329gat));
  NAND2_X1  g497(.A1(new_n461), .A2(new_n463), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n694), .B2(new_n437), .ZN(new_n700));
  INV_X1    g499(.A(new_n436), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n699), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n665), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n700), .A2(KEYINPUT47), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n684), .A2(new_n654), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n705), .A2(new_n699), .B1(new_n665), .B2(new_n702), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n706), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g506(.A1(new_n684), .A2(new_n442), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G50gat), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT48), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n665), .A2(new_n452), .A3(new_n442), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n710), .B1(new_n709), .B2(new_n711), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(G1331gat));
  AND2_X1   g513(.A1(new_n679), .A2(new_n680), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n622), .A2(new_n542), .A3(new_n640), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n438), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT106), .B(G57gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1332gat));
  AND2_X1   g519(.A1(new_n715), .A2(new_n716), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n394), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n723), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT107), .B1(new_n717), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n724), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1333gat));
  OR3_X1    g530(.A1(new_n717), .A2(G71gat), .A3(new_n701), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n733));
  OAI21_X1  g532(.A(G71gat), .B1(new_n717), .B2(new_n655), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(G1334gat));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n442), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G78gat), .ZN(G1335gat));
  INV_X1    g538(.A(new_n621), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(new_n543), .A3(new_n641), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT108), .Z(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(new_n682), .B2(new_n683), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n744), .A2(new_n554), .A3(new_n438), .ZN(new_n745));
  AND2_X1   g544(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n746));
  INV_X1    g545(.A(new_n592), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n677), .A2(KEYINPUT109), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n621), .A2(new_n542), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT109), .B1(new_n677), .B2(new_n747), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n746), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n677), .A2(new_n747), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n746), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n755), .A2(new_n748), .A3(new_n749), .A4(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n752), .A2(new_n641), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n666), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n745), .B1(new_n761), .B2(new_n554), .ZN(G1336gat));
  NAND2_X1  g561(.A1(new_n691), .A2(new_n550), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n572), .B1(new_n743), .B2(new_n691), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n765), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n767), .B(new_n768), .C1(new_n759), .C2(new_n763), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(G1337gat));
  INV_X1    g569(.A(G99gat), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n744), .A2(new_n771), .A3(new_n655), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n760), .A2(new_n436), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(new_n771), .ZN(G1338gat));
  NOR2_X1   g573(.A1(new_n389), .A2(G106gat), .ZN(new_n775));
  AND4_X1   g574(.A1(new_n641), .A2(new_n752), .A3(new_n758), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(KEYINPUT111), .B(G106gat), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n743), .B2(new_n442), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT53), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n743), .A2(KEYINPUT112), .A3(new_n442), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT112), .B1(new_n743), .B2(new_n442), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n780), .A2(new_n781), .A3(new_n777), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  INV_X1    g582(.A(new_n775), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n759), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n779), .B1(new_n782), .B2(new_n785), .ZN(G1339gat));
  NOR3_X1   g585(.A1(new_n622), .A2(new_n542), .A3(new_n641), .ZN(new_n787));
  INV_X1    g586(.A(new_n524), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n503), .A2(new_n505), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(G229gat), .A3(G233gat), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n510), .A2(new_n511), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n518), .ZN(new_n794));
  AOI22_X1  g593(.A1(KEYINPUT18), .A2(new_n794), .B1(new_n531), .B2(new_n515), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n534), .B1(new_n795), .B2(new_n533), .ZN(new_n796));
  INV_X1    g595(.A(new_n535), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n641), .B(new_n793), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT114), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n566), .A2(new_n624), .A3(new_n567), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n624), .B1(new_n566), .B2(new_n567), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n625), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n576), .A2(new_n577), .A3(new_n626), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n803), .A3(new_n632), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n631), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n632), .B1(new_n802), .B2(new_n803), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n636), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n808), .A3(KEYINPUT55), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n809), .A2(KEYINPUT113), .A3(new_n637), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT113), .B1(new_n809), .B2(new_n637), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT55), .B1(new_n805), .B2(new_n808), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n542), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n792), .B1(new_n529), .B2(new_n535), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n816), .A3(new_n641), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n799), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n592), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n813), .A2(new_n588), .A3(new_n815), .A4(new_n591), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n787), .B1(new_n821), .B2(new_n740), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n438), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n691), .A2(new_n442), .A3(new_n701), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n222), .B1(new_n825), .B2(new_n542), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT115), .Z(new_n827));
  NOR3_X1   g626(.A1(new_n822), .A2(new_n438), .A3(new_n445), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n394), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n542), .A2(new_n222), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(G1340gat));
  NAND2_X1  g630(.A1(new_n825), .A2(new_n641), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G120gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n641), .A2(new_n223), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT116), .ZN(G1341gat));
  INV_X1    g635(.A(new_n825), .ZN(new_n837));
  OAI21_X1  g636(.A(G127gat), .B1(new_n837), .B2(new_n740), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n740), .A2(G127gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n829), .B2(new_n839), .ZN(G1342gat));
  INV_X1    g639(.A(G134gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n747), .A2(new_n394), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT117), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT56), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT118), .ZN(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n837), .B2(new_n592), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n847), .B(new_n848), .C1(KEYINPUT56), .C2(new_n845), .ZN(G1343gat));
  NAND3_X1  g648(.A1(new_n437), .A2(new_n666), .A3(new_n394), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n852), .B(new_n853), .C1(new_n822), .C2(new_n389), .ZN(new_n854));
  INV_X1    g653(.A(new_n812), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n637), .A3(new_n809), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n536), .B2(new_n541), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n640), .B(new_n792), .C1(new_n529), .C2(new_n535), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n592), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n621), .B1(new_n859), .B2(new_n820), .ZN(new_n860));
  OAI211_X1 g659(.A(KEYINPUT57), .B(new_n442), .C1(new_n860), .C2(new_n787), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n787), .ZN(new_n863));
  INV_X1    g662(.A(new_n820), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(new_n818), .B2(new_n592), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n863), .B1(new_n865), .B2(new_n621), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n866), .B2(new_n442), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(new_n852), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n851), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G141gat), .B1(new_n869), .B2(new_n543), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n823), .A2(new_n442), .A3(new_n655), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n691), .ZN(new_n872));
  INV_X1    g671(.A(G141gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n542), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT58), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n870), .A2(new_n877), .A3(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1344gat));
  OAI211_X1 g678(.A(new_n641), .B(new_n851), .C1(new_n862), .C2(new_n868), .ZN(new_n880));
  INV_X1    g679(.A(G148gat), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(KEYINPUT59), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n866), .A2(KEYINPUT57), .A3(new_n442), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n442), .B1(new_n860), .B2(new_n787), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT120), .B1(new_n884), .B2(new_n853), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n866), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n442), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n886), .A2(new_n641), .A3(new_n851), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G148gat), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n880), .A2(new_n882), .B1(new_n889), .B2(KEYINPUT59), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n881), .A3(new_n641), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT121), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n894));
  INV_X1    g693(.A(new_n882), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n867), .A2(new_n852), .ZN(new_n896));
  INV_X1    g695(.A(new_n861), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n867), .B2(new_n852), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n850), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n895), .B1(new_n899), .B2(new_n641), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n888), .B2(G148gat), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n891), .B(new_n894), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n893), .A2(new_n903), .ZN(G1345gat));
  OAI21_X1  g703(.A(G155gat), .B1(new_n869), .B2(new_n740), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n872), .A2(new_n209), .A3(new_n621), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1346gat));
  OAI21_X1  g706(.A(G162gat), .B1(new_n869), .B2(new_n592), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n844), .A2(new_n210), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n871), .B2(new_n909), .ZN(G1347gat));
  NAND2_X1  g709(.A1(new_n691), .A2(new_n438), .ZN(new_n911));
  OR3_X1    g710(.A1(new_n911), .A2(KEYINPUT124), .A3(new_n701), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT124), .B1(new_n911), .B2(new_n701), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n389), .A3(new_n866), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(new_n315), .A3(new_n543), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n822), .A2(new_n666), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n445), .A2(new_n394), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n918), .B(KEYINPUT122), .Z(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT123), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n542), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n916), .B1(new_n924), .B2(new_n315), .ZN(G1348gat));
  OAI21_X1  g724(.A(G176gat), .B1(new_n915), .B2(new_n640), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n921), .A2(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n641), .A2(new_n316), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(G1349gat));
  OAI21_X1  g728(.A(G183gat), .B1(new_n915), .B2(new_n740), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n621), .A2(new_n309), .A3(new_n305), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n920), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g732(.A(G190gat), .B1(new_n915), .B2(new_n592), .ZN(new_n934));
  XOR2_X1   g733(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n936), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n747), .A2(new_n294), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n937), .B(new_n938), .C1(new_n927), .C2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT126), .ZN(G1351gat));
  NOR3_X1   g740(.A1(new_n654), .A2(new_n394), .A3(new_n389), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n917), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(G197gat), .B1(new_n943), .B2(new_n542), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n886), .A2(new_n887), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n654), .A2(new_n911), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n542), .A2(G197gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G1352gat));
  INV_X1    g748(.A(G204gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n943), .A2(new_n950), .A3(new_n641), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT62), .Z(new_n952));
  AND3_X1   g751(.A1(new_n945), .A2(new_n641), .A3(new_n946), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n950), .B2(new_n953), .ZN(G1353gat));
  NAND3_X1  g753(.A1(new_n943), .A2(new_n264), .A3(new_n621), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n945), .A2(new_n621), .A3(new_n946), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n265), .A3(new_n747), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n947), .A2(new_n747), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(new_n265), .ZN(G1355gat));
endmodule


