//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(G125), .A2(G140), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT72), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT72), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n190), .B1(new_n195), .B2(G140), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT73), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT73), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(new_n192), .B2(new_n194), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n199), .B(KEYINPUT16), .C1(new_n201), .C2(new_n190), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT72), .B(G125), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n204), .A2(KEYINPUT16), .A3(G140), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(G146), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G125), .B(G140), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT19), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n190), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n204), .B2(new_n200), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n210), .B1(new_n212), .B2(new_n209), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT93), .ZN(new_n214));
  OR3_X1    g028(.A1(new_n213), .A2(new_n214), .A3(G146), .ZN(new_n215));
  INV_X1    g029(.A(G237), .ZN(new_n216));
  INV_X1    g030(.A(G953), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G143), .A4(G214), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n216), .A2(new_n217), .A3(G214), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n218), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT92), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT92), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n228), .A3(G131), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n230), .B(new_n218), .C1(new_n223), .C2(new_n224), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT91), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT64), .B(G143), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n216), .A2(new_n217), .A3(G214), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT91), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n235), .A2(new_n236), .A3(new_n230), .A4(new_n218), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n227), .A2(new_n229), .A3(new_n232), .A4(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n214), .B1(new_n213), .B2(G146), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n207), .A2(new_n215), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT90), .ZN(new_n241));
  INV_X1    g055(.A(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n208), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n241), .B(new_n243), .C1(new_n212), .C2(new_n242), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n196), .A2(KEYINPUT90), .A3(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT18), .A2(G131), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n235), .A2(new_n246), .A3(new_n218), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n225), .A2(KEYINPUT18), .A3(G131), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n244), .A2(new_n245), .A3(new_n247), .A4(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n189), .B1(new_n240), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT94), .ZN(new_n252));
  INV_X1    g066(.A(new_n249), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT17), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n227), .B2(new_n229), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n232), .A2(new_n237), .ZN(new_n256));
  AOI211_X1 g070(.A(KEYINPUT92), .B(new_n230), .C1(new_n235), .C2(new_n218), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n228), .B1(new_n225), .B2(G131), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n255), .B1(new_n259), .B2(new_n254), .ZN(new_n260));
  AOI21_X1  g074(.A(G146), .B1(new_n203), .B2(new_n206), .ZN(new_n261));
  AOI211_X1 g075(.A(new_n242), .B(new_n205), .C1(new_n198), .C2(new_n202), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n253), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n252), .B1(new_n264), .B2(new_n189), .ZN(new_n265));
  INV_X1    g079(.A(new_n202), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n199), .B1(new_n212), .B2(KEYINPUT16), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n206), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n242), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n207), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT17), .B1(new_n257), .B2(new_n258), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n238), .B2(KEYINPUT17), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n189), .B(new_n249), .C1(new_n270), .C2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(KEYINPUT94), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n251), .B1(new_n265), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT20), .ZN(new_n276));
  NOR2_X1   g090(.A1(G475), .A2(G902), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(KEYINPUT94), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n260), .A2(new_n263), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n280), .A2(new_n252), .A3(new_n189), .A4(new_n249), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n250), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n277), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT20), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n265), .A2(new_n274), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n264), .A2(new_n189), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n278), .A2(new_n284), .B1(new_n288), .B2(G475), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n217), .A2(G952), .ZN(new_n290));
  NAND2_X1  g104(.A1(G234), .A2(G237), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(G902), .A3(G953), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT21), .B(G898), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G478), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(KEYINPUT15), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT96), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT13), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n233), .A2(new_n303), .A3(G128), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n233), .A2(G128), .ZN(new_n305));
  INV_X1    g119(.A(G128), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G143), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(G134), .B(new_n304), .C1(new_n308), .C2(new_n303), .ZN(new_n309));
  INV_X1    g123(.A(G134), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n305), .A2(new_n310), .A3(new_n307), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT76), .B(G107), .ZN(new_n312));
  XNOR2_X1  g126(.A(G116), .B(G122), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n309), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT95), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT95), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n309), .A2(new_n317), .A3(new_n311), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n308), .A2(G134), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n311), .ZN(new_n320));
  INV_X1    g134(.A(G107), .ZN(new_n321));
  INV_X1    g135(.A(G116), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n322), .A2(G122), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n321), .B1(new_n323), .B2(KEYINPUT14), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT14), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n313), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n324), .A2(new_n326), .B1(new_n312), .B2(new_n313), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n320), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n316), .A2(new_n318), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT9), .B(G234), .ZN(new_n330));
  INV_X1    g144(.A(G217), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n330), .A2(new_n331), .A3(G953), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n316), .A2(new_n318), .A3(new_n328), .A4(new_n332), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n302), .B1(new_n336), .B2(new_n285), .ZN(new_n337));
  AOI211_X1 g151(.A(KEYINPUT96), .B(G902), .C1(new_n334), .C2(new_n335), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n301), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n285), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n300), .B1(new_n340), .B2(KEYINPUT96), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n289), .A2(new_n298), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(G210), .B1(G237), .B2(G902), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OR2_X1    g161(.A1(KEYINPUT0), .A2(G128), .ZN(new_n348));
  NAND2_X1  g162(.A1(KEYINPUT0), .A2(G128), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n223), .A2(new_n242), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n242), .A2(G143), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n219), .A2(G146), .ZN(new_n355));
  AOI211_X1 g169(.A(new_n355), .B(new_n349), .C1(new_n233), .C2(G146), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n195), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n242), .A2(G143), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT1), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G128), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n358), .B(new_n361), .C1(new_n223), .C2(new_n242), .ZN(new_n362));
  OAI21_X1  g176(.A(G128), .B1(new_n355), .B2(new_n359), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT66), .ZN(new_n364));
  AOI21_X1  g178(.A(G146), .B1(new_n220), .B2(new_n222), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n363), .B(new_n364), .C1(new_n365), .C2(new_n352), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n353), .B1(new_n233), .B2(G146), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n364), .B1(new_n368), .B2(new_n363), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n362), .B(new_n204), .C1(new_n367), .C2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(KEYINPUT85), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n372));
  INV_X1    g186(.A(new_n362), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n352), .B1(new_n223), .B2(new_n242), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n306), .B1(new_n358), .B2(KEYINPUT1), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT66), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n373), .B1(new_n376), .B2(new_n366), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n372), .B1(new_n377), .B2(new_n204), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n357), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n217), .A2(G224), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT7), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n357), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n370), .A2(KEYINPUT85), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n377), .A2(new_n372), .A3(new_n204), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n382), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT87), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G110), .B(G122), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT8), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n321), .A2(G104), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n321), .A2(KEYINPUT76), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT76), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G107), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n395), .B1(new_n399), .B2(new_n188), .ZN(new_n400));
  INV_X1    g214(.A(G101), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n393), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n394), .B1(new_n312), .B2(G104), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT80), .A3(G101), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT75), .B1(new_n188), .B2(KEYINPUT3), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT75), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT3), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n406), .A2(new_n396), .A3(new_n398), .A4(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n408), .B1(G104), .B2(new_n321), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(G101), .B1(new_n188), .B2(G107), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G116), .B(G119), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT5), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n322), .A2(KEYINPUT5), .A3(G119), .ZN(new_n417));
  INV_X1    g231(.A(G113), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT2), .B(G113), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n416), .A2(new_n419), .B1(new_n421), .B2(new_n415), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n405), .A2(new_n414), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n422), .B1(new_n405), .B2(new_n414), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n392), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(KEYINPUT86), .B(new_n392), .C1(new_n423), .C2(new_n424), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n357), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n358), .B1(new_n223), .B2(new_n242), .ZN(new_n431));
  OAI22_X1  g245(.A1(new_n431), .A2(new_n349), .B1(new_n374), .B2(new_n350), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT84), .A3(new_n195), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n386), .B2(new_n385), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n427), .A2(new_n428), .B1(new_n435), .B2(new_n388), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n390), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n408), .A2(G104), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(KEYINPUT75), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n411), .B1(new_n441), .B2(new_n312), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n188), .A2(G107), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n401), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n414), .A2(KEYINPUT4), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT77), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n410), .A2(new_n443), .A3(new_n412), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G101), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT77), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT4), .A4(new_n414), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n415), .B(new_n420), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT78), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n447), .A2(KEYINPUT78), .A3(new_n453), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n423), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n391), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n438), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n437), .B1(new_n390), .B2(new_n436), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n459), .B2(new_n391), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n391), .B2(new_n459), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n435), .B(new_n381), .ZN(new_n467));
  OR3_X1    g281(.A1(new_n459), .A2(KEYINPUT6), .A3(new_n391), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n285), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n347), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n390), .A2(new_n436), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT88), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n460), .A3(new_n438), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n474), .A2(new_n285), .A3(new_n469), .A4(new_n346), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(KEYINPUT89), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G214), .B1(G237), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n347), .C1(new_n463), .C2(new_n470), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n345), .A2(new_n476), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G469), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT81), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n362), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n355), .B1(new_n233), .B2(G146), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(KEYINPUT81), .A3(new_n361), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n306), .B1(new_n351), .B2(KEYINPUT1), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n483), .B(new_n485), .C1(new_n486), .C2(new_n484), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n414), .A3(new_n405), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n405), .A2(new_n414), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n362), .B1(new_n367), .B2(new_n369), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT11), .B1(new_n310), .B2(G137), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT11), .ZN(new_n493));
  INV_X1    g307(.A(G137), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(G134), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT65), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n494), .B2(G134), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n310), .A2(KEYINPUT65), .A3(G137), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G131), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n498), .A2(new_n499), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n230), .A3(new_n496), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n491), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT12), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT67), .ZN(new_n507));
  INV_X1    g321(.A(new_n503), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n230), .B1(new_n502), .B2(new_n496), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n501), .A2(KEYINPUT67), .A3(new_n503), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(KEYINPUT12), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n491), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT10), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n377), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n489), .A2(new_n517), .B1(new_n488), .B2(new_n516), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n432), .B1(new_n456), .B2(new_n457), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n451), .A2(KEYINPUT79), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT79), .B1(new_n451), .B2(new_n519), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n512), .B(new_n518), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT82), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n451), .A2(new_n519), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT79), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n451), .A2(KEYINPUT79), .A3(new_n519), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n529), .A2(KEYINPUT82), .A3(new_n512), .A4(new_n518), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n515), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G110), .B(G140), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n217), .A2(G227), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n524), .A2(new_n530), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n512), .B1(new_n529), .B2(new_n518), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n535), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT83), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n538), .B1(new_n524), .B2(new_n530), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n543), .A2(KEYINPUT83), .A3(new_n535), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n481), .B(new_n285), .C1(new_n542), .C2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n481), .A2(new_n285), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n537), .A2(new_n535), .A3(new_n539), .ZN(new_n547));
  INV_X1    g361(.A(new_n515), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n535), .B1(new_n537), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n546), .B1(new_n550), .B2(G469), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G221), .ZN(new_n553));
  INV_X1    g367(.A(new_n330), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n554), .B2(new_n285), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n480), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT22), .B(G137), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n217), .A2(G221), .A3(G234), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n559), .B(new_n560), .Z(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT23), .ZN(new_n563));
  INV_X1    g377(.A(G119), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(G128), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n306), .A2(KEYINPUT23), .A3(G119), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n565), .B(new_n566), .C1(G119), .C2(new_n306), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G110), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT24), .B(G110), .Z(new_n569));
  XNOR2_X1  g383(.A(G119), .B(G128), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n269), .B2(new_n207), .ZN(new_n573));
  OAI22_X1  g387(.A1(new_n567), .A2(G110), .B1(new_n570), .B2(new_n569), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n243), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n262), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n562), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n572), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n261), .B2(new_n262), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n207), .A2(new_n243), .A3(new_n574), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n561), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n285), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT25), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n577), .A2(KEYINPUT25), .A3(new_n581), .A4(new_n285), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n331), .B1(G234), .B2(new_n285), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n586), .A2(KEYINPUT74), .A3(new_n587), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n587), .A2(G902), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n577), .A2(new_n581), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT70), .ZN(new_n595));
  INV_X1    g409(.A(G472), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n285), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT31), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n494), .A2(G134), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n310), .A2(G137), .ZN(new_n600));
  OAI21_X1  g414(.A(G131), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n503), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT68), .B1(new_n377), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT68), .ZN(new_n604));
  INV_X1    g418(.A(new_n602), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n490), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n354), .A2(new_n356), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n510), .A2(new_n607), .A3(new_n511), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n603), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT30), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n504), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT30), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n611), .B(new_n612), .C1(new_n377), .C2(new_n602), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n452), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n603), .A2(new_n606), .A3(new_n452), .A4(new_n608), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n216), .A2(new_n217), .A3(G210), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT27), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT26), .B(G101), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n598), .B1(new_n614), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n615), .A2(new_n619), .ZN(new_n622));
  INV_X1    g436(.A(new_n613), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(KEYINPUT30), .B2(new_n609), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n622), .B(KEYINPUT31), .C1(new_n624), .C2(new_n452), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n490), .A2(new_n605), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n608), .A2(new_n627), .A3(new_n452), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT28), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n628), .A2(KEYINPUT69), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT69), .B1(new_n628), .B2(new_n629), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n627), .A2(new_n611), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n615), .B1(new_n633), .B2(new_n452), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT28), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n619), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n597), .B1(new_n626), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n595), .B1(new_n639), .B2(KEYINPUT32), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT32), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n621), .A2(new_n625), .B1(new_n636), .B2(new_n637), .ZN(new_n642));
  OAI211_X1 g456(.A(KEYINPUT70), .B(new_n641), .C1(new_n642), .C2(new_n597), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n639), .A2(KEYINPUT32), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n615), .B1(new_n624), .B2(new_n452), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n637), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n632), .A2(new_n635), .A3(new_n619), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT29), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n628), .A2(new_n629), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT69), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n628), .A2(KEYINPUT69), .A3(new_n629), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n452), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n609), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n629), .B1(new_n656), .B2(new_n615), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n637), .A2(new_n648), .ZN(new_n659));
  AOI21_X1  g473(.A(G902), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n649), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G472), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n640), .A2(new_n643), .A3(new_n644), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT71), .ZN(new_n664));
  AOI22_X1  g478(.A1(G472), .A2(new_n661), .B1(new_n639), .B2(KEYINPUT32), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT71), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n640), .A4(new_n643), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n594), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n558), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G101), .ZN(G3));
  INV_X1    g484(.A(new_n639), .ZN(new_n671));
  AOI21_X1  g485(.A(G902), .B1(new_n626), .B2(new_n638), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n671), .B1(new_n596), .B2(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n557), .A2(new_n594), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n287), .B1(new_n281), .B2(new_n279), .ZN(new_n675));
  OAI21_X1  g489(.A(G475), .B1(new_n675), .B2(G902), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n276), .B1(new_n275), .B2(new_n277), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n282), .A2(KEYINPUT20), .A3(new_n283), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n299), .A2(new_n285), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n681), .B1(new_n340), .B2(G478), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n336), .B(KEYINPUT33), .Z(new_n683));
  AOI21_X1  g497(.A(new_n682), .B1(new_n683), .B2(G478), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n297), .ZN(new_n686));
  INV_X1    g500(.A(new_n477), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n471), .B2(new_n475), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n674), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT34), .B(G104), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G6));
  OAI211_X1 g506(.A(new_n342), .B(new_n676), .C1(new_n677), .C2(new_n678), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n297), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n674), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT35), .B(G107), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  AOI21_X1  g512(.A(KEYINPUT74), .B1(new_n586), .B2(new_n587), .ZN(new_n699));
  INV_X1    g513(.A(new_n587), .ZN(new_n700));
  AOI211_X1 g514(.A(new_n589), .B(new_n700), .C1(new_n584), .C2(new_n585), .ZN(new_n701));
  INV_X1    g515(.A(new_n592), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT97), .B1(new_n573), .B2(new_n576), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT97), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n579), .A2(new_n704), .A3(new_n580), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(KEYINPUT36), .B2(new_n562), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n703), .A2(new_n708), .A3(new_n705), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n702), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n699), .A2(new_n701), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n480), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n557), .A2(new_n673), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT37), .B(G110), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G12));
  NAND2_X1  g530(.A1(new_n664), .A2(new_n667), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n292), .B(KEYINPUT98), .Z(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(G900), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n719), .B1(new_n720), .B2(new_n295), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT99), .B1(new_n693), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n711), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT99), .ZN(new_n724));
  INV_X1    g538(.A(new_n721), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n289), .A2(new_n724), .A3(new_n342), .A4(new_n725), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n688), .A2(new_n722), .A3(new_n723), .A4(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n555), .B1(new_n545), .B2(new_n551), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n717), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G128), .ZN(G30));
  OAI21_X1  g544(.A(new_n622), .B1(new_n624), .B2(new_n452), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n619), .B1(new_n656), .B2(new_n615), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n731), .B1(KEYINPUT101), .B2(new_n732), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n732), .A2(KEYINPUT101), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n285), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n639), .A2(KEYINPUT32), .B1(new_n735), .B2(G472), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n736), .A2(new_n640), .A3(new_n643), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT102), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(new_n640), .A3(new_n643), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n342), .A2(new_n477), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n289), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n743), .A2(new_n723), .A3(new_n746), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n721), .B(KEYINPUT39), .Z(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n557), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n476), .A2(new_n479), .ZN(new_n754));
  XNOR2_X1  g568(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n747), .A2(new_n752), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n223), .ZN(G45));
  NAND3_X1  g572(.A1(new_n679), .A2(new_n684), .A3(new_n725), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n688), .A2(new_n760), .A3(new_n723), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n717), .A2(new_n728), .A3(new_n761), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT104), .B(G146), .Z(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G48));
  NAND2_X1  g578(.A1(new_n537), .A2(new_n539), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n541), .A3(new_n534), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT83), .B1(new_n543), .B2(new_n535), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n767), .A3(new_n536), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n768), .A2(new_n481), .A3(new_n285), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n481), .B1(new_n768), .B2(new_n285), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n769), .A2(new_n770), .A3(new_n555), .ZN(new_n771));
  INV_X1    g585(.A(new_n594), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n717), .A2(new_n771), .A3(new_n689), .A4(new_n772), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT41), .B(G113), .Z(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT105), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n773), .B(new_n775), .ZN(G15));
  NAND4_X1  g590(.A1(new_n717), .A2(new_n771), .A3(new_n772), .A4(new_n695), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G116), .ZN(G18));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n345), .A2(new_n723), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n664), .B2(new_n667), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n285), .B1(new_n542), .B2(new_n544), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(G469), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n556), .A3(new_n545), .A4(new_n688), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n779), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n781), .A2(new_n779), .A3(new_n785), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(KEYINPUT107), .B(G119), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G21));
  NAND2_X1  g605(.A1(new_n471), .A2(new_n475), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n745), .A3(new_n298), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n594), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n590), .A2(KEYINPUT109), .A3(new_n591), .A4(new_n593), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g613(.A(KEYINPUT108), .B(G472), .Z(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n654), .A2(new_n657), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n802), .A2(new_n637), .B1(new_n621), .B2(new_n625), .ZN(new_n803));
  OAI22_X1  g617(.A1(new_n672), .A2(new_n801), .B1(new_n803), .B2(new_n597), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n795), .B1(new_n799), .B2(new_n805), .ZN(new_n806));
  AOI211_X1 g620(.A(KEYINPUT110), .B(new_n804), .C1(new_n797), .C2(new_n798), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n771), .B(new_n794), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G122), .ZN(G24));
  NAND2_X1  g623(.A1(new_n759), .A2(KEYINPUT111), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n804), .A2(new_n711), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n679), .A2(new_n812), .A3(new_n684), .A4(new_n725), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n784), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(new_n191), .ZN(G27));
  NAND2_X1  g630(.A1(new_n556), .A2(new_n477), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(new_n476), .B2(new_n479), .ZN(new_n818));
  INV_X1    g632(.A(new_n546), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n537), .A2(new_n548), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n534), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT112), .B1(new_n531), .B2(new_n535), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n543), .A2(new_n535), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n823), .A3(G469), .A4(new_n824), .ZN(new_n825));
  AND4_X1   g639(.A1(KEYINPUT113), .A2(new_n545), .A3(new_n819), .A4(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n825), .A2(new_n819), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT113), .B1(new_n827), .B2(new_n545), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n818), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n665), .B1(KEYINPUT32), .B2(new_n639), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n799), .A3(new_n810), .A4(new_n813), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT42), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n825), .A2(new_n819), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n833), .B1(new_n769), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n827), .A2(KEYINPUT113), .A3(new_n545), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n810), .A2(new_n813), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(KEYINPUT42), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n837), .A2(new_n668), .A3(new_n818), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(new_n230), .ZN(G33));
  AND2_X1   g656(.A1(new_n722), .A2(new_n726), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n837), .A2(new_n668), .A3(new_n843), .A4(new_n818), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(G134), .ZN(G36));
  OAI21_X1  g659(.A(new_n824), .B1(new_n535), .B2(new_n531), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT45), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n481), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n848), .A2(KEYINPUT114), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(KEYINPUT114), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT45), .A4(new_n824), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n819), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT46), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n769), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n852), .A2(KEYINPUT46), .A3(new_n819), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n556), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT115), .B1(new_n858), .B2(new_n749), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n555), .B1(new_n855), .B2(new_n856), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n861), .A3(new_n748), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n289), .A2(new_n684), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT116), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT43), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n864), .A2(KEYINPUT116), .A3(KEYINPUT43), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n673), .A3(new_n723), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT44), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n687), .B1(new_n476), .B2(new_n479), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n863), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(G137), .ZN(G39));
  INV_X1    g691(.A(KEYINPUT47), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n858), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n860), .A2(KEYINPUT47), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR4_X1   g695(.A1(new_n717), .A2(new_n874), .A3(new_n772), .A4(new_n759), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(G140), .ZN(G42));
  NOR2_X1   g698(.A1(new_n769), .A2(new_n770), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n886), .A2(KEYINPUT49), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(KEYINPUT49), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n756), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n864), .A2(new_n817), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n743), .A3(new_n799), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n867), .A2(new_n719), .A3(new_n868), .ZN(new_n893));
  INV_X1    g707(.A(new_n806), .ZN(new_n894));
  INV_X1    g708(.A(new_n807), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n743), .A2(new_n772), .A3(new_n293), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n771), .A2(new_n873), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI221_X1 g714(.A(new_n290), .B1(new_n784), .B2(new_n897), .C1(new_n900), .C2(new_n685), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n830), .A2(new_n799), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n899), .A2(new_n902), .A3(new_n893), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT48), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NOR4_X1   g719(.A1(new_n898), .A2(new_n679), .A3(new_n684), .A4(new_n899), .ZN(new_n906));
  NOR4_X1   g720(.A1(new_n899), .A2(new_n893), .A3(new_n711), .A4(new_n804), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n756), .A2(new_n477), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n771), .A3(new_n896), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT50), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n885), .A2(new_n555), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n879), .A2(new_n880), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n897), .A2(new_n874), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n905), .B1(new_n918), .B2(KEYINPUT51), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT51), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n914), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n892), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n918), .A2(KEYINPUT51), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n921), .B1(new_n920), .B2(new_n914), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT123), .A4(new_n905), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n754), .A2(new_n477), .A3(new_n686), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n476), .A2(new_n694), .A3(new_n477), .A4(new_n479), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n929), .A2(new_n930), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n674), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n668), .A2(new_n558), .B1(new_n712), .B2(new_n713), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT118), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT118), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n940), .B(new_n818), .C1(new_n826), .C2(new_n828), .ZN(new_n941));
  NOR4_X1   g755(.A1(new_n711), .A2(new_n679), .A3(new_n342), .A4(new_n721), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n717), .A2(new_n728), .A3(new_n873), .A4(new_n942), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n832), .A3(new_n840), .A4(new_n844), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n668), .B(new_n771), .C1(new_n689), .C2(new_n695), .ZN(new_n946));
  INV_X1    g760(.A(new_n788), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n808), .B(new_n946), .C1(new_n947), .C2(new_n786), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n557), .B1(new_n667), .B2(new_n664), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n815), .B1(new_n950), .B2(new_n727), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT52), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n721), .A2(KEYINPUT119), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n721), .A2(KEYINPUT119), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n953), .A2(new_n556), .A3(new_n954), .ZN(new_n955));
  NOR4_X1   g769(.A1(new_n699), .A2(new_n701), .A3(new_n710), .A4(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n792), .A2(new_n745), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n737), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n826), .B2(new_n828), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n951), .A2(new_n952), .A3(new_n762), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n940), .A2(new_n771), .A3(new_n688), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n729), .A2(new_n762), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT52), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n939), .A2(new_n949), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n962), .A2(new_n951), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n969));
  OAI22_X1  g783(.A1(new_n968), .A2(KEYINPUT53), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT54), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n844), .A2(new_n941), .A3(new_n943), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n841), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n808), .A2(new_n773), .A3(new_n777), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n788), .B2(new_n787), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n973), .A2(new_n975), .A3(new_n963), .A4(new_n960), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT118), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n977), .A2(new_n936), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n969), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT121), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT54), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n964), .A2(new_n948), .A3(new_n945), .ZN(new_n982));
  INV_X1    g796(.A(new_n967), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n982), .A2(KEYINPUT53), .A3(new_n939), .A4(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT121), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n985), .B(new_n969), .C1(new_n976), .C2(new_n978), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n980), .A2(new_n981), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n971), .A2(KEYINPUT122), .A3(new_n987), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n987), .A2(KEYINPUT122), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n927), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(G952), .A2(G953), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n891), .B1(new_n990), .B2(new_n991), .ZN(G75));
  NAND3_X1  g806(.A1(new_n980), .A2(new_n984), .A3(new_n986), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(G210), .A3(G902), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT56), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n466), .A2(new_n468), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(new_n467), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT55), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n994), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n998), .B1(new_n994), .B2(new_n995), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n217), .A2(G952), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(G51));
  INV_X1    g816(.A(new_n852), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n993), .A2(G902), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n768), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n984), .A2(new_n986), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n985), .B1(new_n966), .B2(new_n969), .ZN(new_n1008));
  OAI21_X1  g822(.A(KEYINPUT54), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n987), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n546), .B(KEYINPUT57), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1006), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1005), .B1(new_n1012), .B2(KEYINPUT124), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT124), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1011), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n1009), .B2(new_n987), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1014), .B1(new_n1016), .B2(new_n1006), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1001), .B1(new_n1013), .B2(new_n1017), .ZN(G54));
  NAND2_X1  g832(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT125), .Z(new_n1020));
  NAND3_X1  g834(.A1(new_n993), .A2(G902), .A3(new_n1020), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1021), .A2(new_n282), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1021), .A2(new_n282), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n1022), .A2(new_n1023), .A3(new_n1001), .ZN(G60));
  XNOR2_X1  g838(.A(new_n680), .B(KEYINPUT59), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n683), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1010), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1001), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1025), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n988), .A2(new_n989), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1029), .B1(new_n683), .B2(new_n1031), .ZN(G63));
  NAND2_X1  g846(.A1(G217), .A2(G902), .ZN(new_n1033));
  XOR2_X1   g847(.A(new_n1033), .B(KEYINPUT60), .Z(new_n1034));
  NAND2_X1  g848(.A1(new_n993), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n577), .A2(new_n581), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n707), .A2(new_n709), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n993), .A2(new_n1038), .A3(new_n1034), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1037), .A2(new_n1028), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT61), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n1040), .B(new_n1041), .ZN(G66));
  INV_X1    g856(.A(G224), .ZN(new_n1043));
  OAI21_X1  g857(.A(G953), .B1(new_n296), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n939), .A2(new_n975), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1044), .B1(new_n1046), .B2(G953), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n996), .B1(G898), .B2(new_n217), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1047), .B(new_n1048), .ZN(G69));
  AOI22_X1  g863(.A1(new_n863), .A2(new_n875), .B1(new_n881), .B2(new_n882), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n685), .A2(new_n693), .ZN(new_n1051));
  AND4_X1   g865(.A1(new_n668), .A2(new_n750), .A3(new_n873), .A4(new_n1051), .ZN(new_n1052));
  AND2_X1   g866(.A1(new_n951), .A2(new_n762), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n757), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g868(.A(KEYINPUT62), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n757), .A2(new_n1053), .A3(KEYINPUT62), .ZN(new_n1057));
  AOI21_X1  g871(.A(new_n1052), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1050), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1059), .A2(new_n217), .ZN(new_n1060));
  XOR2_X1   g874(.A(new_n624), .B(new_n213), .Z(new_n1061));
  NAND3_X1  g875(.A1(new_n1060), .A2(KEYINPUT126), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g876(.A(KEYINPUT126), .ZN(new_n1063));
  AOI21_X1  g877(.A(G953), .B1(new_n1050), .B2(new_n1058), .ZN(new_n1064));
  INV_X1    g878(.A(new_n1061), .ZN(new_n1065));
  OAI21_X1  g879(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n217), .B1(G227), .B2(G900), .ZN(new_n1068));
  OR2_X1    g882(.A1(new_n1068), .A2(KEYINPUT127), .ZN(new_n1069));
  NAND2_X1  g883(.A1(new_n1053), .A2(new_n844), .ZN(new_n1070));
  AOI211_X1 g884(.A(new_n746), .B(new_n902), .C1(new_n471), .C2(new_n475), .ZN(new_n1071));
  AOI211_X1 g885(.A(new_n841), .B(new_n1070), .C1(new_n863), .C2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g886(.A1(new_n1072), .A2(new_n217), .A3(new_n1050), .ZN(new_n1073));
  AOI21_X1  g887(.A(new_n1061), .B1(G900), .B2(G953), .ZN(new_n1074));
  AOI22_X1  g888(.A1(new_n1073), .A2(new_n1074), .B1(KEYINPUT127), .B2(new_n1068), .ZN(new_n1075));
  NAND3_X1  g889(.A1(new_n1067), .A2(new_n1069), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g890(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g891(.A(new_n1069), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1078));
  NOR2_X1   g892(.A1(new_n1077), .A2(new_n1078), .ZN(G72));
  NAND3_X1  g893(.A1(new_n1072), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1080));
  NAND2_X1  g894(.A1(G472), .A2(G902), .ZN(new_n1081));
  XOR2_X1   g895(.A(new_n1081), .B(KEYINPUT63), .Z(new_n1082));
  AOI211_X1 g896(.A(new_n619), .B(new_n645), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g897(.A1(new_n646), .A2(new_n731), .ZN(new_n1084));
  AND3_X1   g898(.A1(new_n970), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g899(.A1(new_n645), .A2(new_n619), .ZN(new_n1086));
  NAND3_X1  g900(.A1(new_n1050), .A2(new_n1046), .A3(new_n1058), .ZN(new_n1087));
  AOI21_X1  g901(.A(new_n1086), .B1(new_n1087), .B2(new_n1082), .ZN(new_n1088));
  NOR4_X1   g902(.A1(new_n1083), .A2(new_n1085), .A3(new_n1088), .A4(new_n1001), .ZN(G57));
endmodule


