

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587;

  XOR2_X1 U320 ( .A(G127GAT), .B(G15GAT), .Z(n439) );
  INV_X1 U321 ( .A(n379), .ZN(n352) );
  AND2_X1 U322 ( .A1(G227GAT), .A2(G233GAT), .ZN(n288) );
  XNOR2_X1 U323 ( .A(n356), .B(KEYINPUT64), .ZN(n357) );
  XNOR2_X1 U324 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U325 ( .A(n390), .B(KEYINPUT48), .ZN(n391) );
  OR2_X1 U326 ( .A1(n567), .A2(n434), .ZN(n436) );
  XNOR2_X1 U327 ( .A(n392), .B(n391), .ZN(n531) );
  XNOR2_X1 U328 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U329 ( .A(n443), .B(n288), .ZN(n444) );
  XNOR2_X1 U330 ( .A(n355), .B(n354), .ZN(n381) );
  XNOR2_X1 U331 ( .A(n445), .B(n444), .ZN(n446) );
  INV_X1 U332 ( .A(G43GAT), .ZN(n478) );
  XNOR2_X1 U333 ( .A(n477), .B(n476), .ZN(n505) );
  XNOR2_X1 U334 ( .A(n450), .B(G176GAT), .ZN(n451) );
  XNOR2_X1 U335 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U336 ( .A(n452), .B(n451), .ZN(G1349GAT) );
  XNOR2_X1 U337 ( .A(n481), .B(n480), .ZN(G1330GAT) );
  XNOR2_X1 U338 ( .A(G85GAT), .B(KEYINPUT72), .ZN(n289) );
  XNOR2_X1 U339 ( .A(n289), .B(G92GAT), .ZN(n335) );
  XNOR2_X1 U340 ( .A(G148GAT), .B(G106GAT), .ZN(n290) );
  XNOR2_X1 U341 ( .A(n290), .B(G78GAT), .ZN(n428) );
  XNOR2_X1 U342 ( .A(n335), .B(n428), .ZN(n302) );
  XOR2_X1 U343 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n292) );
  NAND2_X1 U344 ( .A1(G230GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U346 ( .A(n293), .B(KEYINPUT31), .Z(n297) );
  XNOR2_X1 U347 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n294) );
  XNOR2_X1 U348 ( .A(n294), .B(KEYINPUT71), .ZN(n320) );
  XNOR2_X1 U349 ( .A(G120GAT), .B(G99GAT), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n295), .B(G71GAT), .ZN(n437) );
  XNOR2_X1 U351 ( .A(n320), .B(n437), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U353 ( .A(n298), .B(KEYINPUT33), .Z(n300) );
  XOR2_X1 U354 ( .A(G64GAT), .B(G204GAT), .Z(n308) );
  XNOR2_X1 U355 ( .A(G176GAT), .B(n308), .ZN(n299) );
  XNOR2_X1 U356 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n576) );
  XNOR2_X1 U358 ( .A(n576), .B(KEYINPUT41), .ZN(n552) );
  INV_X1 U359 ( .A(KEYINPUT54), .ZN(n394) );
  XOR2_X1 U360 ( .A(KEYINPUT88), .B(G197GAT), .Z(n304) );
  XNOR2_X1 U361 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U363 ( .A(G211GAT), .B(n305), .Z(n430) );
  XOR2_X1 U364 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n307) );
  NAND2_X1 U365 ( .A1(G226GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U366 ( .A(n307), .B(n306), .ZN(n311) );
  XNOR2_X1 U367 ( .A(G36GAT), .B(G92GAT), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U369 ( .A(n311), .B(n310), .Z(n318) );
  XOR2_X1 U370 ( .A(G169GAT), .B(KEYINPUT17), .Z(n313) );
  XNOR2_X1 U371 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U373 ( .A(n314), .B(KEYINPUT18), .Z(n316) );
  XNOR2_X1 U374 ( .A(G190GAT), .B(G176GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n447) );
  XNOR2_X1 U376 ( .A(G8GAT), .B(n447), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U378 ( .A(n430), .B(n319), .Z(n522) );
  XOR2_X1 U379 ( .A(G155GAT), .B(G22GAT), .Z(n421) );
  XNOR2_X1 U380 ( .A(n421), .B(n439), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n321), .B(n320), .ZN(n326) );
  XNOR2_X1 U382 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n322), .B(G8GAT), .ZN(n370) );
  XOR2_X1 U384 ( .A(KEYINPUT12), .B(n370), .Z(n324) );
  NAND2_X1 U385 ( .A1(G231GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U387 ( .A(n326), .B(n325), .Z(n334) );
  XOR2_X1 U388 ( .A(G71GAT), .B(G183GAT), .Z(n328) );
  XNOR2_X1 U389 ( .A(G78GAT), .B(G211GAT), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U391 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n330) );
  XNOR2_X1 U392 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U395 ( .A(n334), .B(n333), .Z(n558) );
  XOR2_X1 U396 ( .A(n335), .B(G99GAT), .Z(n337) );
  NAND2_X1 U397 ( .A1(G232GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U399 ( .A(G134GAT), .B(G43GAT), .Z(n443) );
  XOR2_X1 U400 ( .A(n443), .B(KEYINPUT76), .Z(n340) );
  XNOR2_X1 U401 ( .A(G162GAT), .B(G50GAT), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n338), .B(KEYINPUT75), .ZN(n425) );
  XNOR2_X1 U403 ( .A(G218GAT), .B(n425), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n355) );
  XOR2_X1 U406 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n344) );
  XNOR2_X1 U407 ( .A(KEYINPUT79), .B(KEYINPUT11), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U409 ( .A(G106GAT), .B(G190GAT), .Z(n346) );
  XNOR2_X1 U410 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n345) );
  XNOR2_X1 U411 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U412 ( .A(n348), .B(n347), .Z(n353) );
  XOR2_X1 U413 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n350) );
  XNOR2_X1 U414 ( .A(KEYINPUT68), .B(G36GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U416 ( .A(G29GAT), .B(n351), .ZN(n379) );
  XOR2_X1 U417 ( .A(KEYINPUT36), .B(n381), .Z(n585) );
  AND2_X1 U418 ( .A1(n558), .A2(n585), .ZN(n358) );
  INV_X1 U419 ( .A(KEYINPUT45), .ZN(n356) );
  NOR2_X1 U420 ( .A1(n359), .A2(n576), .ZN(n361) );
  INV_X1 U421 ( .A(KEYINPUT113), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n380) );
  XOR2_X1 U423 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n363) );
  XNOR2_X1 U424 ( .A(KEYINPUT65), .B(KEYINPUT70), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n377) );
  XOR2_X1 U426 ( .A(G197GAT), .B(G22GAT), .Z(n365) );
  XNOR2_X1 U427 ( .A(G141GAT), .B(G113GAT), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U429 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n367) );
  XNOR2_X1 U430 ( .A(G15GAT), .B(G169GAT), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U432 ( .A(n369), .B(n368), .Z(n375) );
  XOR2_X1 U433 ( .A(n370), .B(G43GAT), .Z(n372) );
  NAND2_X1 U434 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U436 ( .A(G50GAT), .B(n373), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U438 ( .A(n377), .B(n376), .Z(n378) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n571) );
  NAND2_X1 U440 ( .A1(n380), .A2(n571), .ZN(n389) );
  INV_X1 U441 ( .A(n381), .ZN(n560) );
  INV_X1 U442 ( .A(n558), .ZN(n582) );
  NOR2_X1 U443 ( .A1(n571), .A2(n552), .ZN(n383) );
  XNOR2_X1 U444 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n384) );
  NAND2_X1 U446 ( .A1(n582), .A2(n384), .ZN(n385) );
  NOR2_X1 U447 ( .A1(n560), .A2(n385), .ZN(n387) );
  XNOR2_X1 U448 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n387), .B(n386), .ZN(n388) );
  NAND2_X1 U450 ( .A1(n389), .A2(n388), .ZN(n392) );
  INV_X1 U451 ( .A(KEYINPUT114), .ZN(n390) );
  NOR2_X1 U452 ( .A1(n522), .A2(n531), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n567) );
  XOR2_X1 U454 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n396) );
  XNOR2_X1 U455 ( .A(KEYINPUT90), .B(KEYINPUT92), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n402) );
  XOR2_X1 U457 ( .A(G141GAT), .B(KEYINPUT2), .Z(n398) );
  XNOR2_X1 U458 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n431) );
  XOR2_X1 U460 ( .A(n431), .B(KEYINPUT4), .Z(n400) );
  NAND2_X1 U461 ( .A1(G225GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n417) );
  XOR2_X1 U464 ( .A(G127GAT), .B(G120GAT), .Z(n404) );
  XNOR2_X1 U465 ( .A(G148GAT), .B(G155GAT), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U467 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n406) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(G57GAT), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U470 ( .A(n408), .B(n407), .Z(n415) );
  XOR2_X1 U471 ( .A(G113GAT), .B(KEYINPUT83), .Z(n410) );
  XNOR2_X1 U472 ( .A(KEYINPUT82), .B(KEYINPUT0), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n438) );
  XOR2_X1 U474 ( .A(G85GAT), .B(n438), .Z(n412) );
  XNOR2_X1 U475 ( .A(G29GAT), .B(G134GAT), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U477 ( .A(G162GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U479 ( .A(n417), .B(n416), .Z(n566) );
  INV_X1 U480 ( .A(n566), .ZN(n519) );
  XOR2_X1 U481 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n419) );
  XNOR2_X1 U482 ( .A(KEYINPUT86), .B(G204GAT), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U484 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U487 ( .A(n424), .B(KEYINPUT23), .Z(n427) );
  XNOR2_X1 U488 ( .A(n425), .B(KEYINPUT87), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U490 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n465) );
  NAND2_X1 U493 ( .A1(n519), .A2(n465), .ZN(n434) );
  XNOR2_X1 U494 ( .A(KEYINPUT122), .B(KEYINPUT55), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n448) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n439), .B(KEYINPUT20), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n440), .B(KEYINPUT84), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n445) );
  XOR2_X1 U500 ( .A(n447), .B(n446), .Z(n533) );
  INV_X1 U501 ( .A(n533), .ZN(n463) );
  AND2_X1 U502 ( .A1(n448), .A2(n463), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n449), .B(KEYINPUT123), .ZN(n564) );
  NOR2_X1 U504 ( .A1(n552), .A2(n564), .ZN(n452) );
  XNOR2_X1 U505 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n450) );
  XOR2_X1 U506 ( .A(KEYINPUT105), .B(KEYINPUT38), .Z(n477) );
  NOR2_X1 U507 ( .A1(n576), .A2(n571), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n453), .B(KEYINPUT74), .ZN(n490) );
  XNOR2_X1 U509 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n475) );
  INV_X1 U510 ( .A(n522), .ZN(n457) );
  NAND2_X1 U511 ( .A1(n463), .A2(n457), .ZN(n454) );
  XNOR2_X1 U512 ( .A(KEYINPUT96), .B(n454), .ZN(n455) );
  NAND2_X1 U513 ( .A1(n455), .A2(n465), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT25), .ZN(n460) );
  XOR2_X1 U515 ( .A(n457), .B(KEYINPUT27), .Z(n464) );
  NOR2_X1 U516 ( .A1(n465), .A2(n463), .ZN(n458) );
  XOR2_X1 U517 ( .A(KEYINPUT26), .B(n458), .Z(n568) );
  NOR2_X1 U518 ( .A1(n464), .A2(n568), .ZN(n459) );
  NOR2_X1 U519 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT97), .ZN(n462) );
  NAND2_X1 U521 ( .A1(n462), .A2(n519), .ZN(n470) );
  XNOR2_X1 U522 ( .A(n463), .B(KEYINPUT85), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n519), .A2(n464), .ZN(n529) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT28), .ZN(n535) );
  NAND2_X1 U525 ( .A1(n529), .A2(n535), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n466), .B(KEYINPUT95), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT98), .ZN(n488) );
  NAND2_X1 U530 ( .A1(n488), .A2(n582), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n472), .B(KEYINPUT103), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n473), .A2(n585), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n475), .B(n474), .ZN(n517) );
  NAND2_X1 U534 ( .A1(n490), .A2(n517), .ZN(n476) );
  NOR2_X1 U535 ( .A1(n533), .A2(n505), .ZN(n481) );
  XNOR2_X1 U536 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n479) );
  NOR2_X1 U537 ( .A1(n564), .A2(n381), .ZN(n483) );
  XNOR2_X1 U538 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n483), .B(n482), .ZN(n485) );
  INV_X1 U540 ( .A(G190GAT), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n485), .B(n484), .ZN(G1351GAT) );
  NAND2_X1 U542 ( .A1(n558), .A2(n381), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n486), .B(KEYINPUT16), .ZN(n487) );
  XNOR2_X1 U544 ( .A(KEYINPUT81), .B(n487), .ZN(n489) );
  AND2_X1 U545 ( .A1(n489), .A2(n488), .ZN(n508) );
  NAND2_X1 U546 ( .A1(n508), .A2(n490), .ZN(n499) );
  NOR2_X1 U547 ( .A1(n519), .A2(n499), .ZN(n492) );
  XNOR2_X1 U548 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(n493), .ZN(G1324GAT) );
  NOR2_X1 U551 ( .A1(n522), .A2(n499), .ZN(n494) );
  XOR2_X1 U552 ( .A(KEYINPUT100), .B(n494), .Z(n495) );
  XNOR2_X1 U553 ( .A(G8GAT), .B(n495), .ZN(G1325GAT) );
  NOR2_X1 U554 ( .A1(n533), .A2(n499), .ZN(n497) );
  XNOR2_X1 U555 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U557 ( .A(G15GAT), .B(n498), .Z(G1326GAT) );
  NOR2_X1 U558 ( .A1(n535), .A2(n499), .ZN(n500) );
  XOR2_X1 U559 ( .A(KEYINPUT102), .B(n500), .Z(n501) );
  XNOR2_X1 U560 ( .A(G22GAT), .B(n501), .ZN(G1327GAT) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n503) );
  NOR2_X1 U562 ( .A1(n519), .A2(n505), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n522), .A2(n505), .ZN(n504) );
  XOR2_X1 U565 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  NOR2_X1 U566 ( .A1(n505), .A2(n535), .ZN(n506) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n506), .Z(G1331GAT) );
  INV_X1 U568 ( .A(n571), .ZN(n548) );
  NOR2_X1 U569 ( .A1(n548), .A2(n552), .ZN(n507) );
  XOR2_X1 U570 ( .A(KEYINPUT107), .B(n507), .Z(n518) );
  NAND2_X1 U571 ( .A1(n518), .A2(n508), .ZN(n513) );
  NOR2_X1 U572 ( .A1(n519), .A2(n513), .ZN(n509) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n509), .Z(n510) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n522), .A2(n513), .ZN(n511) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n533), .A2(n513), .ZN(n512) );
  XOR2_X1 U578 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U579 ( .A1(n535), .A2(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n526) );
  NOR2_X1 U584 ( .A1(n519), .A2(n526), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n526), .ZN(n523) );
  XOR2_X1 U588 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U589 ( .A1(n533), .A2(n526), .ZN(n524) );
  XOR2_X1 U590 ( .A(KEYINPUT110), .B(n524), .Z(n525) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  NOR2_X1 U592 ( .A1(n535), .A2(n526), .ZN(n527) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(n527), .Z(n528) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  INV_X1 U595 ( .A(n529), .ZN(n530) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U597 ( .A(KEYINPUT115), .B(n532), .ZN(n547) );
  NOR2_X1 U598 ( .A1(n533), .A2(n547), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n534), .B(KEYINPUT116), .ZN(n536) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n544) );
  NOR2_X1 U601 ( .A1(n571), .A2(n544), .ZN(n537) );
  XOR2_X1 U602 ( .A(G113GAT), .B(n537), .Z(G1340GAT) );
  NOR2_X1 U603 ( .A1(n552), .A2(n544), .ZN(n539) );
  XNOR2_X1 U604 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U606 ( .A(G120GAT), .B(n540), .Z(G1341GAT) );
  NOR2_X1 U607 ( .A1(n582), .A2(n544), .ZN(n542) );
  XNOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U610 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  NOR2_X1 U611 ( .A1(n381), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n550) );
  NOR2_X1 U615 ( .A1(n568), .A2(n547), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n561), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT121), .Z(n555) );
  INV_X1 U620 ( .A(n552), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n561), .A2(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U623 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n561), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U629 ( .A1(n571), .A2(n564), .ZN(n563) );
  XOR2_X1 U630 ( .A(G169GAT), .B(n563), .Z(G1348GAT) );
  NOR2_X1 U631 ( .A1(n582), .A2(n564), .ZN(n565) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n565), .Z(G1350GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n570) );
  INV_X1 U634 ( .A(n568), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n581) );
  NOR2_X1 U636 ( .A1(n571), .A2(n581), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n575) );
  XOR2_X1 U639 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  INV_X1 U641 ( .A(n581), .ZN(n584) );
  AND2_X1 U642 ( .A1(n584), .A2(n576), .ZN(n580) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n578) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(G211GAT), .B(n583), .Z(G1354GAT) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

