//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT11), .A2(G134), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G137), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n196), .A2(KEYINPUT65), .A3(KEYINPUT11), .A4(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G134), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n202), .A3(G137), .ZN(new_n203));
  AOI21_X1  g017(.A(G137), .B1(new_n200), .B2(new_n202), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n198), .B(new_n203), .C1(new_n204), .C2(KEYINPUT11), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G131), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT64), .B(G134), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G137), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n209), .A2(new_n210), .A3(new_n198), .A4(new_n203), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT78), .A2(G104), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT78), .A2(G104), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n213), .A2(new_n214), .A3(G107), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n216), .B1(G104), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT81), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n214), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n221));
  INV_X1    g035(.A(G107), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT78), .A2(G104), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G107), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G107), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n226), .B1(G104), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n228), .A3(new_n216), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n220), .A2(new_n222), .A3(new_n224), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(new_n217), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n219), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G143), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT1), .A3(G146), .ZN(new_n235));
  XNOR2_X1  g049(.A(G143), .B(G146), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G128), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n239));
  INV_X1    g053(.A(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G143), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n234), .A2(G146), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n236), .A2(KEYINPUT66), .A3(new_n239), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n237), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n233), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n233), .A2(new_n247), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n212), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT82), .B1(new_n233), .B2(new_n247), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT10), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT10), .ZN(new_n255));
  OAI211_X1 g069(.A(KEYINPUT82), .B(new_n255), .C1(new_n233), .C2(new_n247), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n212), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT79), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n213), .A2(new_n227), .A3(new_n214), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n221), .A2(new_n222), .A3(G104), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT3), .A2(G107), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n259), .B(G101), .C1(new_n260), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT4), .A3(new_n229), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n216), .B1(new_n225), .B2(new_n228), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(new_n259), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT80), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n229), .A2(KEYINPUT4), .ZN(new_n269));
  OAI21_X1  g083(.A(G101), .B1(new_n260), .B2(new_n263), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT79), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT80), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n269), .A2(new_n271), .A3(new_n272), .A4(new_n264), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n266), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n241), .A2(new_n242), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT0), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n238), .ZN(new_n279));
  NOR2_X1   g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n236), .B1(new_n278), .B2(new_n238), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n276), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n274), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n257), .A2(new_n258), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n192), .B1(new_n252), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n258), .B1(new_n257), .B2(new_n286), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n254), .A2(new_n256), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n284), .B1(new_n268), .B2(new_n273), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n191), .B1(new_n292), .B2(new_n258), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT83), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n289), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n290), .A2(new_n291), .A3(new_n212), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT83), .B1(new_n296), .B2(new_n191), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n288), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n187), .B(G469), .C1(new_n298), .C2(G902), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT85), .B1(new_n296), .B2(new_n191), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n287), .A2(new_n301), .A3(new_n192), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n252), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n191), .B1(new_n289), .B2(new_n296), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT86), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n212), .B1(new_n290), .B2(new_n291), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n287), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT86), .A3(new_n191), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n303), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G469), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n252), .A2(new_n287), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n191), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n287), .A2(new_n294), .A3(new_n192), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n307), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n293), .A2(new_n294), .ZN(new_n318));
  OAI211_X1 g132(.A(G469), .B(new_n315), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(G469), .A2(G902), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(KEYINPUT84), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n299), .A2(new_n313), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G221), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT9), .B(G234), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n323), .B1(new_n325), .B2(new_n312), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n326), .B(KEYINPUT77), .Z(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT87), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n322), .A2(KEYINPUT87), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G234), .ZN(new_n334));
  OAI21_X1  g148(.A(G217), .B1(new_n334), .B2(G902), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT74), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n337), .A2(KEYINPUT16), .A3(G140), .ZN(new_n338));
  XNOR2_X1  g152(.A(G125), .B(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT16), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n338), .A2(new_n341), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G146), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n240), .B1(new_n342), .B2(new_n343), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(KEYINPUT76), .A3(new_n346), .ZN(new_n347));
  OR3_X1    g161(.A1(new_n344), .A2(KEYINPUT76), .A3(G146), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n238), .A2(G119), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n238), .A2(G119), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT24), .B(G110), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT23), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n238), .A2(KEYINPUT23), .A3(G119), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n355), .A2(new_n349), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G110), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n347), .A2(new_n348), .A3(new_n353), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n358), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n351), .A2(new_n352), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n361), .A2(new_n362), .B1(new_n240), .B2(new_n339), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n345), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT22), .B(G137), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n323), .A2(new_n334), .A3(G953), .ZN(new_n367));
  XOR2_X1   g181(.A(new_n366), .B(new_n367), .Z(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n360), .B2(new_n364), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT25), .B1(new_n372), .B2(new_n312), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n374));
  NOR4_X1   g188(.A1(new_n370), .A2(new_n371), .A3(new_n374), .A4(G902), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n336), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n372), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n335), .A2(new_n312), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G472), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n245), .A2(new_n246), .ZN(new_n381));
  INV_X1    g195(.A(new_n237), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n199), .A2(G137), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(new_n208), .B2(G137), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n381), .A2(new_n382), .B1(G131), .B2(new_n384), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n212), .A2(new_n283), .B1(new_n385), .B2(new_n211), .ZN(new_n386));
  OR2_X1    g200(.A1(KEYINPUT67), .A2(KEYINPUT30), .ZN(new_n387));
  NAND2_X1  g201(.A1(KEYINPUT67), .A2(KEYINPUT30), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n211), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n384), .A2(G131), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n390), .A2(new_n247), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n283), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n393), .B1(new_n206), .B2(new_n211), .ZN(new_n394));
  OAI211_X1 g208(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n392), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT2), .B(G113), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G116), .B(G119), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n212), .A2(new_n283), .ZN(new_n404));
  INV_X1    g218(.A(new_n402), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n385), .A2(new_n211), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT26), .B(G101), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G237), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n189), .A3(G210), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT69), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n411), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT73), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT73), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n408), .A2(new_n418), .A3(new_n415), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n392), .A2(new_n394), .A3(new_n402), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(KEYINPUT28), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n386), .A2(new_n405), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n422), .A2(new_n420), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n421), .B1(new_n423), .B2(KEYINPUT28), .ZN(new_n424));
  INV_X1    g238(.A(new_n415), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT29), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n419), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT28), .B1(new_n422), .B2(new_n420), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(KEYINPUT28), .B2(new_n420), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(new_n415), .ZN(new_n430));
  AOI21_X1  g244(.A(G902), .B1(new_n430), .B2(KEYINPUT29), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n380), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT71), .ZN(new_n433));
  AOI211_X1 g247(.A(KEYINPUT70), .B(new_n415), .C1(new_n386), .C2(new_n405), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT70), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n407), .B2(new_n425), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n405), .B1(new_n389), .B2(new_n395), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n403), .B(KEYINPUT71), .C1(new_n436), .C2(new_n434), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT31), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT72), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT70), .B1(new_n420), .B2(new_n415), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n407), .A2(new_n435), .A3(new_n425), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n438), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT31), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n445), .A2(new_n446), .B1(new_n429), .B2(new_n415), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n441), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n442), .B1(new_n441), .B2(new_n447), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT32), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n451), .A2(G472), .A3(G902), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n432), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n441), .A2(new_n447), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT72), .ZN(new_n455));
  NOR2_X1   g269(.A1(G472), .A2(G902), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n441), .A2(new_n447), .A3(new_n442), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n451), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n379), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(G475), .A2(G902), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n461), .B(KEYINPUT93), .Z(new_n462));
  NAND3_X1  g276(.A1(new_n412), .A2(new_n189), .A3(G214), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n234), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(KEYINPUT18), .B2(G131), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n463), .B(G143), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT18), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n466), .A2(new_n467), .A3(new_n210), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n339), .B(G146), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n347), .A2(new_n348), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n464), .A2(G131), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT17), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT91), .B1(new_n464), .B2(G131), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT91), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n466), .A2(new_n476), .A3(new_n210), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n475), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n474), .B1(new_n478), .B2(new_n473), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n470), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  INV_X1    g295(.A(G104), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT19), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n339), .B(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(G146), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(new_n344), .B2(G146), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n475), .A2(new_n472), .A3(new_n477), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n470), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n485), .B1(new_n491), .B2(new_n483), .ZN(new_n492));
  INV_X1    g306(.A(new_n483), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n489), .A2(new_n490), .ZN(new_n494));
  OAI211_X1 g308(.A(KEYINPUT92), .B(new_n493), .C1(new_n494), .C2(new_n470), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n462), .B1(new_n484), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT20), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT20), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(new_n462), .C1(new_n484), .C2(new_n496), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT94), .ZN(new_n501));
  OR3_X1    g315(.A1(new_n480), .A2(new_n501), .A3(new_n483), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n501), .B1(new_n480), .B2(new_n483), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n502), .B(new_n312), .C1(new_n484), .C2(new_n503), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n498), .A2(new_n500), .B1(new_n504), .B2(G475), .ZN(new_n505));
  INV_X1    g319(.A(G952), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(G953), .ZN(new_n507));
  NAND2_X1  g321(.A1(G234), .A2(G237), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT21), .B(G898), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(G902), .A3(G953), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n234), .A2(G128), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n238), .A2(G143), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n516), .B(new_n208), .Z(new_n517));
  INV_X1    g331(.A(G116), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT14), .A3(G122), .ZN(new_n519));
  XNOR2_X1  g333(.A(G116), .B(G122), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(G107), .B(new_n519), .C1(new_n521), .C2(KEYINPUT14), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n517), .B(new_n522), .C1(G107), .C2(new_n521), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT13), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n515), .B1(new_n514), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT13), .B1(new_n234), .B2(G128), .ZN(new_n526));
  OAI21_X1  g340(.A(G134), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT95), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n208), .A2(new_n514), .A3(new_n515), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n521), .A2(G107), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n520), .A2(new_n222), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n523), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n325), .A2(G217), .A3(new_n189), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n312), .ZN(new_n536));
  INV_X1    g350(.A(G478), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(KEYINPUT15), .ZN(new_n538));
  XOR2_X1   g352(.A(new_n536), .B(new_n538), .Z(new_n539));
  NAND3_X1  g353(.A1(new_n505), .A2(new_n513), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G214), .B1(G237), .B2(G902), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n402), .A2(new_n276), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n274), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n399), .A2(KEYINPUT5), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n518), .A2(G119), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n544), .B(G113), .C1(KEYINPUT5), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n401), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(new_n233), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G110), .B(G122), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n543), .A2(new_n552), .A3(new_n550), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(KEYINPUT6), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT88), .B1(new_n393), .B2(G125), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n247), .A2(new_n337), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n393), .A2(KEYINPUT88), .A3(G125), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT89), .ZN(new_n562));
  INV_X1    g376(.A(G224), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n562), .B1(new_n563), .B2(G953), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n189), .A2(KEYINPUT89), .A3(G224), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n566), .B(KEYINPUT90), .Z(new_n567));
  XOR2_X1   g381(.A(new_n561), .B(new_n567), .Z(new_n568));
  INV_X1    g382(.A(KEYINPUT6), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n551), .A2(new_n569), .A3(new_n553), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n556), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G210), .B1(G237), .B2(G902), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n564), .A2(KEYINPUT7), .A3(new_n565), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n559), .A2(new_n560), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n559), .B2(new_n560), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n552), .B(KEYINPUT8), .Z(new_n576));
  NAND2_X1  g390(.A1(new_n548), .A2(new_n233), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n550), .B2(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n579), .B2(new_n555), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n571), .A2(new_n572), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n572), .B1(new_n571), .B2(new_n580), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n541), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n540), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n333), .A2(new_n460), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  NAND3_X1  g401(.A1(new_n455), .A2(new_n312), .A3(new_n457), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G472), .ZN(new_n589));
  INV_X1    g403(.A(new_n379), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n458), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n541), .ZN(new_n593));
  INV_X1    g407(.A(new_n583), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n594), .B2(new_n581), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n513), .ZN(new_n596));
  INV_X1    g410(.A(new_n505), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n533), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n534), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT33), .B1(new_n599), .B2(new_n600), .ZN(new_n603));
  OR3_X1    g417(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT97), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n535), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT97), .B1(new_n602), .B2(new_n603), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n537), .A2(G902), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n536), .A2(new_n537), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n597), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n596), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n592), .A2(new_n333), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  INV_X1    g431(.A(new_n539), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n505), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n596), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n592), .A2(new_n333), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G107), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  AOI22_X1  g437(.A1(G472), .A2(new_n588), .B1(new_n450), .B2(new_n456), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n369), .A2(KEYINPUT36), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n365), .B(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(new_n312), .A3(new_n335), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n376), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n333), .A2(new_n585), .A3(new_n624), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT37), .B(G110), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G12));
  NAND2_X1  g445(.A1(new_n453), .A2(new_n459), .ZN(new_n632));
  INV_X1    g446(.A(new_n619), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n512), .A2(G900), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n509), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n595), .A2(new_n628), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n333), .A2(new_n632), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n238), .ZN(G30));
  XNOR2_X1  g454(.A(new_n635), .B(KEYINPUT39), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n333), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT40), .Z(new_n643));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n455), .A2(new_n457), .A3(new_n452), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n439), .A2(new_n440), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n423), .A2(new_n415), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(G472), .B1(new_n649), .B2(G902), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n459), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n376), .A2(new_n627), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n594), .A2(new_n581), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT38), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n597), .A2(new_n618), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n653), .A2(new_n656), .A3(new_n593), .A4(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n658), .B1(new_n643), .B2(new_n644), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n645), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n234), .ZN(G45));
  INV_X1    g475(.A(new_n635), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n637), .A2(new_n613), .A3(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n333), .A2(new_n632), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT99), .B(G146), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G48));
  NAND2_X1  g480(.A1(new_n310), .A2(new_n312), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G469), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(KEYINPUT100), .A3(new_n313), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n670), .A3(G469), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n326), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n460), .A2(new_n614), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT41), .B(G113), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G15));
  NAND3_X1  g489(.A1(new_n460), .A2(new_n620), .A3(new_n672), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G116), .ZN(G18));
  NOR2_X1   g491(.A1(new_n540), .A2(new_n652), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT32), .B1(new_n450), .B2(new_n456), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n427), .A2(new_n431), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(G472), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n646), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n678), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n326), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n313), .A2(KEYINPUT100), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n311), .B1(new_n310), .B2(new_n312), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n671), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n684), .B(new_n595), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT101), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  AOI211_X1 g504(.A(new_n326), .B(new_n584), .C1(new_n669), .C2(new_n671), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n628), .A2(new_n513), .A3(new_n539), .A4(new_n505), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n453), .B2(new_n459), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  AOI22_X1  g511(.A1(new_n588), .A2(G472), .B1(new_n456), .B2(new_n454), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n698), .A2(new_n590), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n596), .A2(new_n657), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n672), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  NAND2_X1  g516(.A1(new_n454), .A2(new_n456), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n589), .A2(new_n628), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n698), .A2(KEYINPUT102), .A3(new_n628), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n613), .A2(new_n662), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n691), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n582), .A2(new_n593), .A3(new_n583), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n320), .B(KEYINPUT103), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n298), .B2(G469), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n326), .B1(new_n313), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n713), .B1(new_n717), .B2(KEYINPUT104), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n719), .B(new_n326), .C1(new_n313), .C2(new_n716), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n712), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n319), .A2(new_n714), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT86), .B1(new_n308), .B2(new_n191), .ZN(new_n723));
  AOI211_X1 g537(.A(new_n305), .B(new_n192), .C1(new_n287), .C2(new_n307), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(G902), .B1(new_n725), .B2(new_n303), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n722), .B1(new_n726), .B2(new_n311), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n719), .B1(new_n727), .B2(new_n326), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n717), .A2(KEYINPUT104), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(KEYINPUT105), .A3(new_n729), .A4(new_n713), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n721), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n590), .B1(new_n679), .B2(new_n682), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n460), .A2(KEYINPUT106), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n731), .A2(new_n709), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n732), .B1(new_n721), .B2(new_n730), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n613), .A2(KEYINPUT42), .A3(new_n662), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n736), .A2(KEYINPUT42), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G131), .ZN(G33));
  INV_X1    g554(.A(new_n636), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NOR2_X1   g557(.A1(new_n298), .A2(KEYINPUT45), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n311), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n298), .A2(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n714), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(KEYINPUT107), .A3(new_n313), .ZN(new_n749));
  INV_X1    g563(.A(new_n747), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n715), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n749), .B1(KEYINPUT46), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT107), .B1(new_n748), .B2(new_n313), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n684), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n641), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n505), .A2(KEYINPUT108), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n505), .A2(KEYINPUT108), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n612), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT43), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n612), .A2(new_n761), .A3(new_n505), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n624), .A3(new_n652), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(KEYINPUT44), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(KEYINPUT44), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n594), .A2(new_n541), .A3(new_n581), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n756), .A2(new_n765), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n196), .ZN(G39));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n754), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(KEYINPUT47), .B(new_n684), .C1(new_n752), .C2(new_n753), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n709), .A2(new_n379), .A3(new_n713), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n632), .A3(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(G140), .Z(G42));
  NOR3_X1   g590(.A1(new_n651), .A2(new_n379), .A3(new_n509), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n669), .A2(new_n671), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n684), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n767), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n597), .A3(new_n612), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n763), .A2(new_n509), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n699), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n782), .B(new_n507), .C1(new_n689), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n783), .A2(new_n780), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n734), .A2(new_n735), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT48), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n785), .A2(new_n786), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n787), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n779), .A2(KEYINPUT116), .A3(new_n541), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n672), .B2(new_n593), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n784), .A2(new_n655), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT50), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n597), .A2(new_n612), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n781), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n804), .A2(new_n805), .B1(new_n788), .B2(new_n708), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(KEYINPUT117), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n801), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n788), .A2(new_n708), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n781), .A2(new_n805), .A3(new_n802), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n801), .A2(new_n809), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n800), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n778), .A2(new_n327), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n771), .A2(new_n772), .A3(new_n813), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n814), .A2(KEYINPUT119), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n784), .A2(new_n767), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(KEYINPUT119), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT51), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n773), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n813), .B(KEYINPUT115), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n816), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n806), .A2(new_n807), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n800), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n794), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT109), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n596), .B2(new_n619), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n633), .A2(new_n595), .A3(KEYINPUT109), .A4(new_n513), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n592), .A2(new_n333), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n629), .A3(new_n615), .A4(new_n586), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n690), .A2(new_n695), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n460), .B(new_n672), .C1(new_n614), .C2(new_n620), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n701), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n835), .A2(new_n739), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n505), .A2(new_n539), .A3(new_n635), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n837), .A2(new_n652), .A3(new_n767), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n632), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n737), .A2(new_n741), .B1(new_n333), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n708), .A2(new_n731), .A3(new_n709), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n840), .A2(KEYINPUT110), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n657), .A2(new_n584), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n635), .B(KEYINPUT111), .Z(new_n848));
  AND2_X1   g662(.A1(new_n717), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n651), .A2(new_n652), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n333), .B(new_n632), .C1(new_n638), .C2(new_n663), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n698), .A2(KEYINPUT102), .A3(new_n628), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT102), .B1(new_n698), .B2(new_n628), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n691), .A2(new_n709), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n850), .B(new_n851), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT52), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n710), .A2(new_n858), .A3(new_n851), .A4(new_n850), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n836), .A2(new_n846), .A3(KEYINPUT53), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n835), .A2(new_n739), .A3(new_n857), .A4(new_n859), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n839), .A2(new_n333), .ZN(new_n864));
  AND4_X1   g678(.A1(KEYINPUT110), .A2(new_n742), .A3(new_n841), .A4(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT110), .B1(new_n840), .B2(new_n841), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n862), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n861), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(KEYINPUT112), .B(new_n862), .C1(new_n863), .C2(new_n867), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(KEYINPUT54), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT113), .B1(new_n832), .B2(new_n834), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT113), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n696), .A2(new_n874), .A3(new_n701), .A4(new_n833), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n739), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n831), .A2(new_n862), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n879), .A2(new_n857), .A3(new_n859), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n873), .A2(new_n739), .A3(KEYINPUT114), .A4(new_n875), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n878), .A2(new_n846), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n882), .A2(new_n868), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n826), .A2(new_n872), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n506), .A2(new_n189), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n328), .A2(new_n541), .ZN(new_n888));
  OR4_X1    g702(.A1(new_n379), .A2(new_n655), .A3(new_n759), .A4(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n778), .B(KEYINPUT49), .Z(new_n890));
  OR3_X1    g704(.A1(new_n889), .A2(new_n890), .A3(new_n651), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n887), .A2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n189), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n312), .B1(new_n882), .B2(new_n868), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(G210), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n556), .A2(new_n570), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT121), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n568), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n894), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n896), .B2(new_n901), .ZN(G51));
  NAND2_X1  g717(.A1(new_n882), .A2(new_n868), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(KEYINPUT122), .A3(new_n884), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n904), .A2(new_n907), .A3(KEYINPUT54), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n714), .B(KEYINPUT57), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n310), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n895), .A2(new_n750), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n893), .B1(new_n911), .B2(new_n912), .ZN(G54));
  NOR2_X1   g727(.A1(new_n484), .A2(new_n496), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(KEYINPUT58), .A2(G475), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT123), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n895), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n915), .B1(new_n895), .B2(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n893), .ZN(G60));
  NAND2_X1  g734(.A1(G478), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT59), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n906), .A2(new_n608), .A3(new_n908), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n894), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n872), .A2(new_n884), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n608), .B1(new_n925), .B2(new_n922), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n926), .ZN(G63));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT60), .Z(new_n929));
  XOR2_X1   g743(.A(new_n626), .B(KEYINPUT124), .Z(new_n930));
  NAND3_X1  g744(.A1(new_n904), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n904), .A2(new_n929), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n894), .B(new_n931), .C1(new_n932), .C2(new_n372), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT61), .B1(new_n931), .B2(KEYINPUT125), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G66));
  XNOR2_X1  g749(.A(new_n835), .B(KEYINPUT126), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n189), .ZN(new_n937));
  OAI21_X1  g751(.A(G953), .B1(new_n510), .B2(new_n563), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n898), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(G898), .B2(new_n189), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n939), .B(new_n941), .ZN(G69));
  AOI21_X1  g756(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n396), .B(new_n487), .Z(new_n944));
  NAND2_X1  g758(.A1(G900), .A2(G953), .ZN(new_n945));
  INV_X1    g759(.A(new_n742), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n710), .A2(new_n851), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n768), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n775), .ZN(new_n949));
  INV_X1    g763(.A(new_n756), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n790), .A3(new_n847), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n948), .A2(new_n739), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n944), .B(new_n945), .C1(new_n952), .C2(G953), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n947), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n645), .B2(new_n659), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n956), .A2(KEYINPUT62), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(KEYINPUT62), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n613), .A2(new_n619), .ZN(new_n959));
  NOR4_X1   g773(.A1(new_n642), .A2(new_n732), .A3(new_n767), .A4(new_n959), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n775), .A2(new_n768), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n944), .B1(new_n962), .B2(new_n189), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n943), .B1(new_n954), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n943), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n962), .A2(new_n189), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n965), .B(new_n953), .C1(new_n966), .C2(new_n944), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(G72));
  XNOR2_X1  g782(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n380), .A2(new_n312), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n962), .B2(new_n936), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n972), .A2(new_n425), .A3(new_n408), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n647), .A2(new_n419), .A3(new_n417), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n870), .A2(new_n871), .A3(new_n971), .A4(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n971), .B1(new_n952), .B2(new_n936), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n408), .A2(new_n425), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n893), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n973), .A2(new_n975), .A3(new_n978), .ZN(G57));
endmodule


