//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067;
  AND2_X1   g000(.A1(KEYINPUT78), .A2(G140), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT78), .A2(G140), .ZN(new_n188));
  OAI21_X1  g002(.A(G125), .B1(new_n187), .B2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT79), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT79), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n194), .B(G125), .C1(new_n187), .C2(new_n188), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n190), .A2(KEYINPUT16), .A3(new_n193), .A4(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(G125), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT16), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT80), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT78), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n191), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT78), .A2(G140), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n192), .B1(new_n206), .B2(new_n194), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n207), .A2(new_n199), .A3(KEYINPUT16), .A4(new_n190), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n201), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT65), .B(G131), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(G237), .A2(G953), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(G143), .A3(G214), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(G143), .B1(new_n213), .B2(G214), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n212), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n216), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(new_n211), .A3(new_n214), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  MUX2_X1   g034(.A(new_n220), .B(new_n217), .S(KEYINPUT17), .Z(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n201), .A2(new_n222), .A3(new_n208), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n210), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n214), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT18), .A2(G131), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n225), .B(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n195), .A2(new_n193), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n204), .A2(new_n205), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n194), .B1(new_n230), .B2(G125), .ZN(new_n231));
  OAI21_X1  g045(.A(G146), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT91), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n193), .A2(new_n197), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G146), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n232), .A2(new_n233), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n233), .B1(new_n232), .B2(new_n240), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n228), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(G113), .B(G122), .ZN(new_n245));
  INV_X1    g059(.A(G104), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n224), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n247), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT19), .B1(new_n229), .B2(new_n231), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT64), .B(G146), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n234), .A2(KEYINPUT19), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n220), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n222), .B1(new_n201), .B2(new_n208), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n222), .B1(new_n207), .B2(new_n190), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT91), .B1(new_n257), .B2(new_n239), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n227), .B1(new_n258), .B2(new_n241), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n249), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n248), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(G475), .A2(G902), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT92), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT20), .ZN(new_n265));
  INV_X1    g079(.A(new_n262), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n248), .B2(new_n260), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT20), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT92), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n262), .A2(KEYINPUT93), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n262), .A2(KEYINPUT93), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT20), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT94), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n261), .A2(KEYINPUT94), .A3(new_n272), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n265), .A2(new_n269), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n224), .A2(new_n244), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n249), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n248), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G475), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G116), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT14), .A3(G122), .ZN(new_n286));
  XOR2_X1   g100(.A(G116), .B(G122), .Z(new_n287));
  OAI211_X1 g101(.A(G107), .B(new_n286), .C1(new_n287), .C2(KEYINPUT14), .ZN(new_n288));
  OR2_X1    g102(.A1(KEYINPUT82), .A2(G107), .ZN(new_n289));
  NAND2_X1  g103(.A1(KEYINPUT82), .A2(G107), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G143), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G128), .ZN(new_n293));
  INV_X1    g107(.A(G128), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G143), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G134), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n296), .A2(new_n297), .ZN(new_n299));
  OAI221_X1 g113(.A(new_n288), .B1(new_n291), .B2(new_n287), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n287), .B(new_n291), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT13), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n293), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n295), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n293), .A2(new_n302), .ZN(new_n305));
  OAI21_X1  g119(.A(G134), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n296), .A2(new_n297), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n301), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT9), .B(G234), .ZN(new_n309));
  INV_X1    g123(.A(G217), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n309), .A2(new_n310), .A3(G953), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n300), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT95), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n300), .A2(new_n308), .ZN(new_n315));
  INV_X1    g129(.A(new_n311), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n300), .A2(new_n308), .A3(KEYINPUT95), .A4(new_n311), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n314), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT76), .B(G902), .Z(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G478), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n322), .A2(KEYINPUT15), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n284), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G221), .B1(new_n309), .B2(G902), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G110), .B(G140), .ZN(new_n329));
  INV_X1    g143(.A(G227), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G953), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n329), .B(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT84), .ZN(new_n333));
  INV_X1    g147(.A(G101), .ZN(new_n334));
  AND2_X1   g148(.A1(KEYINPUT82), .A2(G107), .ZN(new_n335));
  NOR2_X1   g149(.A1(KEYINPUT82), .A2(G107), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n246), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G107), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G104), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n334), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n335), .A2(new_n336), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n338), .B2(G104), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n341), .A2(new_n342), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT83), .B(G101), .Z(new_n346));
  AOI22_X1  g160(.A1(new_n333), .A2(new_n340), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(G104), .B1(new_n289), .B2(new_n290), .ZN(new_n348));
  INV_X1    g162(.A(new_n339), .ZN(new_n349));
  OAI21_X1  g163(.A(G101), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT84), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n235), .A2(new_n237), .A3(G143), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n292), .A2(G146), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n352), .A2(new_n353), .A3(G128), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n222), .A2(G143), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n294), .B1(new_n356), .B2(KEYINPUT1), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n352), .B2(new_n354), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n355), .B1(new_n358), .B2(KEYINPUT85), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n360));
  AOI211_X1 g174(.A(new_n360), .B(new_n357), .C1(new_n352), .C2(new_n354), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n347), .B(new_n351), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n294), .B1(new_n352), .B2(KEYINPUT1), .ZN(new_n363));
  INV_X1    g177(.A(new_n356), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n238), .B2(new_n292), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n333), .B(G101), .C1(new_n348), .C2(new_n349), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n342), .A2(new_n289), .A3(new_n290), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n344), .A2(new_n339), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n346), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n340), .A2(new_n333), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n366), .B(new_n355), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n362), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT11), .B1(new_n297), .B2(G137), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT11), .ZN(new_n376));
  INV_X1    g190(.A(G137), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(G134), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n297), .A2(G137), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n211), .ZN(new_n381));
  INV_X1    g195(.A(G131), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n375), .A2(new_n378), .B1(new_n297), .B2(G137), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n374), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT12), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n374), .A2(KEYINPUT12), .A3(new_n384), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT86), .B(KEYINPUT10), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n362), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n356), .B1(new_n251), .B2(G143), .ZN(new_n392));
  XOR2_X1   g206(.A(KEYINPUT0), .B(G128), .Z(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n352), .A2(KEYINPUT0), .A3(G128), .A4(new_n354), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n334), .B1(new_n368), .B2(new_n369), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n370), .B(KEYINPUT4), .C1(new_n345), .C2(new_n334), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n384), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n371), .A2(new_n372), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n355), .B1(new_n363), .B2(new_n365), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT70), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(KEYINPUT70), .B(new_n355), .C1(new_n363), .C2(new_n365), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n403), .A2(new_n406), .A3(KEYINPUT10), .A4(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n391), .A2(new_n401), .A3(new_n402), .A4(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT87), .B1(new_n389), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT12), .B1(new_n374), .B2(new_n384), .ZN(new_n411));
  AOI211_X1 g225(.A(new_n386), .B(new_n402), .C1(new_n362), .C2(new_n373), .ZN(new_n412));
  OAI211_X1 g226(.A(KEYINPUT87), .B(new_n409), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n332), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n332), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n362), .A2(new_n390), .B1(new_n399), .B2(new_n400), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n402), .B1(new_n418), .B2(new_n408), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n415), .A2(G469), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G469), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(new_n281), .ZN(new_n424));
  INV_X1    g238(.A(new_n320), .ZN(new_n425));
  INV_X1    g239(.A(new_n409), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n332), .B1(new_n419), .B2(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n416), .B(new_n409), .C1(new_n411), .C2(new_n412), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n424), .B1(new_n429), .B2(new_n423), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n328), .B1(new_n422), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G113), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n285), .A2(G119), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT5), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G119), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G116), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n285), .A2(G119), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT5), .ZN(new_n439));
  XNOR2_X1  g253(.A(G116), .B(G119), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n432), .A2(KEYINPUT2), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT2), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G113), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n435), .A2(new_n439), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n351), .A2(new_n370), .A3(new_n367), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n398), .A2(new_n397), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n436), .A2(G116), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n441), .B(new_n443), .C1(new_n433), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n444), .A2(new_n440), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT68), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT68), .B1(new_n449), .B2(new_n450), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n447), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n370), .A2(KEYINPUT4), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(new_n398), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n446), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G110), .B(G122), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n457), .B(new_n446), .C1(new_n453), .C2(new_n455), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT6), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(KEYINPUT6), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n400), .B(new_n447), .C1(new_n452), .C2(new_n451), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n457), .B1(new_n464), .B2(new_n446), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n456), .A2(new_n467), .A3(new_n458), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT88), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n462), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G224), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(G953), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n202), .B(new_n355), .C1(new_n363), .C2(new_n365), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n202), .B1(new_n394), .B2(new_n395), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT89), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n396), .A2(G125), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n478), .B1(new_n479), .B2(new_n474), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n473), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT89), .B1(new_n475), .B2(new_n476), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n478), .A3(new_n474), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n472), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n470), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G210), .B1(G237), .B2(G902), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n475), .A2(new_n476), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n473), .A2(KEYINPUT7), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n457), .B(KEYINPUT8), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n403), .A2(new_n445), .ZN(new_n493));
  INV_X1    g307(.A(new_n446), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n490), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n491), .A2(new_n495), .A3(new_n461), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n281), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n487), .A2(new_n488), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n488), .ZN(new_n501));
  OAI211_X1 g315(.A(KEYINPUT88), .B(new_n468), .C1(new_n463), .C2(new_n465), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n485), .B1(new_n502), .B2(new_n462), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n501), .B1(new_n503), .B2(new_n498), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(KEYINPUT90), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n488), .B1(new_n487), .B2(new_n499), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G953), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n510), .A2(G952), .ZN(new_n511));
  INV_X1    g325(.A(G234), .ZN(new_n512));
  INV_X1    g326(.A(G237), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AOI211_X1 g329(.A(new_n510), .B(new_n320), .C1(G234), .C2(G237), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT21), .B(G898), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G214), .B1(G237), .B2(G902), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AND4_X1   g335(.A1(new_n326), .A2(new_n431), .A3(new_n509), .A4(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT77), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT28), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT66), .B1(new_n377), .B2(G134), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT66), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n297), .A3(G137), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n377), .A2(G134), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(G131), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n381), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n529), .B2(G131), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n406), .A2(new_n534), .A3(new_n407), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n384), .A2(new_n395), .A3(new_n394), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT69), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT69), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n384), .A2(new_n538), .A3(new_n395), .A4(new_n394), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n451), .A2(new_n452), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n535), .A2(new_n541), .A3(new_n537), .A4(new_n539), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n524), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n536), .A2(new_n541), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT28), .B1(new_n546), .B2(new_n535), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n213), .A2(G210), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT27), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT26), .B(G101), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT29), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n545), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n523), .B1(new_n553), .B2(new_n425), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n543), .A2(new_n544), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT28), .ZN(new_n556));
  INV_X1    g370(.A(new_n547), .ZN(new_n557));
  INV_X1    g371(.A(new_n552), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(KEYINPUT77), .A3(new_n320), .ZN(new_n560));
  INV_X1    g374(.A(new_n551), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n540), .A2(KEYINPUT30), .ZN(new_n562));
  INV_X1    g376(.A(new_n404), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n529), .A2(G131), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT67), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n381), .A3(new_n531), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n536), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(KEYINPUT30), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n541), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n544), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n561), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT75), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n567), .A2(new_n542), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n544), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(new_n547), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n572), .A2(new_n573), .B1(new_n551), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n573), .A3(new_n551), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT29), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n554), .B(new_n560), .C1(new_n578), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G472), .ZN(new_n583));
  NOR2_X1   g397(.A1(G472), .A2(G902), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n584), .A2(KEYINPUT32), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n561), .B1(new_n576), .B2(new_n547), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT74), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(KEYINPUT74), .B(new_n561), .C1(new_n576), .C2(new_n547), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n544), .A2(new_n551), .ZN(new_n591));
  OAI211_X1 g405(.A(KEYINPUT71), .B(KEYINPUT31), .C1(new_n570), .C2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n591), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n568), .B1(KEYINPUT30), .B2(new_n540), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n594), .B1(new_n595), .B2(new_n541), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT71), .B1(new_n596), .B2(KEYINPUT31), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n590), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n562), .A2(new_n569), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n591), .B1(new_n599), .B2(new_n542), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT72), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT31), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n594), .B(new_n602), .C1(new_n595), .C2(new_n541), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT72), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n585), .B1(new_n598), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n584), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT71), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n600), .B2(new_n602), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n610), .A2(new_n592), .B1(new_n588), .B2(new_n589), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n603), .A2(new_n605), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n583), .B(new_n607), .C1(new_n613), .C2(KEYINPUT32), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT24), .B(G110), .Z(new_n615));
  XNOR2_X1  g429(.A(G119), .B(G128), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT23), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n436), .B2(G128), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n294), .A2(KEYINPUT23), .A3(G119), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n619), .B(new_n620), .C1(G119), .C2(new_n294), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G110), .ZN(new_n622));
  INV_X1    g436(.A(new_n223), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n617), .B(new_n622), .C1(new_n623), .C2(new_n255), .ZN(new_n624));
  OAI22_X1  g438(.A1(new_n621), .A2(G110), .B1(new_n616), .B2(new_n615), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n240), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n255), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT22), .B(G137), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n510), .A2(G221), .A3(G234), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n629), .B(new_n630), .Z(new_n631));
  NAND3_X1  g445(.A1(new_n624), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n631), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n622), .A2(new_n617), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n210), .B2(new_n223), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n635), .B2(new_n627), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n632), .A2(new_n636), .A3(new_n320), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT81), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT25), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n310), .B1(new_n320), .B2(G234), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n637), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n632), .A2(new_n636), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n641), .A2(G902), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n522), .A2(new_n614), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(new_n346), .Z(G3));
  INV_X1    g464(.A(G472), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n610), .A2(new_n592), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n612), .A3(new_n590), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n651), .B1(new_n653), .B2(new_n320), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n654), .A2(new_n613), .A3(new_n647), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT33), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n315), .B2(new_n316), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n319), .A2(new_n656), .B1(new_n312), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n425), .A2(new_n322), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n658), .A2(new_n659), .B1(new_n322), .B2(new_n321), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n277), .B2(new_n283), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n520), .B1(new_n500), .B2(new_n504), .ZN(new_n663));
  INV_X1    g477(.A(new_n518), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n655), .A2(new_n431), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  OAI211_X1 g483(.A(new_n265), .B(new_n269), .C1(KEYINPUT20), .C2(new_n263), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n325), .A3(new_n283), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n655), .A2(new_n431), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n338), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NOR2_X1   g490(.A1(new_n654), .A2(new_n613), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT97), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n624), .A2(new_n678), .A3(new_n628), .ZN(new_n679));
  OAI21_X1  g493(.A(KEYINPUT97), .B1(new_n635), .B2(new_n627), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n633), .A2(KEYINPUT36), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n681), .B1(new_n679), .B2(new_n680), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n645), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT98), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT98), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n686), .B(new_n645), .C1(new_n682), .C2(new_n683), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n643), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n522), .A2(new_n677), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  XNOR2_X1  g505(.A(KEYINPUT99), .B(G900), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n515), .B1(new_n516), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n671), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT87), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n416), .B1(new_n697), .B2(new_n413), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n423), .A3(new_n420), .ZN(new_n699));
  INV_X1    g513(.A(new_n428), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n391), .A2(new_n401), .A3(new_n408), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n384), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n416), .B1(new_n702), .B2(new_n409), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n423), .B(new_n320), .C1(new_n700), .C2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n424), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n327), .B(new_n663), .C1(new_n699), .C2(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n643), .A2(new_n685), .A3(new_n687), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n614), .A2(new_n694), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G128), .ZN(G30));
  NAND2_X1  g525(.A1(new_n505), .A2(new_n508), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT38), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n284), .A2(new_n325), .A3(new_n519), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n713), .A2(new_n688), .A3(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n693), .B(KEYINPUT39), .Z(new_n716));
  NAND2_X1  g530(.A1(new_n431), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n570), .A2(new_n571), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n561), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n281), .B1(new_n555), .B2(new_n551), .ZN(new_n722));
  OAI21_X1  g536(.A(G472), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n607), .B(new_n723), .C1(new_n613), .C2(KEYINPUT32), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n715), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(new_n725), .B(KEYINPUT101), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  NOR2_X1   g541(.A1(new_n662), .A2(new_n693), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n614), .A2(new_n709), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  OAI21_X1  g544(.A(new_n320), .B1(new_n700), .B2(new_n703), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G469), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n327), .A3(new_n704), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT102), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT102), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n732), .A2(new_n735), .A3(new_n327), .A4(new_n704), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n614), .A2(new_n737), .A3(new_n648), .A4(new_n666), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G15));
  NAND4_X1  g554(.A1(new_n614), .A2(new_n737), .A3(new_n648), .A4(new_n672), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  AND3_X1   g556(.A1(new_n732), .A2(new_n327), .A3(new_n704), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n663), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(new_n708), .A3(new_n518), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n614), .A3(new_n326), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  AOI21_X1  g561(.A(new_n551), .B1(new_n556), .B2(new_n557), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(KEYINPUT31), .B2(new_n596), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n608), .B1(new_n749), .B2(new_n612), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n654), .A2(new_n647), .A3(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n734), .A2(new_n664), .A3(new_n736), .ZN(new_n752));
  INV_X1    g566(.A(new_n283), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n264), .B1(new_n263), .B2(KEYINPUT20), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n267), .A2(KEYINPUT92), .A3(new_n268), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n275), .A2(new_n276), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n503), .A2(new_n501), .A3(new_n498), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n325), .B(new_n519), .C1(new_n506), .C2(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT103), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n324), .B(new_n520), .C1(new_n500), .C2(new_n504), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT103), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n284), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n751), .A2(new_n752), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT104), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT104), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n751), .A2(new_n752), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G122), .ZN(G24));
  NOR2_X1   g585(.A1(new_n654), .A2(new_n750), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n743), .A2(new_n688), .A3(new_n663), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n728), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G125), .ZN(G27));
  NAND2_X1  g589(.A1(new_n712), .A2(new_n519), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n327), .B1(new_n699), .B2(new_n706), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n614), .A2(new_n778), .A3(new_n648), .A4(new_n728), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT105), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n382), .ZN(G33));
  AND4_X1   g599(.A1(new_n614), .A2(new_n778), .A3(new_n648), .A4(new_n694), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n297), .ZN(G36));
  OR3_X1    g601(.A1(new_n284), .A2(KEYINPUT43), .A3(new_n660), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT43), .B1(new_n284), .B2(new_n660), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT107), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n688), .B1(new_n654), .B2(new_n613), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT108), .B1(new_n794), .B2(KEYINPUT44), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT44), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n796), .B(new_n797), .C1(new_n792), .C2(new_n793), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n794), .A2(KEYINPUT44), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n415), .A2(new_n421), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n423), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n415), .A2(KEYINPUT45), .A3(new_n421), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n705), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT46), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT106), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n805), .A2(KEYINPUT46), .A3(new_n705), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(new_n704), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n806), .A2(KEYINPUT106), .A3(new_n807), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n814), .A2(new_n327), .ZN(new_n815));
  INV_X1    g629(.A(new_n776), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n800), .A2(new_n716), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n799), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(new_n377), .ZN(G39));
  NAND2_X1  g633(.A1(new_n814), .A2(new_n327), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT47), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n814), .A2(KEYINPUT47), .A3(new_n327), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n728), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n825), .A2(new_n614), .A3(new_n648), .A4(new_n776), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n829));
  NOR2_X1   g643(.A1(G952), .A2(G953), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n328), .B(new_n693), .C1(new_n422), .C2(new_n430), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n607), .A2(new_n723), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT32), .B1(new_n653), .B2(new_n584), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n708), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n758), .A2(new_n760), .A3(KEYINPUT103), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n763), .B1(new_n762), .B2(new_n284), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n832), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n777), .A2(new_n688), .A3(new_n693), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n765), .A2(new_n841), .A3(new_n724), .A4(KEYINPUT110), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n710), .A2(new_n729), .A3(new_n774), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT52), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n710), .A2(new_n774), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT52), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n779), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT42), .B1(new_n779), .B2(KEYINPUT105), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n852), .A2(new_n853), .A3(new_n786), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n284), .A2(new_n324), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT109), .B1(new_n855), .B2(new_n661), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n661), .A2(KEYINPUT109), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n431), .A2(new_n509), .A3(new_n521), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n655), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n738), .A3(new_n741), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n746), .A2(new_n649), .A3(new_n689), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n778), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n708), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n670), .A2(new_n283), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n866), .A2(new_n325), .A3(new_n693), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n614), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n772), .A2(new_n728), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n854), .A2(new_n770), .A3(new_n863), .A4(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n831), .B1(new_n851), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n847), .B1(new_n843), .B2(new_n844), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT111), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT111), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n846), .A2(new_n876), .A3(new_n848), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n860), .A2(new_n738), .A3(new_n741), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n746), .A2(new_n649), .A3(new_n689), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n770), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n786), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n782), .A2(new_n783), .A3(new_n870), .A4(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n875), .A2(new_n877), .A3(new_n883), .A4(KEYINPUT53), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n872), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n875), .A2(new_n877), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n831), .ZN(new_n888));
  XNOR2_X1  g702(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n873), .A2(new_n874), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n883), .A2(new_n890), .A3(KEYINPUT53), .A4(new_n850), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n724), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n776), .A2(new_n733), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(new_n648), .A3(new_n515), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n788), .A2(new_n515), .A3(new_n789), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n751), .ZN(new_n899));
  OAI221_X1 g713(.A(new_n511), .B1(new_n896), .B2(new_n662), .C1(new_n899), .C2(new_n744), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n897), .A2(new_n733), .A3(new_n776), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n614), .A2(new_n648), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g718(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n900), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n898), .A2(new_n751), .A3(new_n816), .ZN(new_n909));
  INV_X1    g723(.A(new_n823), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT47), .B1(new_n814), .B2(new_n327), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n732), .A2(new_n704), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n328), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n909), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT115), .ZN(new_n916));
  INV_X1    g730(.A(new_n660), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n284), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n916), .B1(new_n896), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n724), .A2(new_n647), .A3(new_n514), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n921), .A2(KEYINPUT115), .A3(new_n895), .A4(new_n918), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n901), .A2(new_n688), .A3(new_n772), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n713), .A2(new_n520), .A3(new_n743), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT114), .B1(new_n899), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT50), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(KEYINPUT114), .B(KEYINPUT50), .C1(new_n899), .C2(new_n926), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n925), .A2(KEYINPUT51), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n908), .B1(new_n915), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT116), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT51), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n914), .B(KEYINPUT113), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n909), .B1(new_n912), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n929), .A2(new_n930), .A3(new_n923), .A4(new_n924), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n933), .B(new_n934), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n822), .A2(new_n823), .A3(new_n935), .ZN(new_n939));
  INV_X1    g753(.A(new_n909), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT116), .B1(new_n941), .B2(KEYINPUT51), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n932), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n830), .B1(new_n893), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT49), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n328), .B(new_n520), .C1(new_n913), .C2(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n946), .B(new_n648), .C1(new_n945), .C2(new_n913), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n947), .A2(new_n284), .A3(new_n660), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n894), .A3(new_n713), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n829), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n943), .A2(new_n886), .A3(new_n892), .ZN(new_n952));
  INV_X1    g766(.A(new_n830), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(KEYINPUT118), .A3(new_n949), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n951), .A2(new_n955), .ZN(G75));
  AOI21_X1  g770(.A(new_n320), .B1(new_n888), .B2(new_n891), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n501), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT56), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n470), .B(new_n486), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT55), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n960), .A2(new_n962), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n510), .A2(G952), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(G51));
  XNOR2_X1  g780(.A(new_n424), .B(KEYINPUT57), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n889), .B1(new_n888), .B2(new_n891), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT119), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n892), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI211_X1 g784(.A(KEYINPUT119), .B(new_n889), .C1(new_n888), .C2(new_n891), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n427), .A2(new_n428), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n320), .B(new_n805), .C1(new_n888), .C2(new_n891), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT120), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n965), .B1(new_n974), .B2(new_n976), .ZN(G54));
  INV_X1    g791(.A(new_n965), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n957), .A2(KEYINPUT58), .A3(G475), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n261), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n261), .B2(new_n979), .ZN(G60));
  NAND2_X1  g795(.A1(G478), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT59), .Z(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n886), .B2(new_n892), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n978), .B1(new_n984), .B2(new_n658), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n970), .A2(new_n971), .ZN(new_n986));
  INV_X1    g800(.A(new_n983), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n658), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n985), .B1(new_n986), .B2(new_n988), .ZN(G63));
  NAND2_X1  g803(.A1(new_n888), .A2(new_n891), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n682), .A2(new_n683), .ZN(new_n991));
  NAND2_X1  g805(.A1(G217), .A2(G902), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT60), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n990), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(KEYINPUT61), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n993), .B1(new_n888), .B2(new_n891), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n978), .B1(new_n997), .B2(new_n644), .ZN(new_n998));
  OAI21_X1  g812(.A(KEYINPUT122), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n990), .A2(new_n994), .ZN(new_n1000));
  INV_X1    g814(.A(new_n644), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT61), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(new_n997), .B2(new_n991), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT122), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .A4(new_n978), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n995), .A2(KEYINPUT121), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT121), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n997), .A2(new_n1009), .A3(new_n991), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1008), .A2(new_n1002), .A3(new_n978), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n1003), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1007), .A2(new_n1012), .ZN(G66));
  NAND2_X1  g827(.A1(new_n880), .A2(new_n510), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT123), .Z(new_n1015));
  OAI21_X1  g829(.A(G953), .B1(new_n517), .B2(new_n471), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n502), .B(new_n462), .C1(G898), .C2(new_n510), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1017), .B(new_n1018), .ZN(G69));
  NAND4_X1  g833(.A1(new_n903), .A2(new_n716), .A3(new_n778), .A4(new_n858), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n844), .B(KEYINPUT124), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n726), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT62), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(KEYINPUT62), .B1(new_n726), .B2(new_n1021), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1020), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n827), .B1(new_n799), .B2(new_n817), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n510), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n250), .A2(new_n252), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n599), .B(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n510), .A2(G900), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(new_n330), .B2(G953), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1033), .B(KEYINPUT125), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n902), .A2(new_n839), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n815), .A2(new_n716), .A3(new_n1036), .ZN(new_n1037));
  AND2_X1   g851(.A1(new_n1037), .A2(KEYINPUT126), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1037), .A2(KEYINPUT126), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n854), .B(new_n1021), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n510), .B1(new_n1040), .B2(new_n1027), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1032), .ZN(new_n1042));
  AND2_X1   g856(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n1031), .B(new_n1035), .C1(new_n1043), .C2(new_n1030), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1030), .ZN(new_n1045));
  XNOR2_X1  g859(.A(new_n1022), .B(new_n1023), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1027), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1046), .A2(new_n1047), .A3(new_n1020), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1045), .B1(new_n1048), .B2(new_n510), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1030), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1034), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AND2_X1   g865(.A1(new_n1044), .A2(new_n1051), .ZN(G72));
  NOR3_X1   g866(.A1(new_n1040), .A2(new_n880), .A3(new_n1027), .ZN(new_n1053));
  NAND2_X1  g867(.A1(G472), .A2(G902), .ZN(new_n1054));
  XOR2_X1   g868(.A(new_n1054), .B(KEYINPUT63), .Z(new_n1055));
  INV_X1    g869(.A(new_n1055), .ZN(new_n1056));
  OAI211_X1 g870(.A(new_n561), .B(new_n720), .C1(new_n1053), .C2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g871(.A(new_n1056), .B1(new_n572), .B2(new_n596), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n965), .B1(new_n885), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g874(.A(new_n880), .ZN(new_n1061));
  NAND4_X1  g875(.A1(new_n1046), .A2(new_n1047), .A3(new_n1061), .A4(new_n1020), .ZN(new_n1062));
  INV_X1    g876(.A(KEYINPUT127), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n1062), .A2(new_n1063), .A3(new_n1055), .ZN(new_n1064));
  AND2_X1   g878(.A1(new_n1064), .A2(new_n721), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1062), .A2(new_n1055), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1066), .A2(KEYINPUT127), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n1060), .B1(new_n1065), .B2(new_n1067), .ZN(G57));
endmodule


