//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n469), .A2(G137), .A3(new_n461), .ZN(new_n470));
  INV_X1    g045(.A(G101), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT67), .B1(new_n462), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n461), .A3(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NOR3_X1   g050(.A1(new_n468), .A2(new_n470), .A3(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n469), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n469), .A2(new_n461), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n463), .A2(new_n465), .A3(G126), .A4(G2105), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n461), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(new_n495), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n498), .A2(new_n469), .A3(G138), .A4(new_n461), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n486), .A2(KEYINPUT68), .A3(new_n490), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n493), .A2(new_n496), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT70), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n499), .A2(new_n496), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n503), .A2(new_n504), .A3(new_n493), .A4(new_n500), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT71), .B1(new_n507), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n514), .A2(new_n518), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n517), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n522), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(new_n519), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n516), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n520), .A2(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n522), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n516), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n520), .A2(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n522), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  XNOR2_X1  g129(.A(KEYINPUT73), .B(G65), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n514), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G78), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(new_n510), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT74), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n556), .B(new_n560), .C1(new_n557), .C2(new_n510), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(G651), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n522), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G91), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n520), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n562), .A2(new_n564), .A3(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  NAND2_X1  g143(.A1(new_n563), .A2(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n520), .A2(G49), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND4_X1  g147(.A1(new_n512), .A2(G86), .A3(new_n513), .A4(new_n518), .ZN(new_n573));
  INV_X1    g148(.A(G48), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n574), .B2(new_n519), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n512), .A2(G61), .A3(new_n513), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT75), .Z(new_n578));
  AOI21_X1  g153(.A(new_n516), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n516), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n520), .A2(G47), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n522), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n520), .A2(G54), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT76), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n514), .B2(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n590), .B1(new_n593), .B2(new_n516), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(KEYINPUT77), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(KEYINPUT77), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n522), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n563), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n596), .A2(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n589), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n589), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G280));
  XOR2_X1   g182(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  OAI21_X1  g185(.A(KEYINPUT79), .B1(new_n548), .B2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n609), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  MUX2_X1   g188(.A(KEYINPUT79), .B(new_n611), .S(new_n613), .Z(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n480), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n478), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n461), .A2(G111), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT83), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n616), .B(new_n617), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT84), .B(G2096), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n472), .A2(new_n474), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(new_n469), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT82), .B(G2100), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n623), .A2(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT15), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2435), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(G2435), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2443), .B(G2446), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n642), .A2(new_n644), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n634), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n649), .A2(new_n645), .A3(new_n633), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n648), .A2(new_n650), .A3(G14), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT85), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  OAI21_X1  g234(.A(KEYINPUT17), .B1(new_n654), .B2(new_n657), .ZN(new_n660));
  AOI22_X1  g235(.A1(new_n660), .A2(new_n655), .B1(new_n654), .B2(new_n657), .ZN(new_n661));
  OAI211_X1 g236(.A(KEYINPUT17), .B(new_n656), .C1(new_n654), .C2(new_n657), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT86), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT87), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n669), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(KEYINPUT88), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n669), .A2(new_n672), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n677), .A2(new_n671), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT20), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT89), .B(KEYINPUT90), .Z(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n682), .B(new_n687), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G6), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n580), .B2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT32), .ZN(new_n693));
  INV_X1    g268(.A(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(G16), .A2(G22), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G166), .B2(G16), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(G1971), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(G1971), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n690), .A2(G23), .ZN(new_n700));
  INV_X1    g275(.A(G288), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n690), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT92), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n695), .A2(new_n698), .A3(new_n699), .A4(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT34), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n690), .A2(G24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n587), .B2(new_n690), .ZN(new_n709));
  INV_X1    g284(.A(G1986), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n478), .A2(G119), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n480), .A2(G131), .ZN(new_n713));
  OR2_X1    g288(.A1(G95), .A2(G2105), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n714), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G25), .B(new_n718), .S(G29), .Z(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT35), .B(G1991), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n719), .B(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n707), .A2(new_n711), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT36), .Z(new_n724));
  NOR2_X1   g299(.A1(G29), .A2(G35), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G162), .B2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2090), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT94), .B(G2067), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(G26), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n478), .A2(G128), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n480), .A2(G140), .ZN(new_n734));
  OR2_X1    g309(.A1(G104), .A2(G2105), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n735), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n732), .B1(new_n737), .B2(G29), .ZN(new_n738));
  MUX2_X1   g313(.A(new_n732), .B(new_n738), .S(KEYINPUT28), .Z(new_n739));
  AOI21_X1  g314(.A(new_n728), .B1(new_n730), .B2(new_n739), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n478), .A2(G129), .B1(G105), .B2(new_n624), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n480), .A2(G141), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT26), .Z(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G29), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G29), .B2(G32), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n739), .A2(new_n730), .ZN(new_n751));
  OR2_X1    g326(.A1(G29), .A2(G33), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(new_n461), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT95), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n480), .A2(G139), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT25), .Z(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n752), .B1(new_n759), .B2(new_n731), .ZN(new_n760));
  INV_X1    g335(.A(G2072), .ZN(new_n761));
  OR2_X1    g336(.A1(KEYINPUT24), .A2(G34), .ZN(new_n762));
  NAND2_X1  g337(.A1(KEYINPUT24), .A2(G34), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n762), .A2(new_n731), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G160), .B2(new_n731), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n760), .A2(new_n761), .B1(G2084), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n740), .A2(new_n750), .A3(new_n751), .A4(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n760), .A2(new_n761), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n748), .A2(new_n749), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT96), .ZN(new_n771));
  NOR2_X1   g346(.A1(G27), .A2(G29), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G164), .B2(G29), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2078), .ZN(new_n774));
  NOR4_X1   g349(.A1(new_n767), .A2(new_n769), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(KEYINPUT93), .B1(new_n776), .B2(G16), .ZN(new_n777));
  OR3_X1    g352(.A1(new_n776), .A2(KEYINPUT93), .A3(G16), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n777), .B(new_n778), .C1(new_n548), .C2(new_n690), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G1341), .Z(new_n780));
  XOR2_X1   g355(.A(KEYINPUT31), .B(G11), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT97), .B(G28), .ZN(new_n782));
  NOR2_X1   g357(.A1(KEYINPUT98), .A2(KEYINPUT30), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(G29), .B1(KEYINPUT98), .B2(KEYINPUT30), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G5), .A2(G16), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G171), .B2(G16), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n786), .B1(new_n788), .B2(G1961), .ZN(new_n789));
  NAND2_X1  g364(.A1(G168), .A2(G16), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G16), .B2(G21), .ZN(new_n791));
  INV_X1    g366(.A(G1966), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n602), .A2(G16), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G4), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1348), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n791), .A2(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n789), .B(new_n796), .C1(new_n795), .C2(new_n794), .ZN(new_n797));
  NAND2_X1  g372(.A1(G299), .A2(G16), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n690), .A2(KEYINPUT23), .A3(G20), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT23), .ZN(new_n800));
  INV_X1    g375(.A(G20), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(G16), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n798), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1956), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G1961), .B2(new_n788), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n775), .A2(new_n780), .A3(new_n797), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n724), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n765), .A2(G2084), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n621), .A2(new_n731), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n791), .A2(new_n792), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n807), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(G150));
  INV_X1    g387(.A(G150), .ZN(G311));
  AOI22_X1  g388(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(new_n516), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n520), .A2(G55), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n522), .B2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT101), .B(G860), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT37), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n602), .A2(G559), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n819), .A2(new_n548), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n815), .A2(new_n818), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n544), .B2(new_n547), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n825), .B(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n822), .B1(new_n832), .B2(new_n820), .ZN(G145));
  XNOR2_X1  g408(.A(new_n718), .B(new_n627), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n478), .A2(G130), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n480), .A2(G142), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n461), .A2(G118), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT102), .Z(new_n839));
  OAI211_X1 g414(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n834), .B(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n841), .A2(KEYINPUT103), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(KEYINPUT103), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n759), .B(new_n737), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n499), .A2(new_n496), .A3(new_n486), .A4(new_n490), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n745), .B(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n845), .B(new_n847), .Z(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n848), .B1(new_n842), .B2(new_n843), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n484), .B(G160), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n621), .ZN(new_n854));
  AOI21_X1  g429(.A(G37), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n849), .A2(new_n841), .ZN(new_n856));
  INV_X1    g431(.A(new_n854), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n851), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g435(.A(new_n829), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n612), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n602), .B(G299), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(KEYINPUT104), .B1(new_n602), .B2(G299), .ZN(new_n867));
  INV_X1    g442(.A(new_n863), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(KEYINPUT104), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n866), .B1(new_n869), .B2(new_n865), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n864), .B1(new_n870), .B2(new_n862), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT42), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n873), .B(new_n864), .C1(new_n870), .C2(new_n862), .ZN(new_n874));
  XNOR2_X1  g449(.A(G303), .B(G288), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n875), .A2(new_n580), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n580), .ZN(new_n877));
  OR3_X1    g452(.A1(new_n876), .A2(new_n877), .A3(G290), .ZN(new_n878));
  OAI21_X1  g453(.A(G290), .B1(new_n876), .B2(new_n877), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n872), .A2(new_n874), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n872), .B2(new_n874), .ZN(new_n883));
  OAI21_X1  g458(.A(G868), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n819), .A2(new_n605), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n884), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(G295));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n886), .ZN(G331));
  NAND2_X1  g465(.A1(new_n869), .A2(new_n865), .ZN(new_n891));
  INV_X1    g466(.A(new_n866), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n861), .A2(G301), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n829), .A2(G171), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(G286), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(G168), .A3(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n891), .A2(new_n892), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n868), .A3(new_n897), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G37), .B1(new_n901), .B2(new_n881), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n880), .A3(new_n900), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT43), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n880), .B1(new_n899), .B2(new_n900), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n865), .B1(new_n896), .B2(new_n897), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n906), .A2(new_n869), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n880), .B1(new_n906), .B2(new_n863), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n910));
  NOR4_X1   g485(.A1(new_n905), .A2(new_n909), .A3(new_n910), .A4(G37), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT44), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n902), .B2(new_n903), .ZN(new_n913));
  NOR4_X1   g488(.A1(new_n905), .A2(new_n909), .A3(KEYINPUT43), .A4(G37), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n912), .B1(new_n915), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g491(.A(G1384), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n846), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n470), .A2(new_n475), .ZN(new_n921));
  INV_X1    g496(.A(new_n468), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(G40), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n737), .B(G2067), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT107), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n927), .B2(new_n746), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT124), .ZN(new_n929));
  INV_X1    g504(.A(G1996), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT46), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n933), .B(KEYINPUT47), .Z(new_n934));
  XNOR2_X1  g509(.A(new_n745), .B(new_n930), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n718), .A2(new_n720), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n737), .A2(G2067), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n925), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n718), .B(new_n721), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n925), .B1(new_n936), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n587), .A2(new_n710), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n925), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT48), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n934), .A2(new_n940), .A3(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(KEYINPUT109), .B(G8), .C1(new_n923), .C2(new_n918), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(G160), .A2(G40), .A3(new_n846), .A4(new_n917), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT109), .B1(new_n950), .B2(G8), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1976), .ZN(new_n953));
  NOR2_X1   g528(.A1(G288), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT52), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT52), .B1(G288), .B2(new_n953), .ZN(new_n956));
  OAI221_X1 g531(.A(new_n956), .B1(new_n953), .B2(G288), .C1(new_n949), .C2(new_n951), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n580), .A2(new_n694), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT49), .ZN(new_n959));
  OAI21_X1  g534(.A(G1981), .B1(new_n575), .B2(new_n579), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n961), .A2(new_n962), .B1(new_n949), .B2(new_n951), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n955), .A2(new_n957), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(G303), .A2(G8), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G8), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n502), .A2(new_n917), .A3(new_n505), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n923), .B1(new_n971), .B2(new_n919), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n846), .A2(KEYINPUT45), .A3(new_n917), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT108), .B(G1971), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n923), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n918), .B2(KEYINPUT50), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n971), .B2(KEYINPUT50), .ZN(new_n980));
  INV_X1    g555(.A(G2090), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n970), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n964), .A2(new_n969), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n963), .A2(new_n953), .A3(new_n701), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n985), .A2(KEYINPUT110), .A3(new_n958), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT110), .B1(new_n985), .B2(new_n958), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n986), .A2(new_n987), .A3(new_n952), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT63), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n975), .B1(new_n972), .B2(new_n973), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n502), .A2(new_n991), .A3(new_n505), .A4(new_n917), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n923), .B1(new_n918), .B2(KEYINPUT50), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(G2090), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n990), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n969), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n982), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n969), .B(G8), .C1(new_n999), .C2(new_n990), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n964), .A3(new_n1000), .ZN(new_n1001));
  AOI211_X1 g576(.A(G2084), .B(new_n979), .C1(new_n971), .C2(KEYINPUT50), .ZN(new_n1002));
  OR3_X1    g577(.A1(new_n971), .A2(KEYINPUT111), .A3(new_n919), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n923), .B1(new_n918), .B2(new_n919), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT111), .B1(new_n971), .B2(new_n919), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1002), .B1(new_n1006), .B2(new_n792), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G168), .A2(G8), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n989), .B1(new_n1001), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n997), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n989), .B1(new_n1012), .B2(new_n983), .ZN(new_n1013));
  OAI21_X1  g588(.A(G8), .B1(new_n999), .B2(new_n990), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(new_n1011), .A3(new_n997), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1013), .A2(new_n1015), .A3(new_n964), .A4(new_n1016), .ZN(new_n1017));
  AOI211_X1 g592(.A(new_n984), .B(new_n988), .C1(new_n1010), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n971), .A2(new_n919), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT56), .B(G2072), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1019), .A2(new_n978), .A3(new_n1020), .A4(new_n973), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n972), .A2(KEYINPUT115), .A3(new_n1020), .A4(new_n973), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n1026));
  XNOR2_X1  g601(.A(G299), .B(new_n1026), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT113), .B(G1956), .Z(new_n1028));
  NAND2_X1  g603(.A1(new_n994), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT114), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n994), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1025), .A2(new_n1027), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1027), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(KEYINPUT61), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1023), .A2(new_n1024), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT61), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n1027), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n950), .A2(G2067), .ZN(new_n1041));
  OAI211_X1 g616(.A(KEYINPUT60), .B(new_n1041), .C1(new_n980), .C2(G1348), .ZN(new_n1042));
  INV_X1    g617(.A(new_n602), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1042), .A2(KEYINPUT119), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n1042), .B2(KEYINPUT119), .ZN(new_n1045));
  OAI22_X1  g620(.A1(new_n1044), .A2(new_n1045), .B1(KEYINPUT119), .B2(new_n1042), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1041), .B1(new_n980), .B2(G1348), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT117), .B(G1996), .ZN(new_n1050));
  INV_X1    g625(.A(new_n950), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT58), .B(G1341), .ZN(new_n1052));
  OAI22_X1  g627(.A1(new_n974), .A2(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n548), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT59), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1053), .A2(new_n1054), .A3(new_n1057), .A4(new_n548), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1046), .A2(new_n1049), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1035), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT116), .B1(new_n1037), .B2(new_n1027), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1047), .A2(new_n602), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1040), .A2(new_n1059), .B1(new_n1034), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1001), .A2(KEYINPUT121), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n998), .A2(new_n964), .A3(new_n1000), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT51), .B1(new_n1007), .B2(G168), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n970), .B1(new_n1007), .B2(G168), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI211_X1 g647(.A(G286), .B(new_n1002), .C1(new_n1006), .C2(new_n792), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT51), .B1(new_n1073), .B2(new_n970), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n980), .A2(G1961), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n1077));
  INV_X1    g652(.A(G2078), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n972), .A2(new_n1078), .A3(new_n973), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1076), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1004), .A2(KEYINPUT53), .A3(new_n1078), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1003), .A2(new_n1081), .A3(new_n1005), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(G301), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n973), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1086), .A2(new_n1080), .ZN(new_n1087));
  OAI211_X1 g662(.A(KEYINPUT54), .B(new_n1083), .C1(new_n1087), .C2(G301), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1086), .A2(G301), .A3(new_n1080), .ZN(new_n1090));
  AOI21_X1  g665(.A(G301), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1069), .A2(new_n1075), .A3(new_n1088), .A4(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1018), .B1(new_n1065), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1018), .B(KEYINPUT122), .C1(new_n1065), .C2(new_n1093), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1075), .A2(KEYINPUT62), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1075), .A2(KEYINPUT62), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1098), .A2(new_n1069), .A3(new_n1091), .A4(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n943), .A2(KEYINPUT106), .ZN(new_n1103));
  NAND2_X1  g678(.A1(G290), .A2(G1986), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1103), .B(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n942), .B1(new_n924), .B2(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1101), .A2(new_n1102), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1102), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n947), .B1(new_n1107), .B2(new_n1108), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g684(.A1(G227), .A2(new_n459), .ZN(new_n1111));
  NAND2_X1  g685(.A1(new_n651), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g686(.A1(new_n1112), .A2(KEYINPUT125), .ZN(new_n1113));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n1114));
  NAND3_X1  g688(.A1(new_n651), .A2(new_n1114), .A3(new_n1111), .ZN(new_n1115));
  AOI22_X1  g689(.A1(new_n855), .A2(new_n858), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g690(.A(new_n688), .B(new_n1116), .C1(new_n913), .C2(new_n914), .ZN(new_n1117));
  XNOR2_X1  g691(.A(new_n1117), .B(KEYINPUT126), .ZN(G308));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n1119));
  XNOR2_X1  g693(.A(new_n1117), .B(new_n1119), .ZN(G225));
endmodule


