

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U557 ( .A1(n759), .A2(n757), .ZN(n704) );
  XNOR2_X1 U558 ( .A(n737), .B(KEYINPUT32), .ZN(n743) );
  OR2_X1 U559 ( .A1(n742), .A2(n741), .ZN(n523) );
  INV_X1 U560 ( .A(KEYINPUT96), .ZN(n695) );
  XNOR2_X1 U561 ( .A(n696), .B(n695), .ZN(n697) );
  AND2_X1 U562 ( .A1(n743), .A2(n523), .ZN(n783) );
  INV_X1 U563 ( .A(KEYINPUT71), .ZN(n588) );
  INV_X1 U564 ( .A(G651), .ZN(n540) );
  XOR2_X1 U565 ( .A(KEYINPUT15), .B(n592), .Z(n969) );
  NOR2_X1 U566 ( .A1(n620), .A2(n540), .ZN(n636) );
  NOR2_X2 U567 ( .A1(n535), .A2(n534), .ZN(G160) );
  INV_X1 U568 ( .A(G2104), .ZN(n529) );
  NOR2_X4 U569 ( .A1(G2105), .A2(n529), .ZN(n875) );
  NAND2_X1 U570 ( .A1(G101), .A2(n875), .ZN(n524) );
  XNOR2_X1 U571 ( .A(KEYINPUT64), .B(n524), .ZN(n526) );
  INV_X1 U572 ( .A(KEYINPUT23), .ZN(n525) );
  XNOR2_X1 U573 ( .A(n526), .B(n525), .ZN(n528) );
  AND2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n878) );
  NAND2_X1 U575 ( .A1(G113), .A2(n878), .ZN(n527) );
  NAND2_X1 U576 ( .A1(n528), .A2(n527), .ZN(n535) );
  AND2_X1 U577 ( .A1(n529), .A2(G2105), .ZN(n880) );
  NAND2_X1 U578 ( .A1(G125), .A2(n880), .ZN(n533) );
  XNOR2_X1 U579 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n531) );
  NOR2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  XNOR2_X1 U581 ( .A(n531), .B(n530), .ZN(n874) );
  NAND2_X1 U582 ( .A1(G137), .A2(n874), .ZN(n532) );
  NAND2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n620) );
  NOR2_X1 U585 ( .A1(n620), .A2(G651), .ZN(n639) );
  NAND2_X1 U586 ( .A1(G47), .A2(n639), .ZN(n539) );
  NOR2_X1 U587 ( .A1(G543), .A2(n540), .ZN(n536) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n536), .Z(n537) );
  XNOR2_X2 U589 ( .A(KEYINPUT66), .B(n537), .ZN(n643) );
  NAND2_X1 U590 ( .A1(G60), .A2(n643), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n544) );
  NOR2_X1 U592 ( .A1(G543), .A2(G651), .ZN(n640) );
  NAND2_X1 U593 ( .A1(G85), .A2(n640), .ZN(n542) );
  NAND2_X1 U594 ( .A1(G72), .A2(n636), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n543) );
  OR2_X1 U596 ( .A1(n544), .A2(n543), .ZN(G290) );
  XNOR2_X1 U597 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U599 ( .A1(G111), .A2(n878), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G135), .A2(n874), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n880), .A2(G123), .ZN(n547) );
  XOR2_X1 U603 ( .A(KEYINPUT18), .B(n547), .Z(n548) );
  NOR2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U605 ( .A1(n875), .A2(G99), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n923) );
  XNOR2_X1 U607 ( .A(G2096), .B(n923), .ZN(n552) );
  OR2_X1 U608 ( .A1(G2100), .A2(n552), .ZN(G156) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  NAND2_X1 U612 ( .A1(G52), .A2(n639), .ZN(n554) );
  NAND2_X1 U613 ( .A1(G64), .A2(n643), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G90), .A2(n640), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G77), .A2(n636), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n557), .Z(n558) );
  NOR2_X1 U619 ( .A1(n559), .A2(n558), .ZN(G171) );
  NAND2_X1 U620 ( .A1(n640), .A2(G89), .ZN(n560) );
  XNOR2_X1 U621 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G76), .A2(n636), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U624 ( .A(n563), .B(KEYINPUT5), .ZN(n568) );
  NAND2_X1 U625 ( .A1(G51), .A2(n639), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G63), .A2(n643), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U628 ( .A(KEYINPUT6), .B(n566), .Z(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U630 ( .A(n569), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n827) );
  NAND2_X1 U635 ( .A1(n827), .A2(G567), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  NAND2_X1 U637 ( .A1(n640), .A2(G81), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G68), .A2(n636), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT13), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G43), .A2(n639), .ZN(n576) );
  XOR2_X1 U643 ( .A(KEYINPUT68), .B(n576), .Z(n579) );
  NAND2_X1 U644 ( .A1(n643), .A2(G56), .ZN(n577) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n577), .Z(n578) );
  NOR2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT69), .ZN(n977) );
  NAND2_X1 U649 ( .A1(n977), .A2(G860), .ZN(G153) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U652 ( .A1(G54), .A2(n639), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G79), .A2(n636), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G66), .A2(n643), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n640), .A2(G92), .ZN(n585) );
  XNOR2_X1 U657 ( .A(n585), .B(KEYINPUT70), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U659 ( .A(n589), .B(n588), .ZN(n590) );
  NOR2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n592) );
  INV_X1 U661 ( .A(n969), .ZN(n701) );
  INV_X1 U662 ( .A(G868), .ZN(n658) );
  NAND2_X1 U663 ( .A1(n701), .A2(n658), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U665 ( .A1(n640), .A2(G91), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G65), .A2(n643), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G53), .A2(n639), .ZN(n597) );
  XNOR2_X1 U669 ( .A(KEYINPUT67), .B(n597), .ZN(n598) );
  NOR2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n636), .A2(G78), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(G299) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n602), .B(KEYINPUT72), .ZN(n604) );
  NOR2_X1 U675 ( .A1(n658), .A2(G286), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n603), .ZN(G297) );
  INV_X1 U677 ( .A(G860), .ZN(n611) );
  NAND2_X1 U678 ( .A1(n611), .A2(G559), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n605), .A2(n969), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n606), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G559), .A2(n701), .ZN(n607) );
  NOR2_X1 U682 ( .A1(n658), .A2(n607), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n977), .A2(G868), .ZN(n608) );
  OR2_X1 U684 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G559), .A2(n969), .ZN(n610) );
  XNOR2_X1 U686 ( .A(n610), .B(n977), .ZN(n655) );
  NAND2_X1 U687 ( .A1(n611), .A2(n655), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n640), .A2(G93), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G67), .A2(n643), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G55), .A2(n639), .ZN(n614) );
  XNOR2_X1 U692 ( .A(KEYINPUT73), .B(n614), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n636), .A2(G80), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n657) );
  XNOR2_X1 U696 ( .A(n619), .B(n657), .ZN(G145) );
  NAND2_X1 U697 ( .A1(G87), .A2(n620), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G49), .A2(n639), .ZN(n622) );
  NAND2_X1 U699 ( .A1(G74), .A2(G651), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U701 ( .A1(n643), .A2(n623), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U703 ( .A(n626), .B(KEYINPUT74), .ZN(G288) );
  NAND2_X1 U704 ( .A1(n639), .A2(G50), .ZN(n627) );
  XOR2_X1 U705 ( .A(KEYINPUT77), .B(n627), .Z(n629) );
  NAND2_X1 U706 ( .A1(G62), .A2(n643), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U708 ( .A(KEYINPUT78), .B(n630), .ZN(n635) );
  NAND2_X1 U709 ( .A1(G88), .A2(n640), .ZN(n632) );
  NAND2_X1 U710 ( .A1(G75), .A2(n636), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U712 ( .A(KEYINPUT79), .B(n633), .Z(n634) );
  NOR2_X1 U713 ( .A1(n635), .A2(n634), .ZN(G166) );
  NAND2_X1 U714 ( .A1(n636), .A2(G73), .ZN(n638) );
  XNOR2_X1 U715 ( .A(KEYINPUT2), .B(KEYINPUT76), .ZN(n637) );
  XNOR2_X1 U716 ( .A(n638), .B(n637), .ZN(n648) );
  NAND2_X1 U717 ( .A1(G48), .A2(n639), .ZN(n642) );
  NAND2_X1 U718 ( .A1(G86), .A2(n640), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U720 ( .A1(G61), .A2(n643), .ZN(n644) );
  XNOR2_X1 U721 ( .A(KEYINPUT75), .B(n644), .ZN(n645) );
  NOR2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(G305) );
  INV_X1 U724 ( .A(G299), .ZN(n710) );
  XNOR2_X1 U725 ( .A(n710), .B(n657), .ZN(n654) );
  XNOR2_X1 U726 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n650) );
  XNOR2_X1 U727 ( .A(G290), .B(G166), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U729 ( .A(G288), .B(n651), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n652), .B(G305), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n654), .B(n653), .ZN(n897) );
  XNOR2_X1 U732 ( .A(n655), .B(n897), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n656), .A2(G868), .ZN(n660) );
  NAND2_X1 U734 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U736 ( .A1(G2078), .A2(G2084), .ZN(n661) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n662), .ZN(n664) );
  XOR2_X1 U739 ( .A(KEYINPUT21), .B(KEYINPUT81), .Z(n663) );
  XNOR2_X1 U740 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n665), .A2(G2072), .ZN(n666) );
  XNOR2_X1 U742 ( .A(n666), .B(KEYINPUT82), .ZN(G158) );
  NAND2_X1 U743 ( .A1(G69), .A2(G120), .ZN(n667) );
  NOR2_X1 U744 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U745 ( .A1(G108), .A2(n668), .ZN(n918) );
  NAND2_X1 U746 ( .A1(G567), .A2(n918), .ZN(n669) );
  XNOR2_X1 U747 ( .A(n669), .B(KEYINPUT83), .ZN(n674) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n670) );
  XNOR2_X1 U749 ( .A(KEYINPUT22), .B(n670), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n671), .A2(G96), .ZN(n672) );
  OR2_X1 U751 ( .A1(G218), .A2(n672), .ZN(n919) );
  AND2_X1 U752 ( .A1(G2106), .A2(n919), .ZN(n673) );
  NOR2_X1 U753 ( .A1(n674), .A2(n673), .ZN(G319) );
  INV_X1 U754 ( .A(G319), .ZN(n676) );
  NAND2_X1 U755 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U756 ( .A1(n676), .A2(n675), .ZN(n830) );
  NAND2_X1 U757 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U758 ( .A1(G138), .A2(n874), .ZN(n678) );
  NAND2_X1 U759 ( .A1(G102), .A2(n875), .ZN(n677) );
  NAND2_X1 U760 ( .A1(n678), .A2(n677), .ZN(n684) );
  NAND2_X1 U761 ( .A1(n880), .A2(G126), .ZN(n679) );
  XNOR2_X1 U762 ( .A(n679), .B(KEYINPUT84), .ZN(n681) );
  NAND2_X1 U763 ( .A1(G114), .A2(n878), .ZN(n680) );
  NAND2_X1 U764 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U765 ( .A(KEYINPUT85), .B(n682), .Z(n683) );
  NOR2_X1 U766 ( .A1(n684), .A2(n683), .ZN(G164) );
  XOR2_X1 U767 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NOR2_X1 U768 ( .A1(G164), .A2(G1384), .ZN(n759) );
  NAND2_X1 U769 ( .A1(G40), .A2(G160), .ZN(n685) );
  XNOR2_X1 U770 ( .A(KEYINPUT87), .B(n685), .ZN(n757) );
  INV_X1 U771 ( .A(n704), .ZN(n728) );
  INV_X1 U772 ( .A(G1961), .ZN(n993) );
  NAND2_X1 U773 ( .A1(n728), .A2(n993), .ZN(n687) );
  XNOR2_X1 U774 ( .A(G2078), .B(KEYINPUT25), .ZN(n956) );
  NAND2_X1 U775 ( .A1(n704), .A2(n956), .ZN(n686) );
  NAND2_X1 U776 ( .A1(n687), .A2(n686), .ZN(n722) );
  AND2_X1 U777 ( .A1(n722), .A2(G171), .ZN(n688) );
  XNOR2_X1 U778 ( .A(n688), .B(KEYINPUT95), .ZN(n717) );
  INV_X1 U779 ( .A(n704), .ZN(n718) );
  NAND2_X1 U780 ( .A1(G1348), .A2(n718), .ZN(n690) );
  NAND2_X1 U781 ( .A1(n704), .A2(G2067), .ZN(n689) );
  NAND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U783 ( .A(n691), .B(KEYINPUT97), .Z(n700) );
  OR2_X1 U784 ( .A1(n701), .A2(n700), .ZN(n699) );
  NAND2_X1 U785 ( .A1(n704), .A2(G1996), .ZN(n692) );
  XNOR2_X1 U786 ( .A(n692), .B(KEYINPUT26), .ZN(n694) );
  NAND2_X1 U787 ( .A1(G1341), .A2(n728), .ZN(n693) );
  NAND2_X1 U788 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U789 ( .A1(n977), .A2(n697), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n709) );
  NAND2_X1 U793 ( .A1(n704), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U794 ( .A(n705), .B(KEYINPUT27), .ZN(n707) );
  AND2_X1 U795 ( .A1(G1956), .A2(n728), .ZN(n706) );
  NOR2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U797 ( .A1(n711), .A2(n710), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n714) );
  NOR2_X1 U799 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U800 ( .A(n712), .B(KEYINPUT28), .Z(n713) );
  NAND2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U802 ( .A(n715), .B(KEYINPUT29), .Z(n716) );
  NAND2_X1 U803 ( .A1(n717), .A2(n716), .ZN(n727) );
  NAND2_X1 U804 ( .A1(G8), .A2(n718), .ZN(n791) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n791), .ZN(n742) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n728), .ZN(n738) );
  NOR2_X1 U807 ( .A1(n742), .A2(n738), .ZN(n719) );
  NAND2_X1 U808 ( .A1(G8), .A2(n719), .ZN(n720) );
  XNOR2_X1 U809 ( .A(KEYINPUT30), .B(n720), .ZN(n721) );
  NOR2_X1 U810 ( .A1(G168), .A2(n721), .ZN(n724) );
  NOR2_X1 U811 ( .A1(G171), .A2(n722), .ZN(n723) );
  NOR2_X1 U812 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U813 ( .A(KEYINPUT31), .B(n725), .Z(n726) );
  NAND2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n740) );
  NAND2_X1 U815 ( .A1(n740), .A2(G286), .ZN(n736) );
  INV_X1 U816 ( .A(G8), .ZN(n734) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n791), .ZN(n730) );
  NOR2_X1 U818 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U819 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U820 ( .A(KEYINPUT98), .B(n731), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n732), .A2(G303), .ZN(n733) );
  OR2_X1 U822 ( .A1(n734), .A2(n733), .ZN(n735) );
  AND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U824 ( .A1(G8), .A2(n738), .ZN(n739) );
  NAND2_X1 U825 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U826 ( .A1(G303), .A2(G1971), .ZN(n744) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n751) );
  OR2_X1 U828 ( .A1(n744), .A2(n751), .ZN(n988) );
  NOR2_X1 U829 ( .A1(n783), .A2(n988), .ZN(n745) );
  NOR2_X1 U830 ( .A1(n745), .A2(n791), .ZN(n748) );
  INV_X1 U831 ( .A(KEYINPUT99), .ZN(n746) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n973) );
  AND2_X1 U833 ( .A1(n746), .A2(n973), .ZN(n747) );
  AND2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n749), .A2(KEYINPUT33), .ZN(n756) );
  NAND2_X1 U836 ( .A1(n751), .A2(KEYINPUT33), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n746), .A2(n750), .ZN(n753) );
  NAND2_X1 U838 ( .A1(n751), .A2(KEYINPUT99), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U840 ( .A1(n791), .A2(n754), .ZN(n755) );
  NOR2_X1 U841 ( .A1(n756), .A2(n755), .ZN(n782) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n984) );
  INV_X1 U843 ( .A(n757), .ZN(n758) );
  NOR2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n822) );
  NAND2_X1 U845 ( .A1(G117), .A2(n878), .ZN(n761) );
  NAND2_X1 U846 ( .A1(G141), .A2(n874), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n765) );
  NAND2_X1 U848 ( .A1(G105), .A2(n875), .ZN(n762) );
  XNOR2_X1 U849 ( .A(n762), .B(KEYINPUT93), .ZN(n763) );
  XNOR2_X1 U850 ( .A(n763), .B(KEYINPUT38), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n880), .A2(G129), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n887) );
  NAND2_X1 U854 ( .A1(G1996), .A2(n887), .ZN(n778) );
  NAND2_X1 U855 ( .A1(G131), .A2(n874), .ZN(n768) );
  XOR2_X1 U856 ( .A(KEYINPUT92), .B(n768), .Z(n774) );
  NAND2_X1 U857 ( .A1(n880), .A2(G119), .ZN(n769) );
  XNOR2_X1 U858 ( .A(n769), .B(KEYINPUT90), .ZN(n771) );
  NAND2_X1 U859 ( .A1(G107), .A2(n878), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U861 ( .A(KEYINPUT91), .B(n772), .Z(n773) );
  NOR2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n875), .A2(G95), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n893) );
  NAND2_X1 U865 ( .A1(G1991), .A2(n893), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n926) );
  NAND2_X1 U867 ( .A1(n822), .A2(n926), .ZN(n811) );
  XNOR2_X1 U868 ( .A(G1986), .B(G290), .ZN(n972) );
  NAND2_X1 U869 ( .A1(n822), .A2(n972), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n811), .A2(n779), .ZN(n795) );
  INV_X1 U871 ( .A(n795), .ZN(n780) );
  AND2_X1 U872 ( .A1(n984), .A2(n780), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n797) );
  INV_X1 U874 ( .A(n783), .ZN(n786) );
  NOR2_X1 U875 ( .A1(G2090), .A2(G303), .ZN(n784) );
  NAND2_X1 U876 ( .A1(G8), .A2(n784), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n787) );
  AND2_X1 U878 ( .A1(n787), .A2(n791), .ZN(n793) );
  NOR2_X1 U879 ( .A1(G1981), .A2(G305), .ZN(n788) );
  XOR2_X1 U880 ( .A(n788), .B(KEYINPUT94), .Z(n789) );
  XNOR2_X1 U881 ( .A(KEYINPUT24), .B(n789), .ZN(n790) );
  NOR2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n794) );
  OR2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n809) );
  XNOR2_X1 U886 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  NAND2_X1 U887 ( .A1(G128), .A2(n880), .ZN(n799) );
  NAND2_X1 U888 ( .A1(G116), .A2(n878), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U890 ( .A(KEYINPUT35), .B(n800), .ZN(n806) );
  NAND2_X1 U891 ( .A1(G140), .A2(n874), .ZN(n802) );
  NAND2_X1 U892 ( .A1(G104), .A2(n875), .ZN(n801) );
  NAND2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n804) );
  XOR2_X1 U894 ( .A(KEYINPUT34), .B(KEYINPUT88), .Z(n803) );
  XNOR2_X1 U895 ( .A(n804), .B(n803), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U897 ( .A(KEYINPUT36), .B(n807), .Z(n888) );
  OR2_X1 U898 ( .A1(n819), .A2(n888), .ZN(n808) );
  XNOR2_X1 U899 ( .A(n808), .B(KEYINPUT89), .ZN(n943) );
  NAND2_X1 U900 ( .A1(n822), .A2(n943), .ZN(n817) );
  NAND2_X1 U901 ( .A1(n809), .A2(n817), .ZN(n810) );
  XNOR2_X1 U902 ( .A(n810), .B(KEYINPUT100), .ZN(n825) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n887), .ZN(n928) );
  INV_X1 U904 ( .A(n811), .ZN(n814) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n893), .ZN(n922) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n922), .A2(n812), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U909 ( .A1(n928), .A2(n815), .ZN(n816) );
  XNOR2_X1 U910 ( .A(n816), .B(KEYINPUT39), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n888), .A2(n819), .ZN(n930) );
  NAND2_X1 U913 ( .A1(n820), .A2(n930), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U915 ( .A(KEYINPUT101), .B(n823), .Z(n824) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U917 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U920 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(G188) );
  XOR2_X1 U923 ( .A(G2100), .B(G2096), .Z(n832) );
  XNOR2_X1 U924 ( .A(KEYINPUT42), .B(G2678), .ZN(n831) );
  XNOR2_X1 U925 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U926 ( .A(KEYINPUT43), .B(G2090), .Z(n834) );
  XNOR2_X1 U927 ( .A(G2067), .B(G2072), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U929 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U930 ( .A(G2078), .B(G2084), .ZN(n837) );
  XNOR2_X1 U931 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U932 ( .A(G1966), .B(G1986), .Z(n840) );
  XNOR2_X1 U933 ( .A(G1996), .B(G1991), .ZN(n839) );
  XNOR2_X1 U934 ( .A(n840), .B(n839), .ZN(n850) );
  XOR2_X1 U935 ( .A(KEYINPUT104), .B(KEYINPUT41), .Z(n842) );
  XNOR2_X1 U936 ( .A(G1956), .B(G2474), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U938 ( .A(G1976), .B(G1981), .Z(n844) );
  XNOR2_X1 U939 ( .A(G1961), .B(G1971), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U941 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U942 ( .A(KEYINPUT106), .B(KEYINPUT105), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U944 ( .A(n850), .B(n849), .ZN(G229) );
  NAND2_X1 U945 ( .A1(G124), .A2(n880), .ZN(n851) );
  XOR2_X1 U946 ( .A(KEYINPUT44), .B(n851), .Z(n852) );
  XNOR2_X1 U947 ( .A(n852), .B(KEYINPUT107), .ZN(n854) );
  NAND2_X1 U948 ( .A1(G112), .A2(n878), .ZN(n853) );
  NAND2_X1 U949 ( .A1(n854), .A2(n853), .ZN(n858) );
  NAND2_X1 U950 ( .A1(G136), .A2(n874), .ZN(n856) );
  NAND2_X1 U951 ( .A1(G100), .A2(n875), .ZN(n855) );
  NAND2_X1 U952 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U953 ( .A1(n858), .A2(n857), .ZN(G162) );
  XOR2_X1 U954 ( .A(KEYINPUT112), .B(KEYINPUT48), .Z(n860) );
  XNOR2_X1 U955 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U957 ( .A(KEYINPUT109), .B(n861), .ZN(n872) );
  NAND2_X1 U958 ( .A1(G130), .A2(n880), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G118), .A2(n878), .ZN(n862) );
  NAND2_X1 U960 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U961 ( .A1(G142), .A2(n874), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G106), .A2(n875), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U964 ( .A(KEYINPUT45), .B(n866), .Z(n867) );
  XNOR2_X1 U965 ( .A(KEYINPUT108), .B(n867), .ZN(n868) );
  NOR2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U967 ( .A(n923), .B(n870), .ZN(n871) );
  XNOR2_X1 U968 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U969 ( .A(G162), .B(n873), .ZN(n892) );
  NAND2_X1 U970 ( .A1(G139), .A2(n874), .ZN(n877) );
  NAND2_X1 U971 ( .A1(G103), .A2(n875), .ZN(n876) );
  NAND2_X1 U972 ( .A1(n877), .A2(n876), .ZN(n886) );
  NAND2_X1 U973 ( .A1(n878), .A2(G115), .ZN(n879) );
  XNOR2_X1 U974 ( .A(n879), .B(KEYINPUT110), .ZN(n882) );
  NAND2_X1 U975 ( .A1(G127), .A2(n880), .ZN(n881) );
  NAND2_X1 U976 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U977 ( .A(KEYINPUT47), .B(n883), .ZN(n884) );
  XNOR2_X1 U978 ( .A(KEYINPUT111), .B(n884), .ZN(n885) );
  NOR2_X1 U979 ( .A1(n886), .A2(n885), .ZN(n933) );
  XNOR2_X1 U980 ( .A(n887), .B(n933), .ZN(n890) );
  XOR2_X1 U981 ( .A(G160), .B(n888), .Z(n889) );
  XNOR2_X1 U982 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U983 ( .A(n892), .B(n891), .ZN(n895) );
  XOR2_X1 U984 ( .A(n893), .B(G164), .Z(n894) );
  XNOR2_X1 U985 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U986 ( .A1(G37), .A2(n896), .ZN(G395) );
  XOR2_X1 U987 ( .A(n897), .B(G286), .Z(n899) );
  XNOR2_X1 U988 ( .A(n977), .B(G171), .ZN(n898) );
  XNOR2_X1 U989 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U990 ( .A(n900), .B(n969), .ZN(n901) );
  NOR2_X1 U991 ( .A1(G37), .A2(n901), .ZN(G397) );
  XNOR2_X1 U992 ( .A(G2446), .B(G2443), .ZN(n911) );
  XOR2_X1 U993 ( .A(G2430), .B(KEYINPUT103), .Z(n903) );
  XNOR2_X1 U994 ( .A(G2454), .B(G2435), .ZN(n902) );
  XNOR2_X1 U995 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U996 ( .A(G2438), .B(G2427), .Z(n905) );
  XNOR2_X1 U997 ( .A(G1348), .B(G1341), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U999 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1000 ( .A(KEYINPUT102), .B(G2451), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1002 ( .A(n911), .B(n910), .ZN(n912) );
  NAND2_X1 U1003 ( .A1(n912), .A2(G14), .ZN(n920) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n920), .ZN(n915) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1007 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1009 ( .A1(n917), .A2(n916), .ZN(G225) );
  XOR2_X1 U1010 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  INV_X1 U1012 ( .A(G120), .ZN(G236) );
  INV_X1 U1013 ( .A(G96), .ZN(G221) );
  INV_X1 U1014 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(G325) );
  INV_X1 U1016 ( .A(G325), .ZN(G261) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(n920), .ZN(G401) );
  XOR2_X1 U1019 ( .A(G160), .B(G2084), .Z(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n941) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1025 ( .A(KEYINPUT51), .B(n929), .Z(n931) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n939) );
  XNOR2_X1 U1027 ( .A(G164), .B(G2078), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(n932), .B(KEYINPUT115), .ZN(n935) );
  XOR2_X1 U1029 ( .A(G2072), .B(n933), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1031 ( .A(KEYINPUT116), .B(n936), .Z(n937) );
  XNOR2_X1 U1032 ( .A(KEYINPUT50), .B(n937), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n944), .ZN(n945) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n1025) );
  NAND2_X1 U1038 ( .A1(n945), .A2(n1025), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n946), .A2(G29), .ZN(n1032) );
  XNOR2_X1 U1040 ( .A(G25), .B(G1991), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(n947), .B(KEYINPUT117), .ZN(n955) );
  XNOR2_X1 U1042 ( .A(G2067), .B(G26), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(G28), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G32), .B(G1996), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(KEYINPUT118), .B(n951), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1050 ( .A(G27), .B(n956), .Z(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(KEYINPUT119), .B(n959), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n960), .B(KEYINPUT53), .ZN(n966) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(G34), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n961), .B(KEYINPUT120), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(G2084), .B(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G2090), .B(G35), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n1026) );
  NOR2_X1 U1060 ( .A1(G29), .A2(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n1026), .A2(n967), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n968), .ZN(n1030) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XNOR2_X1 U1064 ( .A(n969), .B(G1348), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(G1971), .A2(G303), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n983) );
  INV_X1 U1067 ( .A(n972), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(G1956), .B(G299), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n981) );
  XOR2_X1 U1071 ( .A(n977), .B(G1341), .Z(n979) );
  XNOR2_X1 U1072 ( .A(G301), .B(G1961), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n990) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G168), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1078 ( .A(KEYINPUT57), .B(n986), .Z(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n1023) );
  INV_X1 U1082 ( .A(G16), .ZN(n1021) );
  XOR2_X1 U1083 ( .A(G1966), .B(G21), .Z(n995) );
  XNOR2_X1 U1084 ( .A(n993), .B(G5), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n1008) );
  XNOR2_X1 U1086 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n996), .B(KEYINPUT60), .ZN(n1006) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(n997), .B(G4), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(G6), .B(G1981), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XOR2_X1 U1094 ( .A(KEYINPUT121), .B(G1956), .Z(n1002) );
  XNOR2_X1 U1095 ( .A(G20), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(n1006), .B(n1005), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT124), .B(n1009), .ZN(n1018) );
  XOR2_X1 U1100 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n1016) );
  XNOR2_X1 U1101 ( .A(G1986), .B(G24), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(G22), .B(G1971), .ZN(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(G1976), .B(KEYINPUT125), .ZN(n1012) );
  XNOR2_X1 U1105 ( .A(n1012), .B(G23), .ZN(n1013) );
  NAND2_X1 U1106 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1107 ( .A(n1016), .B(n1015), .ZN(n1017) );
  NAND2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1019), .Z(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1112 ( .A(n1024), .B(KEYINPUT127), .ZN(n1028) );
  OR2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

