//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g001(.A(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G162gat), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G141gat), .B(G148gat), .Z(new_n208));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n212));
  INV_X1    g011(.A(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(G141gat), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT74), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(new_n213), .B2(G141gat), .ZN(new_n218));
  INV_X1    g017(.A(G141gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n216), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT2), .B1(new_n205), .B2(KEYINPUT76), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n222), .A2(new_n204), .A3(new_n206), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n221), .A2(KEYINPUT77), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT77), .B1(new_n221), .B2(new_n223), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n202), .B(new_n211), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n226), .A2(KEYINPUT82), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT82), .B1(new_n226), .B2(new_n227), .ZN(new_n229));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230));
  INV_X1    g029(.A(G211gat), .ZN(new_n231));
  INV_X1    g030(.A(G218gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n230), .B1(KEYINPUT22), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n228), .A2(new_n229), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n211), .B1(new_n224), .B2(new_n225), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT78), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT77), .ZN(new_n241));
  AND2_X1   g040(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n242), .A2(new_n243), .A3(new_n219), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n218), .A2(new_n220), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n207), .A2(new_n222), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n241), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n221), .A2(KEYINPUT77), .A3(new_n223), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT78), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(new_n211), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n202), .B1(new_n236), .B2(KEYINPUT29), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n240), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G228gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT83), .B1(new_n238), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n257), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n251), .B1(new_n250), .B2(new_n211), .ZN(new_n261));
  AOI211_X1 g060(.A(KEYINPUT78), .B(new_n210), .C1(new_n248), .C2(new_n249), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n263), .B2(new_n253), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT83), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n226), .A2(new_n227), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT82), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n226), .A2(KEYINPUT82), .A3(new_n227), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n236), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n264), .A2(new_n265), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n259), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n253), .A2(new_n239), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n237), .B1(new_n226), .B2(new_n227), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n260), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G78gat), .B(G106gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT31), .ZN(new_n278));
  INV_X1    g077(.A(G50gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G22gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT84), .B(G22gat), .Z(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(KEYINPUT85), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n272), .A2(new_n275), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n238), .A2(KEYINPUT83), .A3(new_n258), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n265), .B1(new_n264), .B2(new_n270), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n275), .B(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n285), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n284), .B1(new_n272), .B2(new_n275), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n283), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n294));
  AND2_X1   g093(.A1(G113gat), .A2(G120gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(G113gat), .A2(G120gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G134gat), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G127gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n297), .B1(new_n295), .B2(new_n296), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n299), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(G127gat), .B(G134gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n295), .A2(new_n296), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n303), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n305), .A2(new_n306), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT27), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G183gat), .ZN(new_n318));
  INV_X1    g117(.A(G190gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT27), .B(G183gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(KEYINPUT28), .A3(new_n319), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT65), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT65), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(new_n330), .A3(new_n327), .ZN(new_n331));
  OR3_X1    g130(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n325), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  INV_X1    g135(.A(G169gat), .ZN(new_n337));
  INV_X1    g136(.A(G176gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT23), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  AND4_X1   g140(.A1(new_n336), .A2(new_n339), .A3(new_n341), .A4(new_n327), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n334), .A2(KEYINPUT24), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT24), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(G183gat), .A3(G190gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n315), .A2(new_n319), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT64), .ZN(new_n348));
  OR3_X1    g147(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n343), .A2(new_n345), .B1(new_n315), .B2(new_n319), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n339), .A2(new_n341), .A3(new_n327), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT25), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n314), .B1(new_n335), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT68), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n346), .A2(new_n347), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n339), .A2(new_n341), .A3(new_n327), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n360), .A2(KEYINPUT25), .B1(new_n350), .B2(new_n342), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n325), .A2(new_n333), .A3(new_n334), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n313), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT68), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(new_n313), .A3(new_n362), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n357), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G227gat), .A2(G233gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n294), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT33), .ZN(new_n371));
  XNOR2_X1  g170(.A(G15gat), .B(G43gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G71gat), .B(G99gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n370), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n374), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n366), .B1(new_n363), .B2(new_n364), .ZN(new_n377));
  AOI211_X1 g176(.A(KEYINPUT68), .B(new_n313), .C1(new_n361), .C2(new_n362), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n369), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n371), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n376), .B(new_n380), .C1(new_n370), .C2(KEYINPUT69), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n379), .A2(KEYINPUT69), .A3(KEYINPUT32), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n375), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n357), .A2(new_n365), .A3(new_n368), .A4(new_n366), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n384), .B(KEYINPUT34), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n385), .B(new_n375), .C1(new_n381), .C2(new_n382), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n293), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n335), .A2(new_n355), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(KEYINPUT29), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT72), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(KEYINPUT71), .ZN(new_n395));
  INV_X1    g194(.A(new_n391), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT71), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n335), .B2(new_n355), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT72), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n400), .B(new_n391), .C1(new_n392), .C2(KEYINPUT29), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n394), .A2(new_n399), .A3(new_n237), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n392), .A2(new_n396), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n395), .A2(new_n398), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n391), .A2(new_n227), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n236), .B(new_n403), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(G64gat), .ZN(new_n408));
  INV_X1    g207(.A(G92gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n402), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n402), .A2(new_n406), .ZN(new_n414));
  INV_X1    g213(.A(new_n410), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n402), .A2(new_n406), .A3(KEYINPUT30), .A4(new_n410), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT0), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(G57gat), .ZN(new_n422));
  INV_X1    g221(.A(G85gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n313), .B(new_n211), .C1(new_n224), .C2(new_n225), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT80), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n250), .A2(KEYINPUT80), .A3(new_n211), .A4(new_n313), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n240), .A2(new_n314), .A3(new_n252), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G225gat), .A2(G233gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT81), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT5), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n240), .A2(KEYINPUT3), .A3(new_n252), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n226), .A2(new_n314), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n427), .A2(new_n440), .A3(new_n428), .ZN(new_n441));
  XOR2_X1   g240(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n436), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT81), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n447), .A3(new_n433), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n435), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n437), .A2(new_n438), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n433), .A2(KEYINPUT5), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n425), .A2(new_n443), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n440), .B1(new_n427), .B2(new_n428), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n450), .B(new_n451), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n424), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(KEYINPUT86), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n457));
  AOI211_X1 g256(.A(new_n457), .B(new_n424), .C1(new_n449), .C2(new_n454), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n449), .A2(new_n424), .A3(new_n454), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n456), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n455), .A2(KEYINPUT6), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n390), .B(new_n419), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT35), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n383), .A2(KEYINPUT70), .A3(new_n386), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT70), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n387), .A2(new_n469), .A3(new_n388), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n293), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n463), .B1(new_n461), .B2(new_n455), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n416), .A2(KEYINPUT73), .A3(new_n417), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT73), .B1(new_n416), .B2(new_n417), .ZN(new_n474));
  INV_X1    g273(.A(new_n413), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n472), .A2(KEYINPUT35), .A3(new_n476), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n465), .A2(new_n466), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n456), .A2(new_n458), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT39), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n453), .A2(new_n452), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n437), .A2(new_n438), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n480), .B(new_n433), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n429), .A2(KEYINPUT4), .ZN(new_n484));
  INV_X1    g283(.A(new_n452), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n432), .B1(new_n486), .B2(new_n450), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT39), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n424), .B(new_n483), .C1(new_n487), .C2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT40), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n433), .B1(new_n481), .B2(new_n482), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT39), .A3(new_n488), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n494), .A2(KEYINPUT40), .A3(new_n424), .A4(new_n483), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n492), .A2(new_n495), .A3(new_n418), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n293), .B1(new_n479), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n454), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n447), .B1(new_n431), .B2(new_n433), .ZN(new_n499));
  AOI211_X1 g298(.A(KEYINPUT81), .B(new_n432), .C1(new_n429), .C2(new_n430), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n501), .B2(new_n446), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n457), .B1(new_n502), .B2(new_n424), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT6), .B1(new_n502), .B2(new_n424), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n455), .A2(KEYINPUT86), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT38), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n402), .A2(new_n406), .A3(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n509), .A2(new_n415), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n414), .A2(KEYINPUT37), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n237), .B(new_n403), .C1(new_n404), .C2(new_n405), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n394), .A2(new_n401), .A3(new_n399), .ZN(new_n514));
  OAI211_X1 g313(.A(KEYINPUT37), .B(new_n513), .C1(new_n514), .C2(new_n237), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n515), .A2(new_n509), .A3(new_n507), .A4(new_n415), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n411), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n506), .A2(new_n463), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n497), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n388), .A2(new_n469), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n370), .A2(KEYINPUT69), .ZN(new_n522));
  INV_X1    g321(.A(new_n382), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n374), .B1(new_n379), .B2(new_n371), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n385), .B1(new_n525), .B2(new_n375), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT36), .B1(new_n527), .B2(new_n467), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n389), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n472), .A2(new_n476), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n293), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n520), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n478), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G43gat), .B(G50gat), .Z(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT89), .B(KEYINPUT15), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT90), .ZN(new_n539));
  NOR2_X1   g338(.A1(G29gat), .A2(G36gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT14), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT15), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(G29gat), .B2(G36gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G29gat), .ZN(new_n549));
  INV_X1    g348(.A(G36gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n542), .A2(new_n547), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n544), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT91), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n556), .A3(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559));
  INV_X1    g358(.A(G1gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT16), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(G1gat), .B2(new_n559), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G8gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT93), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n558), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n546), .A2(KEYINPUT17), .A3(new_n553), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(new_n564), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n558), .B2(KEYINPUT17), .ZN(new_n570));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT92), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n567), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT18), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n567), .A2(new_n570), .A3(KEYINPUT94), .A4(new_n573), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n572), .B(KEYINPUT13), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n558), .A2(new_n565), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(new_n566), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n579), .B(new_n582), .C1(new_n577), .C2(new_n574), .ZN(new_n583));
  XOR2_X1   g382(.A(G169gat), .B(G197gat), .Z(new_n584));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT12), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n582), .B(new_n590), .C1(new_n574), .C2(new_n577), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n591), .B1(new_n579), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n576), .A2(KEYINPUT95), .A3(new_n577), .A4(new_n578), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n583), .A2(new_n589), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n535), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n597), .A2(KEYINPUT96), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(KEYINPUT96), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G85gat), .A2(G92gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT7), .ZN(new_n602));
  NAND2_X1  g401(.A1(G99gat), .A2(G106gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(KEYINPUT8), .A2(new_n603), .B1(new_n423), .B2(new_n409), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G99gat), .B(G106gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n568), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n558), .B2(KEYINPUT17), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n555), .A2(new_n557), .A3(new_n607), .ZN(new_n610));
  NAND3_X1  g409(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G190gat), .B(G218gat), .Z(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n609), .A2(new_n610), .A3(new_n611), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G134gat), .B(G162gat), .Z(new_n618));
  AOI21_X1  g417(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n620), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n614), .A2(KEYINPUT100), .A3(new_n623), .A4(new_n616), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT97), .Z(new_n629));
  OR2_X1    g428(.A1(G71gat), .A2(G78gat), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G57gat), .B(G64gat), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n631), .B1(new_n630), .B2(new_n628), .ZN(new_n634));
  AND2_X1   g433(.A1(KEYINPUT98), .A2(G57gat), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n635), .A2(G64gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(G64gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n565), .B1(new_n627), .B2(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n640), .A2(KEYINPUT99), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(KEYINPUT99), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n627), .ZN(new_n644));
  XNOR2_X1  g443(.A(G127gat), .B(G155gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n641), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n651));
  NAND2_X1  g450(.A1(G231gat), .A2(G233gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G183gat), .B(G211gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n647), .A2(new_n649), .A3(new_n655), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n626), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(G230gat), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n256), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n607), .B(new_n639), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n607), .A2(KEYINPUT10), .A3(new_n633), .A4(new_n638), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n662), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n663), .A2(new_n661), .A3(new_n256), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G120gat), .B(G148gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G176gat), .ZN(new_n671));
  INV_X1    g470(.A(G204gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n669), .A2(new_n674), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n660), .A2(KEYINPUT101), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT101), .B1(new_n660), .B2(new_n678), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n600), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n472), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT102), .B(G1gat), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1324gat));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  NAND4_X1  g486(.A1(new_n682), .A2(KEYINPUT42), .A3(new_n418), .A4(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689));
  OAI221_X1 g488(.A(new_n418), .B1(new_n679), .B2(new_n680), .C1(new_n598), .C2(new_n599), .ZN(new_n690));
  INV_X1    g489(.A(new_n687), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(G8gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n688), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT103), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n688), .A2(new_n692), .A3(new_n696), .A4(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1325gat));
  INV_X1    g497(.A(G15gat), .ZN(new_n699));
  INV_X1    g498(.A(new_n389), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n682), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n531), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n682), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n701), .B1(new_n704), .B2(new_n699), .ZN(G1326gat));
  NAND2_X1  g504(.A1(new_n682), .A2(new_n293), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  OR2_X1    g507(.A1(new_n598), .A2(new_n599), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n657), .A2(new_n658), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n710), .A2(new_n625), .A3(new_n677), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n709), .A2(new_n549), .A3(new_n683), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n535), .A2(KEYINPUT105), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n478), .A2(new_n534), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n717));
  NAND4_X1  g516(.A1(new_n714), .A2(new_n626), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n535), .A2(new_n626), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(KEYINPUT44), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n625), .B1(new_n478), .B2(new_n534), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n722), .A2(KEYINPUT104), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n718), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n677), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n725), .A2(new_n596), .A3(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n727), .A2(new_n683), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n713), .B1(new_n549), .B2(new_n728), .ZN(G1328gat));
  NAND4_X1  g528(.A1(new_n709), .A2(new_n550), .A3(new_n418), .A4(new_n711), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT46), .Z(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n418), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G36gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1329gat));
  INV_X1    g533(.A(G43gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n709), .A2(new_n735), .A3(new_n700), .A4(new_n711), .ZN(new_n736));
  AND4_X1   g535(.A1(new_n702), .A2(new_n725), .A3(new_n596), .A4(new_n726), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(new_n735), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(KEYINPUT47), .B(new_n736), .C1(new_n737), .C2(new_n735), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(G1330gat));
  NAND4_X1  g541(.A1(new_n709), .A2(new_n279), .A3(new_n293), .A4(new_n711), .ZN(new_n743));
  AND4_X1   g542(.A1(new_n293), .A2(new_n725), .A3(new_n596), .A4(new_n726), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(new_n279), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT48), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  OAI221_X1 g547(.A(new_n743), .B1(new_n746), .B2(KEYINPUT48), .C1(new_n744), .C2(new_n279), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1331gat));
  AND2_X1   g549(.A1(new_n714), .A2(new_n716), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n595), .A2(new_n660), .A3(new_n677), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n472), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT108), .B(G57gat), .Z(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT109), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n754), .B(new_n756), .ZN(G1332gat));
  NOR2_X1   g556(.A1(new_n753), .A2(new_n419), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  OAI21_X1  g561(.A(G71gat), .B1(new_n753), .B2(new_n531), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n389), .A2(G71gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n753), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT50), .Z(G1334gat));
  INV_X1    g565(.A(new_n293), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n753), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT110), .B(G78gat), .Z(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1335gat));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n595), .A2(new_n659), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n678), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n725), .A2(new_n683), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n720), .A2(new_n772), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT51), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n722), .A2(new_n595), .A3(new_n659), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(KEYINPUT111), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT111), .B1(new_n776), .B2(new_n779), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n683), .A2(new_n423), .A3(new_n677), .ZN(new_n784));
  OAI221_X1 g583(.A(new_n771), .B1(new_n774), .B2(new_n423), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n774), .A2(new_n423), .ZN(new_n786));
  INV_X1    g585(.A(new_n782), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n784), .B1(new_n787), .B2(new_n780), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT112), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(G1336gat));
  AND2_X1   g589(.A1(new_n725), .A2(new_n773), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n409), .B1(new_n791), .B2(new_n418), .ZN(new_n792));
  NOR2_X1   g591(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n777), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n677), .A2(new_n409), .A3(new_n418), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n776), .A2(new_n779), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n801), .B2(new_n796), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n798), .B1(new_n792), .B2(new_n802), .ZN(G1337gat));
  AND2_X1   g602(.A1(new_n791), .A2(new_n702), .ZN(new_n804));
  INV_X1    g603(.A(G99gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n700), .A2(new_n805), .A3(new_n677), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT114), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n804), .A2(new_n805), .B1(new_n783), .B2(new_n807), .ZN(G1338gat));
  NOR3_X1   g607(.A1(new_n767), .A2(G106gat), .A3(new_n678), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT115), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT53), .B1(new_n795), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n725), .A2(new_n293), .A3(new_n773), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(G106gat), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n725), .A2(KEYINPUT116), .A3(new_n293), .A4(new_n773), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(G106gat), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n809), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n813), .B1(new_n819), .B2(new_n820), .ZN(G1339gat));
  NOR2_X1   g620(.A1(new_n595), .A2(G113gat), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n593), .A2(new_n594), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n573), .B1(new_n567), .B2(new_n570), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n581), .A2(new_n566), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n824), .A2(KEYINPUT117), .B1(new_n825), .B2(new_n580), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n588), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n823), .A2(new_n828), .A3(new_n677), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n667), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n665), .A2(new_n666), .A3(new_n662), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n673), .B1(new_n667), .B2(new_n830), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n675), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT55), .B1(new_n833), .B2(new_n834), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n829), .B(new_n625), .C1(new_n595), .C2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n828), .A3(new_n838), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n710), .B1(new_n841), .B2(new_n626), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n595), .A2(new_n660), .A3(new_n678), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(KEYINPUT118), .A3(new_n844), .ZN(new_n848));
  AND4_X1   g647(.A1(new_n683), .A2(new_n847), .A3(new_n419), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n471), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n850), .A2(KEYINPUT119), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(KEYINPUT119), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n822), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n390), .ZN(new_n854));
  OAI21_X1  g653(.A(G113gat), .B1(new_n854), .B2(new_n595), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(G1340gat));
  NOR2_X1   g655(.A1(new_n678), .A2(G120gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n851), .B2(new_n852), .ZN(new_n858));
  OAI21_X1  g657(.A(G120gat), .B1(new_n854), .B2(new_n678), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1341gat));
  OAI21_X1  g659(.A(G127gat), .B1(new_n854), .B2(new_n659), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n710), .A2(new_n299), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n850), .B2(new_n862), .ZN(G1342gat));
  OAI21_X1  g662(.A(G134gat), .B1(new_n854), .B2(new_n625), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n625), .A2(G134gat), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT56), .B1(new_n850), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n849), .A2(new_n868), .A3(new_n471), .A4(new_n865), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n864), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT120), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n864), .A2(new_n867), .A3(new_n869), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1343gat));
  NAND3_X1  g673(.A1(new_n847), .A2(new_n293), .A3(new_n848), .ZN(new_n875));
  XOR2_X1   g674(.A(KEYINPUT122), .B(KEYINPUT57), .Z(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n767), .A2(new_n877), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n875), .A2(new_n876), .B1(new_n845), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n531), .A2(new_n683), .A3(new_n419), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT121), .Z(new_n881));
  NOR2_X1   g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n219), .B1(new_n882), .B2(new_n596), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n702), .A2(new_n767), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n849), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n596), .A2(new_n219), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT58), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n879), .A2(new_n595), .A3(new_n881), .ZN(new_n890));
  OAI221_X1 g689(.A(new_n889), .B1(new_n885), .B2(new_n886), .C1(new_n890), .C2(new_n219), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(G1344gat));
  OAI21_X1  g691(.A(KEYINPUT59), .B1(new_n885), .B2(new_n678), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n214), .A3(new_n215), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n875), .A2(new_n876), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n595), .B1(new_n679), .B2(new_n680), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n897), .A2(new_n843), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n896), .B(new_n877), .C1(new_n898), .C2(new_n767), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n767), .B1(new_n897), .B2(new_n843), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT123), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n677), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  OAI211_X1 g702(.A(KEYINPUT59), .B(G148gat), .C1(new_n903), .C2(new_n881), .ZN(new_n904));
  INV_X1    g703(.A(new_n882), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n678), .A2(KEYINPUT59), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n894), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(G1345gat));
  INV_X1    g706(.A(new_n885), .ZN(new_n908));
  XNOR2_X1  g707(.A(KEYINPUT76), .B(G155gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n710), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n905), .A2(new_n659), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n909), .ZN(G1346gat));
  OAI21_X1  g711(.A(G162gat), .B1(new_n905), .B2(new_n625), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n908), .A2(new_n203), .A3(new_n626), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1347gat));
  AND3_X1   g714(.A1(new_n847), .A2(new_n472), .A3(new_n848), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n418), .A3(new_n390), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n917), .A2(new_n337), .A3(new_n595), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n471), .A2(new_n418), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT124), .Z(new_n920));
  NAND4_X1  g719(.A1(new_n847), .A2(new_n472), .A3(new_n848), .A4(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n596), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n918), .A2(new_n923), .ZN(G1348gat));
  OAI21_X1  g723(.A(G176gat), .B1(new_n917), .B2(new_n678), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n922), .A2(new_n338), .A3(new_n677), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1349gat));
  NAND2_X1  g726(.A1(new_n710), .A2(new_n323), .ZN(new_n928));
  OR3_X1    g727(.A1(new_n921), .A2(KEYINPUT125), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT125), .B1(new_n921), .B2(new_n928), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G183gat), .B1(new_n917), .B2(new_n659), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT60), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n917), .B2(new_n625), .ZN(new_n938));
  NOR2_X1   g737(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n319), .A3(new_n626), .ZN(new_n941));
  XNOR2_X1  g740(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n940), .B(new_n941), .C1(new_n938), .C2(new_n942), .ZN(G1351gat));
  INV_X1    g742(.A(G197gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n916), .A2(new_n418), .A3(new_n884), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n595), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n702), .A2(new_n683), .A3(new_n419), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n595), .A2(new_n944), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n947), .B(new_n948), .C1(new_n895), .C2(new_n902), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(G1352gat));
  INV_X1    g751(.A(new_n947), .ZN(new_n953));
  OAI21_X1  g752(.A(G204gat), .B1(new_n903), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n677), .A2(new_n672), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT62), .B1(new_n945), .B2(new_n955), .ZN(new_n956));
  OR3_X1    g755(.A1(new_n945), .A2(KEYINPUT62), .A3(new_n955), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(G1353gat));
  OAI211_X1 g757(.A(new_n710), .B(new_n947), .C1(new_n895), .C2(new_n902), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n710), .A2(new_n231), .ZN(new_n962));
  OAI22_X1  g761(.A1(new_n960), .A2(new_n961), .B1(new_n945), .B2(new_n962), .ZN(G1354gat));
  OAI21_X1  g762(.A(new_n947), .B1(new_n895), .B2(new_n902), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n964), .A2(new_n232), .A3(new_n625), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n945), .A2(new_n625), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n232), .B2(new_n966), .ZN(G1355gat));
endmodule


