//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n211), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(KEYINPUT3), .ZN(new_n244));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n250), .B1(new_n251), .B2(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n217), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT65), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(KEYINPUT65), .A2(G33), .A3(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(new_n255), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT65), .B1(G33), .B2(G41), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n217), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(new_n274), .B2(new_n263), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n269), .B1(G226), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n260), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G190), .ZN(new_n279));
  OAI21_X1  g0079(.A(G200), .B1(new_n260), .B2(new_n277), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n217), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT66), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT66), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(new_n285), .A3(new_n217), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n209), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G150), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n288), .A2(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n203), .A2(G50), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n209), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n287), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G13), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n297), .A2(new_n209), .A3(G1), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n296), .B1(G50), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n208), .A2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G50), .ZN(new_n302));
  XOR2_X1   g0102(.A(new_n302), .B(KEYINPUT67), .Z(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(new_n284), .A3(new_n286), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT69), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n306), .A2(KEYINPUT9), .B1(new_n307), .B2(KEYINPUT10), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n306), .A2(KEYINPUT9), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n281), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n311), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n281), .A2(new_n313), .A3(new_n308), .A4(new_n309), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n278), .A2(new_n315), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n316), .B1(G169), .B2(new_n278), .C1(new_n305), .C2(new_n300), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT17), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n264), .A2(G232), .A3(new_n265), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G223), .A2(G1698), .ZN(new_n321));
  INV_X1    g0121(.A(G226), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(G1698), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n323), .A2(new_n248), .B1(G33), .B2(G87), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n320), .B(new_n268), .C1(new_n324), .C2(new_n257), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n325), .A2(G200), .ZN(new_n326));
  INV_X1    g0126(.A(G190), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G58), .A2(G68), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT78), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT78), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(G58), .A3(G68), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n333), .A3(new_n203), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n291), .A2(G159), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT79), .ZN(new_n338));
  AND2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT7), .B1(new_n341), .B2(new_n209), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n246), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n247), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(G68), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT79), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n335), .A2(new_n346), .A3(new_n336), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n338), .A2(KEYINPUT16), .A3(new_n345), .A4(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n246), .A2(new_n209), .A3(new_n247), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n202), .B1(new_n352), .B2(new_n343), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n349), .B1(new_n353), .B2(new_n337), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n348), .A2(new_n283), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n288), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n301), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n304), .A2(new_n357), .B1(new_n299), .B2(new_n356), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n329), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n319), .B1(new_n360), .B2(KEYINPUT81), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n354), .A2(new_n283), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n358), .B1(new_n362), .B2(new_n348), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT81), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT17), .A4(new_n329), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT18), .ZN(new_n367));
  INV_X1    g0167(.A(new_n324), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n269), .B1(new_n368), .B2(new_n258), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT80), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n369), .A2(new_n370), .A3(new_n315), .A4(new_n320), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT80), .B1(new_n325), .B2(G179), .ZN(new_n372));
  INV_X1    g0172(.A(G169), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n325), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n367), .B1(new_n363), .B2(new_n375), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n355), .A2(new_n359), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT18), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n356), .A2(new_n291), .B1(G20), .B2(G77), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n289), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(new_n283), .B1(new_n251), .B2(new_n298), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n298), .A2(new_n283), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(G77), .A3(new_n301), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT68), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n390));
  INV_X1    g0190(.A(G107), .ZN(new_n391));
  INV_X1    g0191(.A(G238), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n390), .B1(new_n391), .B2(new_n248), .C1(new_n252), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n258), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n269), .B1(G244), .B2(new_n275), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n389), .B1(new_n397), .B2(G190), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(G200), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n315), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n396), .A2(new_n373), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n389), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NOR4_X1   g0204(.A1(new_n318), .A2(new_n366), .A3(new_n381), .A4(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(G232), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT70), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT70), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n248), .A2(new_n408), .A3(G232), .A4(G1698), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G97), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n248), .A2(G226), .A3(new_n249), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n407), .A2(new_n409), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n258), .ZN(new_n413));
  AND3_X1   g0213(.A1(KEYINPUT65), .A2(G33), .A3(G41), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n414), .A2(new_n273), .A3(new_n217), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n272), .A2(G274), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT71), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT71), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n264), .A2(new_n267), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n417), .A2(new_n419), .B1(G238), .B2(new_n275), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n413), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g0221(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n413), .A2(new_n420), .A3(new_n422), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(KEYINPUT73), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT73), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n421), .A2(new_n427), .A3(new_n423), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G200), .ZN(new_n430));
  INV_X1    g0230(.A(new_n425), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n413), .B2(new_n420), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n431), .A2(new_n327), .A3(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n291), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n251), .B2(new_n289), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n287), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT11), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n298), .A2(new_n202), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT12), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n287), .A2(new_n436), .A3(KEYINPUT11), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n386), .A2(G68), .A3(new_n301), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n439), .A2(new_n441), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT74), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n434), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n430), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT76), .B(KEYINPUT14), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n429), .A2(KEYINPUT77), .A3(G169), .A4(new_n449), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n431), .A2(new_n315), .A3(new_n433), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n426), .A2(G169), .A3(new_n428), .A4(new_n449), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT77), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n426), .A2(G169), .A3(new_n428), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n455), .A2(KEYINPUT75), .A3(KEYINPUT14), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT75), .B1(new_n455), .B2(KEYINPUT14), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n450), .B(new_n454), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n448), .B1(new_n458), .B2(new_n445), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n405), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n283), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n391), .B1(new_n352), .B2(new_n343), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n292), .A2(new_n251), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g0265(.A(G97), .B(G107), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT6), .ZN(new_n467));
  INV_X1    g0267(.A(G97), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n466), .A2(new_n467), .B1(new_n391), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n465), .B1(new_n470), .B2(new_n209), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n463), .B1(new_n471), .B2(KEYINPUT82), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT82), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n473), .B(new_n465), .C1(new_n470), .C2(new_n209), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n462), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n298), .A2(new_n468), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n208), .A2(G33), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n299), .A2(new_n284), .A3(new_n286), .A4(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n478), .B2(new_n468), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT83), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(G97), .A2(G107), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n467), .B1(new_n481), .B2(new_n205), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n391), .A2(KEYINPUT6), .A3(G97), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n209), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT82), .B1(new_n484), .B2(new_n464), .ZN(new_n485));
  OAI21_X1  g0285(.A(G107), .B1(new_n342), .B2(new_n344), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n474), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n283), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT83), .ZN(new_n489));
  INV_X1    g0289(.A(new_n479), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n271), .A2(G1), .ZN(new_n492));
  NOR2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  AND2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n492), .B(G274), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT84), .B1(new_n415), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT84), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n208), .A2(G45), .A3(G274), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  XNOR2_X1  g0299(.A(KEYINPUT5), .B(G41), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n264), .A2(new_n497), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n263), .A2(new_n274), .B1(new_n500), .B2(new_n492), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n496), .A2(new_n501), .B1(new_n502), .B2(G257), .ZN(new_n503));
  OAI211_X1 g0303(.A(G250), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(new_n249), .C1(new_n339), .C2(new_n340), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n504), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n506), .A2(new_n507), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n258), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n503), .A2(G190), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G200), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n503), .B2(new_n510), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n480), .A2(new_n491), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n373), .B1(new_n503), .B2(new_n510), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n503), .A2(G179), .A3(new_n510), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n488), .A2(new_n490), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(G257), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n523));
  OAI211_X1 g0323(.A(G250), .B(new_n249), .C1(new_n339), .C2(new_n340), .ZN(new_n524));
  INV_X1    g0324(.A(G294), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(new_n245), .C2(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(new_n258), .B1(new_n502), .B2(G264), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n496), .A2(new_n501), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n315), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n373), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G116), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(G20), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n209), .B2(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n391), .A2(KEYINPUT23), .A3(G20), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT22), .ZN(new_n538));
  AOI21_X1  g0338(.A(G20), .B1(new_n246), .B2(new_n247), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(G87), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n209), .B(G87), .C1(new_n339), .C2(new_n340), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(KEYINPUT22), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n537), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT24), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n541), .A2(KEYINPUT22), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n248), .A2(new_n538), .A3(new_n209), .A4(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT24), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(new_n537), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n462), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n478), .A2(new_n391), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n298), .A2(new_n391), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT25), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n529), .B(new_n531), .C1(new_n550), .C2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n547), .A2(new_n548), .A3(new_n537), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n548), .B1(new_n547), .B2(new_n537), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n283), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n527), .A2(new_n327), .A3(new_n528), .ZN(new_n560));
  AOI21_X1  g0360(.A(G200), .B1(new_n527), .B2(new_n528), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n559), .B(new_n554), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n248), .A2(new_n209), .A3(G68), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n209), .B1(new_n410), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(G87), .B2(new_n206), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n564), .B1(new_n289), .B2(new_n468), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT85), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT85), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n563), .A2(new_n566), .A3(new_n570), .A4(new_n567), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n283), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n478), .ZN(new_n573));
  INV_X1    g0373(.A(new_n383), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n383), .A2(new_n298), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n572), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n248), .A2(G238), .A3(new_n249), .ZN(new_n578));
  INV_X1    g0378(.A(G244), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n532), .C1(new_n252), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n258), .ZN(new_n581));
  INV_X1    g0381(.A(G250), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n498), .B1(new_n492), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n264), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n373), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n580), .A2(new_n258), .B1(new_n264), .B2(new_n583), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n315), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n577), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n585), .A2(G200), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n462), .B1(new_n568), .B2(KEYINPUT85), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n591), .A2(new_n571), .B1(new_n298), .B2(new_n383), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n573), .A2(G87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n587), .A2(G190), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n590), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n556), .A2(new_n562), .A3(new_n589), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n502), .A2(G270), .ZN(new_n597));
  OAI211_X1 g0397(.A(G264), .B(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n598));
  OAI211_X1 g0398(.A(G257), .B(new_n249), .C1(new_n339), .C2(new_n340), .ZN(new_n599));
  INV_X1    g0399(.A(G303), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(new_n248), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n258), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n528), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G200), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n505), .B(new_n209), .C1(G33), .C2(new_n468), .ZN(new_n605));
  INV_X1    g0405(.A(G116), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G20), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n283), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT20), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n605), .A2(KEYINPUT20), .A3(new_n283), .A4(new_n607), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n607), .A2(G1), .A3(new_n297), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n606), .B1(new_n208), .B2(G33), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n386), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n604), .B(new_n617), .C1(new_n327), .C2(new_n603), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n528), .A2(new_n597), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n315), .B1(new_n601), .B2(new_n258), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT21), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n373), .B1(new_n612), .B2(new_n615), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(new_n603), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n603), .A2(new_n623), .A3(new_n622), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n618), .B(new_n621), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n522), .A2(new_n596), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n461), .A2(new_n627), .ZN(G372));
  NAND2_X1  g0428(.A1(new_n458), .A2(new_n445), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n448), .B2(new_n403), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n361), .A2(new_n365), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT89), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n380), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n376), .A2(new_n379), .A3(KEYINPUT89), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n312), .B(new_n314), .C1(new_n632), .C2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n556), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n621), .B1(new_n625), .B2(new_n624), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT86), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n581), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n580), .A2(KEYINPUT86), .A3(new_n258), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n584), .B(KEYINPUT87), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G200), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n647), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n577), .A2(new_n588), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n646), .A2(new_n373), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n562), .ZN(new_n653));
  NOR4_X1   g0453(.A1(new_n522), .A2(new_n641), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n648), .A2(new_n651), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT88), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n519), .B(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n489), .B1(new_n488), .B2(new_n490), .ZN(new_n659));
  AOI211_X1 g0459(.A(KEYINPUT83), .B(new_n479), .C1(new_n487), .C2(new_n283), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n655), .A2(new_n657), .A3(new_n658), .A4(new_n662), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n517), .A2(new_n518), .B1(new_n488), .B2(new_n490), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(new_n589), .A3(new_n595), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n651), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n461), .B1(new_n654), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n638), .A2(new_n668), .A3(new_n317), .ZN(G369));
  NOR2_X1   g0469(.A1(new_n297), .A2(G1), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n209), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT27), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n672), .A2(KEYINPUT90), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT90), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n671), .B2(KEYINPUT27), .ZN(new_n676));
  OAI221_X1 g0476(.A(G213), .B1(KEYINPUT27), .B2(new_n671), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n617), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT91), .ZN(new_n681));
  INV_X1    g0481(.A(new_n618), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n640), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n640), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n681), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n639), .A2(new_n653), .ZN(new_n689));
  INV_X1    g0489(.A(new_n679), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n550), .B2(new_n555), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n556), .B2(new_n679), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n685), .A2(new_n690), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n689), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n639), .B2(new_n679), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n212), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n208), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n702), .A2(new_n703), .B1(new_n216), .B2(new_n701), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  AND2_X1   g0505(.A1(new_n587), .A2(new_n527), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n503), .A2(new_n510), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n706), .A2(new_n708), .A3(new_n619), .A4(new_n620), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(G179), .B1(new_n527), .B2(new_n528), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n646), .A2(new_n707), .A3(new_n603), .A4(new_n712), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n619), .A2(new_n620), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(KEYINPUT30), .A3(new_n708), .A4(new_n706), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n711), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n716), .B2(new_n690), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT92), .B1(new_n627), .B2(new_n679), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n664), .B1(new_n661), .B2(new_n514), .ZN(new_n721));
  AND4_X1   g0521(.A1(new_n556), .A2(new_n562), .A3(new_n589), .A4(new_n595), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n721), .A2(new_n722), .A3(new_n683), .A4(new_n679), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT92), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n719), .B1(new_n720), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n679), .B1(new_n667), .B2(new_n654), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n657), .A2(new_n662), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT26), .B1(new_n732), .B2(new_n652), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n651), .B(KEYINPUT93), .Z(new_n734));
  OAI211_X1 g0534(.A(new_n733), .B(new_n734), .C1(KEYINPUT26), .C2(new_n665), .ZN(new_n735));
  OAI211_X1 g0535(.A(KEYINPUT29), .B(new_n679), .C1(new_n735), .C2(new_n654), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n728), .B1(new_n731), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n705), .B1(new_n737), .B2(G1), .ZN(G364));
  NOR2_X1   g0538(.A1(new_n297), .A2(G20), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT94), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G45), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n702), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n688), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G330), .B2(new_n686), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n212), .A2(new_n248), .ZN(new_n746));
  INV_X1    g0546(.A(G355), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n746), .A2(new_n747), .B1(G116), .B2(new_n212), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n700), .A2(new_n248), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n271), .B2(new_n216), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n239), .A2(new_n271), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n217), .B1(G20), .B2(new_n373), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n743), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n327), .A2(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n209), .B1(new_n761), .B2(new_n315), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n209), .A2(G179), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n762), .A2(new_n525), .B1(new_n764), .B2(new_n600), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n209), .A2(new_n315), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G190), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(KEYINPUT33), .B(G317), .Z(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n767), .A2(new_n327), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n765), .B(new_n771), .C1(G326), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G190), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n763), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n248), .B1(new_n776), .B2(G329), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n763), .A2(new_n327), .A3(G200), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n766), .B(KEYINPUT95), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n761), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n780), .B1(new_n783), .B2(G322), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n781), .A2(new_n774), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n773), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n786), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G58), .A2(new_n783), .B1(new_n788), .B2(G77), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n762), .A2(new_n468), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G50), .B2(new_n772), .ZN(new_n791));
  INV_X1    g0591(.A(G159), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n775), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT32), .ZN(new_n794));
  INV_X1    g0594(.A(G87), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n764), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n248), .B1(new_n779), .B2(new_n391), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(G68), .C2(new_n768), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n789), .A2(new_n791), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n787), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n760), .B1(new_n800), .B2(new_n757), .ZN(new_n801));
  INV_X1    g0601(.A(new_n756), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n686), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n745), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NAND2_X1  g0605(.A1(new_n690), .A2(new_n389), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n400), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n403), .ZN(new_n808));
  INV_X1    g0608(.A(new_n403), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n679), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n729), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n811), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n679), .B(new_n813), .C1(new_n667), .C2(new_n654), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n743), .B1(new_n815), .B2(new_n727), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n727), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n757), .A2(new_n754), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n742), .B1(new_n251), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n757), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n248), .B(new_n790), .C1(G311), .C2(new_n776), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n821), .B1(new_n606), .B2(new_n786), .C1(new_n525), .C2(new_n782), .ZN(new_n822));
  INV_X1    g0622(.A(new_n772), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n823), .A2(new_n600), .B1(new_n779), .B2(new_n795), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n769), .A2(new_n778), .B1(new_n764), .B2(new_n391), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G50), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n762), .A2(new_n201), .B1(new_n764), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n248), .B1(new_n775), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT96), .ZN(new_n831));
  INV_X1    g0631(.A(new_n779), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n828), .B(new_n831), .C1(G68), .C2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT97), .Z(new_n834));
  AOI22_X1  g0634(.A1(G137), .A2(new_n772), .B1(new_n768), .B2(G150), .ZN(new_n835));
  INV_X1    g0635(.A(G143), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n835), .B1(new_n786), .B2(new_n792), .C1(new_n836), .C2(new_n782), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n826), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n819), .B1(new_n820), .B2(new_n839), .C1(new_n813), .C2(new_n755), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n817), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G384));
  NAND2_X1  g0642(.A1(new_n216), .A2(G77), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n331), .A2(new_n333), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n843), .A2(new_n844), .B1(G50), .B2(new_n202), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(G1), .A3(new_n297), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT98), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT36), .ZN(new_n848));
  INV_X1    g0648(.A(new_n470), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n849), .A2(KEYINPUT35), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(KEYINPUT35), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n850), .A2(new_n851), .A3(G116), .A4(new_n218), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n847), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n848), .B2(new_n852), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT99), .Z(new_n855));
  INV_X1    g0655(.A(new_n445), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(new_n679), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n459), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n629), .B2(new_n679), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n814), .A2(new_n810), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT100), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT100), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n338), .A2(new_n347), .A3(new_n345), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n349), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(new_n287), .A3(new_n348), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n677), .B1(new_n869), .B2(new_n359), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n631), .B2(new_n380), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n360), .A2(KEYINPUT37), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n873), .A2(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n869), .A2(new_n359), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n377), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n377), .A2(new_n378), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n378), .A2(new_n678), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(new_n360), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n866), .B1(new_n872), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n870), .B1(new_n381), .B2(new_n366), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n874), .A2(new_n876), .B1(new_n880), .B2(new_n881), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n864), .A2(new_n865), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n637), .A2(new_n677), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n879), .A2(new_n360), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n363), .A2(new_n375), .ZN(new_n892));
  NOR4_X1   g0692(.A1(new_n891), .A2(new_n892), .A3(new_n633), .A4(new_n881), .ZN(new_n893));
  INV_X1    g0693(.A(new_n891), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n879), .A2(new_n633), .A3(new_n360), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n894), .A2(new_n878), .B1(new_n895), .B2(KEYINPUT37), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n634), .A2(new_n631), .A3(new_n635), .ZN(new_n897));
  INV_X1    g0697(.A(new_n879), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n893), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n887), .B1(new_n899), .B2(KEYINPUT38), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n450), .A2(new_n454), .ZN(new_n903));
  INV_X1    g0703(.A(new_n457), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n455), .A2(KEYINPUT75), .A3(KEYINPUT14), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n856), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n902), .A2(new_n907), .A3(new_n679), .A4(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n889), .A2(new_n890), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n461), .A2(new_n731), .A3(new_n736), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n638), .A2(new_n317), .A3(new_n911), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n910), .B(new_n912), .Z(new_n913));
  NAND2_X1  g0713(.A1(new_n723), .A2(new_n724), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n596), .A2(new_n626), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n915), .A2(KEYINPUT92), .A3(new_n721), .A4(new_n679), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n811), .B1(new_n917), .B2(new_n719), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n900), .A2(new_n860), .A3(KEYINPUT40), .A4(new_n918), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n857), .B(new_n448), .C1(new_n458), .C2(new_n445), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n629), .A2(new_n679), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n918), .B(new_n888), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n461), .A2(new_n726), .ZN(new_n926));
  OAI21_X1  g0726(.A(G330), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n925), .B2(new_n926), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n913), .A2(new_n928), .B1(new_n208), .B2(new_n740), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n913), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n855), .B1(new_n929), .B2(new_n930), .ZN(G367));
  OAI21_X1  g0731(.A(new_n721), .B1(new_n661), .B2(new_n679), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n732), .B2(new_n679), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n697), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT42), .Z(new_n935));
  AND2_X1   g0735(.A1(new_n933), .A2(new_n639), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n679), .B1(new_n936), .B2(new_n664), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n592), .A2(new_n593), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n690), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT101), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(new_n649), .A3(new_n650), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n652), .B2(new_n940), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n935), .A2(new_n937), .B1(KEYINPUT43), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n943), .B(new_n944), .Z(new_n945));
  NAND3_X1  g0745(.A1(new_n688), .A2(new_n693), .A3(new_n933), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT102), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n945), .A2(new_n946), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n741), .A2(G1), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n701), .B(KEYINPUT41), .Z(new_n953));
  NAND2_X1  g0753(.A1(new_n698), .A2(new_n933), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT45), .Z(new_n955));
  NOR2_X1   g0755(.A1(new_n698), .A2(new_n933), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(new_n694), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n688), .A2(KEYINPUT103), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n687), .B(KEYINPUT103), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n696), .B1(new_n693), .B2(new_n695), .ZN(new_n962));
  MUX2_X1   g0762(.A(new_n960), .B(new_n961), .S(new_n962), .Z(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n737), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n959), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n953), .B1(new_n966), .B2(new_n737), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n951), .B1(new_n948), .B2(new_n947), .C1(new_n952), .C2(new_n967), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n758), .B1(new_n212), .B2(new_n383), .C1(new_n750), .C2(new_n235), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n969), .A2(new_n743), .ZN(new_n970));
  INV_X1    g0770(.A(G137), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n248), .B1(new_n775), .B2(new_n971), .C1(new_n251), .C2(new_n779), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n783), .B2(G150), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n827), .B2(new_n786), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n762), .A2(new_n202), .B1(new_n764), .B2(new_n201), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n769), .A2(new_n792), .B1(new_n823), .B2(new_n836), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT107), .Z(new_n978));
  NOR2_X1   g0778(.A1(new_n764), .A2(new_n606), .ZN(new_n979));
  AOI22_X1  g0779(.A1(KEYINPUT46), .A2(new_n979), .B1(new_n768), .B2(G294), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(KEYINPUT46), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT104), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n981), .A2(new_n982), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n980), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT105), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(KEYINPUT105), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n778), .A2(new_n786), .B1(new_n782), .B2(new_n600), .ZN(new_n989));
  XNOR2_X1  g0789(.A(KEYINPUT106), .B(G317), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n341), .B1(new_n775), .B2(new_n990), .C1(new_n762), .C2(new_n391), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n823), .A2(new_n785), .B1(new_n779), .B2(new_n468), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n987), .A2(new_n988), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n978), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT47), .Z(new_n996));
  OAI221_X1 g0796(.A(new_n970), .B1(new_n802), .B2(new_n942), .C1(new_n996), .C2(new_n820), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n968), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT108), .ZN(G387));
  OR2_X1    g0799(.A1(new_n693), .A2(new_n802), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G311), .A2(new_n768), .B1(new_n772), .B2(G322), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n786), .B2(new_n600), .C1(new_n782), .C2(new_n990), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT48), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n762), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n764), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1006), .A2(G283), .B1(new_n1007), .B2(G294), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n779), .A2(new_n606), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n248), .B(new_n1013), .C1(G326), .C2(new_n776), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n762), .A2(new_n383), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n823), .A2(new_n792), .B1(new_n764), .B2(new_n251), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n356), .C2(new_n768), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n248), .B1(new_n775), .B2(new_n290), .C1(new_n468), .C2(new_n779), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n783), .B2(G50), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(new_n202), .C2(new_n786), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n820), .B1(new_n1015), .B2(new_n1021), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n746), .A2(new_n703), .B1(G107), .B2(new_n212), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n232), .A2(new_n271), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT109), .Z(new_n1025));
  INV_X1    g0825(.A(new_n703), .ZN(new_n1026));
  AOI211_X1 g0826(.A(G45), .B(new_n1026), .C1(G68), .C2(G77), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n288), .A2(G50), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT50), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n750), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1023), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n743), .B1(new_n1031), .B2(new_n759), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1022), .A2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n963), .A2(new_n952), .B1(new_n1000), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n964), .A2(new_n701), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n963), .A2(new_n737), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(G393));
  NOR2_X1   g0837(.A1(new_n933), .A2(new_n802), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT110), .Z(new_n1039));
  OAI21_X1  g0839(.A(new_n758), .B1(new_n468), .B2(new_n212), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n749), .B2(new_n242), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n782), .A2(new_n792), .B1(new_n290), .B2(new_n823), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT51), .Z(new_n1043));
  AOI22_X1  g0843(.A1(new_n768), .A2(G50), .B1(new_n1006), .B2(G77), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n202), .B2(new_n764), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n786), .A2(new_n288), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n248), .B1(new_n775), .B2(new_n836), .C1(new_n795), .C2(new_n779), .ZN(new_n1047));
  NOR4_X1   g0847(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1048), .A2(KEYINPUT111), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(KEYINPUT111), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n783), .A2(G311), .B1(G317), .B2(new_n772), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT52), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n764), .A2(new_n778), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n769), .A2(new_n600), .B1(new_n606), .B2(new_n762), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n248), .B1(new_n776), .B2(G322), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n391), .B2(new_n779), .C1(new_n786), .C2(new_n525), .ZN(new_n1056));
  OR4_X1    g0856(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1049), .A2(new_n1050), .A3(new_n1057), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n742), .B(new_n1041), .C1(new_n1058), .C2(new_n757), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n959), .A2(new_n952), .B1(new_n1039), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n966), .A2(new_n701), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n959), .A2(new_n965), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(G390));
  INV_X1    g0863(.A(new_n818), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n743), .B1(new_n356), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n248), .B(new_n796), .C1(G294), .C2(new_n776), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n468), .B2(new_n786), .C1(new_n606), .C2(new_n782), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1006), .A2(G77), .B1(new_n832), .B2(G68), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n391), .B2(new_n769), .C1(new_n778), .C2(new_n823), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n779), .A2(new_n827), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n341), .B(new_n1070), .C1(G125), .C2(new_n776), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(KEYINPUT54), .B(G143), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1071), .B1(new_n786), .B2(new_n1072), .C1(new_n829), .C2(new_n782), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n764), .A2(new_n290), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT53), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n772), .A2(G128), .B1(new_n1006), .B2(G159), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n971), .C2(new_n769), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1067), .A2(new_n1069), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1065), .B1(new_n1078), .B2(new_n757), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n902), .A2(new_n908), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1079), .B1(new_n1081), .B2(new_n755), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n907), .A2(new_n679), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n862), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n860), .A2(G330), .A3(new_n918), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n679), .B(new_n808), .C1(new_n735), .C2(new_n654), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n810), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n860), .A2(KEYINPUT112), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n459), .A2(new_n858), .B1(new_n907), .B2(new_n690), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT112), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1089), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n900), .A2(new_n1083), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1085), .B(new_n1086), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1086), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1098), .B2(new_n1088), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n902), .A2(new_n908), .B1(new_n862), .B2(new_n1083), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n952), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1082), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n460), .A2(new_n727), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT113), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(new_n912), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1089), .A2(new_n1086), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1098), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n728), .A2(KEYINPUT114), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT114), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n727), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1111), .A2(new_n813), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1109), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n726), .A2(new_n813), .ZN(new_n1116));
  INV_X1    g0916(.A(G330), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1091), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1086), .A2(new_n1118), .B1(new_n810), .B2(new_n814), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1108), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1102), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n701), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n1102), .B2(new_n1120), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1104), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(G378));
  NOR2_X1   g0925(.A1(new_n306), .A2(new_n677), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n318), .B(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1127), .B(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT117), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n919), .A2(new_n924), .A3(new_n1130), .A4(G330), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1091), .A2(new_n1116), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n897), .A2(new_n898), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n896), .A2(new_n893), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n866), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n923), .B1(new_n1137), .B2(new_n887), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1117), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1130), .B1(new_n1139), .B2(new_n924), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1129), .B1(new_n1132), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n910), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n919), .A2(new_n924), .A3(G330), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1129), .B1(new_n1143), .B2(KEYINPUT117), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1141), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1129), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n922), .A2(new_n923), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT38), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n887), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT40), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(G330), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(KEYINPUT117), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1147), .B1(new_n1154), .B2(new_n1131), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n910), .B1(new_n1155), .B2(new_n1144), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1146), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n952), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n341), .A2(new_n270), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G283), .B2(new_n776), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n202), .B2(new_n762), .C1(new_n782), .C2(new_n391), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n768), .A2(G97), .B1(new_n1007), .B2(G77), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n201), .B2(new_n779), .C1(new_n606), .C2(new_n823), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(new_n574), .C2(new_n788), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT115), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(KEYINPUT58), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1159), .B(new_n827), .C1(G33), .C2(G41), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G128), .A2(new_n783), .B1(new_n788), .B2(G137), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n772), .A2(G125), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n768), .A2(G132), .B1(new_n1006), .B2(G150), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n764), .A2(new_n1072), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT116), .Z(new_n1173));
  NOR2_X1   g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n832), .A2(G159), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G33), .B(G41), .C1(new_n776), .C2(G124), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1165), .A2(KEYINPUT58), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1166), .A2(new_n1167), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n757), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n742), .B1(new_n827), .B2(new_n818), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n1147), .C2(new_n755), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1158), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1108), .B1(new_n1102), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1157), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT57), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1122), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT118), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1146), .B2(new_n1156), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT118), .B1(new_n1196), .B2(new_n910), .ZN(new_n1197));
  OAI211_X1 g0997(.A(KEYINPUT57), .B(new_n1189), .C1(new_n1195), .C2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1187), .B1(new_n1193), .B2(new_n1199), .ZN(G375));
  OAI21_X1  g1000(.A(new_n952), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT121), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n742), .B1(new_n202), .B2(new_n818), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n769), .A2(new_n606), .B1(new_n823), .B2(new_n525), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1016), .B(new_n1204), .C1(G97), .C2(new_n1007), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n341), .B1(new_n775), .B2(new_n600), .C1(new_n251), .C2(new_n779), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n788), .B2(G107), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(new_n778), .C2(new_n782), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT119), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n248), .B1(new_n201), .B2(new_n779), .C1(new_n782), .C2(new_n971), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G150), .B2(new_n788), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1007), .A2(G159), .B1(new_n776), .B2(G128), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT120), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n829), .A2(new_n823), .B1(new_n769), .B2(new_n1072), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G50), .B2(new_n1006), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1212), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1210), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1203), .B1(new_n820), .B2(new_n1219), .C1(new_n1098), .C2(new_n755), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1201), .A2(new_n1202), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1202), .B1(new_n1201), .B2(new_n1220), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1108), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1188), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n953), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n1120), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1224), .A2(new_n1228), .ZN(G381));
  OR2_X1    g1029(.A1(G375), .A2(G378), .ZN(new_n1230));
  OR4_X1    g1030(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1231));
  OR4_X1    g1031(.A1(G387), .A2(G381), .A3(new_n1230), .A4(new_n1231), .ZN(G407));
  OAI211_X1 g1032(.A(G407), .B(G213), .C1(G343), .C2(new_n1230), .ZN(G409));
  AOI211_X1 g1033(.A(new_n1124), .B(new_n1186), .C1(new_n1192), .C2(new_n1198), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT122), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1142), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1155), .A2(new_n910), .A3(new_n1144), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT118), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1156), .A2(new_n1194), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1103), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1185), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1235), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1190), .A2(new_n953), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n952), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(KEYINPUT122), .A3(new_n1185), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1242), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1234), .B1(new_n1124), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(G213), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(G343), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT124), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT124), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1250), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1241), .B1(new_n1254), .B2(new_n952), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1243), .B1(new_n1255), .B2(KEYINPUT122), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G378), .B1(new_n1256), .B2(new_n1242), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1252), .B(new_n1253), .C1(new_n1257), .C2(new_n1234), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1226), .A2(KEYINPUT123), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1226), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1120), .A2(new_n701), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G384), .B(new_n1224), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n841), .B1(new_n1266), .B2(new_n1223), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1251), .A2(new_n1258), .A3(KEYINPUT62), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1246), .A2(new_n1244), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT122), .B1(new_n1245), .B2(new_n1185), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1124), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G378), .B(new_n1187), .C1(new_n1193), .C2(new_n1199), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1250), .B(new_n1268), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(KEYINPUT125), .B1(new_n1275), .B2(KEYINPUT62), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT125), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1253), .B1(new_n1257), .B2(new_n1234), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1277), .B(new_n1278), .C1(new_n1279), .C2(new_n1268), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1270), .A2(new_n1276), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1251), .A2(new_n1258), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1250), .A2(G2897), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1268), .B(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G393), .B(new_n804), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(G390), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1288), .A2(KEYINPUT108), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n998), .B(new_n1289), .C1(G390), .C2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1289), .B1(new_n1290), .B2(G390), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n997), .A3(new_n968), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT126), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1294), .B(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1286), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1291), .A2(new_n1293), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(new_n1284), .B2(new_n1279), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1275), .A2(KEYINPUT63), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1251), .A2(new_n1258), .A3(KEYINPUT63), .A4(new_n1269), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1298), .A2(KEYINPUT127), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1296), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1304), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1306), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1309), .ZN(G405));
  NAND2_X1  g1110(.A1(G375), .A2(new_n1124), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1274), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1312), .B(new_n1268), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1296), .B(new_n1313), .ZN(G402));
endmodule


