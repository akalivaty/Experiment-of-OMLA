//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT0), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G57gat), .ZN(new_n205));
  INV_X1    g004(.A(G85gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G225gat), .A2(G233gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G120gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G113gat), .ZN(new_n212));
  INV_X1    g011(.A(G113gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G120gat), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT1), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G127gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G113gat), .B(G120gat), .ZN(new_n218));
  OAI21_X1  g017(.A(G127gat), .B1(new_n218), .B2(KEYINPUT1), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n219), .A3(G134gat), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G148gat), .ZN(new_n222));
  INV_X1    g021(.A(G148gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G141gat), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT75), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT2), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(G141gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n221), .A2(G148gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n225), .A2(new_n226), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n233), .B(KEYINPUT74), .Z(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G134gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n215), .A2(new_n216), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n218), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G162gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT76), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT76), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G162gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G155gat), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT2), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n228), .ZN(new_n247));
  INV_X1    g046(.A(new_n232), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n246), .B(new_n247), .C1(new_n233), .C2(new_n248), .ZN(new_n249));
  AND4_X1   g048(.A1(new_n220), .A2(new_n235), .A3(new_n239), .A4(new_n249), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n249), .A2(new_n235), .B1(new_n239), .B2(new_n220), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n210), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n249), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n220), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n235), .A2(new_n249), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n209), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT77), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n235), .A2(new_n239), .A3(new_n249), .A4(new_n220), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(new_n263), .B2(KEYINPUT4), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n235), .A2(new_n249), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n217), .A2(new_n219), .A3(G134gat), .ZN(new_n266));
  AOI21_X1  g065(.A(G134gat), .B1(new_n217), .B2(new_n219), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n265), .A2(KEYINPUT77), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n263), .A2(KEYINPUT4), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n264), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n253), .B1(new_n261), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n274), .A3(new_n209), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT78), .B1(new_n263), .B2(KEYINPUT4), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n276), .A2(new_n271), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT78), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n265), .A2(new_n278), .A3(new_n268), .A4(new_n269), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n208), .B1(new_n273), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n254), .A2(new_n256), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n263), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n274), .B1(new_n283), .B2(new_n210), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n264), .A2(new_n270), .A3(new_n271), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n284), .B1(new_n285), .B2(new_n260), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n276), .A2(new_n279), .A3(new_n271), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n261), .A2(new_n274), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n207), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n281), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI211_X1 g090(.A(KEYINPUT6), .B(new_n208), .C1(new_n273), .C2(new_n280), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n296), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  NOR3_X1   g098(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n294), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT64), .ZN(new_n306));
  INV_X1    g105(.A(G183gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(KEYINPUT27), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n305), .B(new_n308), .C1(new_n309), .C2(new_n306), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(KEYINPUT28), .A3(new_n305), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n295), .A2(new_n297), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT65), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(KEYINPUT66), .B(new_n302), .C1(new_n318), .C2(new_n300), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n314), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G169gat), .ZN(new_n321));
  INV_X1    g120(.A(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT23), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT24), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n303), .A2(new_n325), .B1(G169gat), .B2(G176gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n307), .A2(new_n305), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(KEYINPUT24), .A3(new_n302), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT25), .A4(new_n328), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n320), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT70), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G218gat), .ZN(new_n344));
  INV_X1    g143(.A(G197gat), .ZN(new_n345));
  INV_X1    g144(.A(G204gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G197gat), .A2(G204gat), .ZN(new_n348));
  OR2_X1    g147(.A1(KEYINPUT69), .A2(G211gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(KEYINPUT69), .A2(G211gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(G218gat), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT22), .ZN(new_n352));
  AOI221_X4 g151(.A(G211gat), .B1(new_n347), .B2(new_n348), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G211gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n352), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n347), .A2(new_n348), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n344), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(KEYINPUT69), .A2(G211gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(KEYINPUT69), .A2(G211gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT22), .B1(new_n361), .B2(G218gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n356), .ZN(new_n363));
  OAI21_X1  g162(.A(G211gat), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n355), .A2(new_n354), .A3(new_n356), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(G218gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n334), .A2(KEYINPUT72), .A3(new_n340), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n339), .A2(new_n343), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT73), .ZN(new_n370));
  INV_X1    g169(.A(new_n338), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n334), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT29), .B1(new_n320), .B2(new_n333), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n340), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n367), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT72), .B1(new_n334), .B2(new_n340), .ZN(new_n377));
  INV_X1    g176(.A(new_n340), .ZN(new_n378));
  AOI211_X1 g177(.A(new_n342), .B(new_n378), .C1(new_n320), .C2(new_n333), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT73), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n367), .A4(new_n339), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n370), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G8gat), .B(G36gat), .Z(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(G64gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n385), .B(G92gat), .Z(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n386), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n370), .A2(new_n376), .A3(new_n382), .A4(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(KEYINPUT30), .A3(new_n389), .ZN(new_n390));
  OR3_X1    g189(.A1(new_n383), .A2(KEYINPUT30), .A3(new_n386), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n293), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT31), .ZN(new_n394));
  INV_X1    g193(.A(G50gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n358), .B2(new_n366), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n254), .B1(new_n397), .B2(KEYINPUT3), .ZN(new_n398));
  NAND2_X1  g197(.A1(G228gat), .A2(G233gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n258), .A2(new_n335), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n375), .A2(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n398), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n398), .B2(new_n402), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n403), .A2(new_n404), .A3(G22gat), .ZN(new_n405));
  INV_X1    g204(.A(G22gat), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n353), .A2(new_n357), .A3(new_n344), .ZN(new_n407));
  AOI21_X1  g206(.A(G218gat), .B1(new_n364), .B2(new_n365), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n335), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n265), .B1(new_n409), .B2(new_n257), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n367), .B1(new_n335), .B2(new_n258), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n399), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n398), .A2(new_n400), .A3(new_n402), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n406), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n396), .B1(new_n405), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(KEYINPUT79), .ZN(new_n416));
  OAI21_X1  g215(.A(G22gat), .B1(new_n403), .B2(new_n404), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n406), .A3(new_n413), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n396), .A2(KEYINPUT79), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT80), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n415), .A2(new_n423), .A3(new_n416), .A4(new_n420), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n334), .A2(new_n256), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n320), .A2(new_n268), .A3(new_n333), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G227gat), .ZN(new_n430));
  INV_X1    g229(.A(G233gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n426), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n432), .ZN(new_n434));
  INV_X1    g233(.A(new_n426), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n427), .A2(new_n434), .A3(new_n428), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G15gat), .B(G43gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G71gat), .ZN(new_n439));
  INV_X1    g238(.A(G99gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n434), .B1(new_n427), .B2(new_n428), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(KEYINPUT33), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT32), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  AOI221_X4 g245(.A(new_n444), .B1(KEYINPUT33), .B2(new_n441), .C1(new_n429), .C2(new_n432), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n437), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n448), .A2(KEYINPUT68), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n443), .A2(new_n445), .ZN(new_n450));
  INV_X1    g249(.A(new_n437), .ZN(new_n451));
  INV_X1    g250(.A(new_n447), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n448), .A3(KEYINPUT68), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n392), .A2(new_n425), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n448), .ZN(new_n457));
  AOI211_X1 g256(.A(new_n202), .B(new_n457), .C1(new_n422), .C2(new_n424), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n202), .A2(new_n456), .B1(new_n458), .B2(new_n392), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n453), .A2(new_n448), .A3(KEYINPUT36), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n455), .B2(KEYINPUT36), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n388), .A2(KEYINPUT38), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT37), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n374), .B2(new_n367), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n339), .A2(new_n343), .A3(new_n375), .A4(new_n368), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n465), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n370), .A2(new_n464), .A3(new_n376), .A4(new_n382), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n462), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n465), .A2(new_n466), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT83), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n477), .A2(KEYINPUT84), .A3(new_n471), .A4(new_n463), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n473), .A2(new_n293), .A3(new_n478), .A4(new_n389), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n383), .A2(KEYINPUT37), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n471), .A2(new_n386), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT38), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n390), .A2(new_n391), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT40), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n287), .A2(new_n259), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT39), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n210), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n207), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n282), .A2(new_n209), .A3(new_n263), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT39), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT81), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT81), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(new_n494), .A3(KEYINPUT39), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n209), .B1(new_n287), .B2(new_n259), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n486), .B1(new_n490), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT82), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n487), .A2(new_n210), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(new_n493), .A3(new_n495), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n208), .B1(new_n497), .B2(new_n488), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(KEYINPUT40), .A3(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(KEYINPUT82), .B(new_n486), .C1(new_n490), .C2(new_n498), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n501), .A2(new_n281), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n425), .B1(new_n485), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n461), .B1(new_n484), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n392), .A2(new_n425), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n459), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT16), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n513), .B2(G1gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(G1gat), .B2(new_n512), .ZN(new_n515));
  INV_X1    g314(.A(G8gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G43gat), .B(G50gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(G29gat), .A2(G36gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n520));
  INV_X1    g319(.A(G29gat), .ZN(new_n521));
  INV_X1    g320(.A(G36gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n519), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n525), .A2(KEYINPUT85), .ZN(new_n529));
  OAI211_X1 g328(.A(KEYINPUT15), .B(new_n518), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT86), .ZN(new_n532));
  OAI22_X1  g331(.A1(new_n518), .A2(KEYINPUT15), .B1(KEYINPUT87), .B2(new_n523), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(KEYINPUT87), .B2(new_n526), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT88), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n517), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n530), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT17), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n539), .B2(new_n517), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n538), .B(new_n517), .Z(new_n545));
  XOR2_X1   g344(.A(new_n541), .B(KEYINPUT89), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT13), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n540), .A2(KEYINPUT18), .A3(new_n541), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n544), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G197gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT11), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(new_n321), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT12), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n544), .A2(new_n555), .A3(new_n548), .A4(new_n549), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(KEYINPUT90), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT90), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n550), .A2(new_n560), .A3(new_n556), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT104), .ZN(new_n564));
  NAND2_X1  g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  OR2_X1    g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n569), .A2(KEYINPUT91), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(KEYINPUT91), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT92), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n565), .B(new_n566), .C1(new_n569), .C2(new_n567), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT7), .ZN(new_n579));
  INV_X1    g378(.A(G106gat), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT8), .B1(new_n440), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT97), .B(G92gat), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n579), .B(new_n581), .C1(G85gat), .C2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G99gat), .B(G106gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT98), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n577), .A2(KEYINPUT10), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n575), .B(new_n585), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G230gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(new_n431), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n589), .A2(new_n595), .ZN(new_n597));
  XNOR2_X1  g396(.A(G120gat), .B(G148gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n322), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(new_n346), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n596), .B2(new_n597), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n564), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(KEYINPUT104), .A3(new_n602), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n563), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n575), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(KEYINPUT21), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT96), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT95), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n617), .A3(new_n517), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n617), .B1(new_n616), .B2(new_n517), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(new_n618), .A3(new_n614), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n612), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT93), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT19), .ZN(new_n628));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT20), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n628), .B(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n621), .A2(new_n623), .A3(new_n612), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n625), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n631), .ZN(new_n634));
  INV_X1    g433(.A(new_n632), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n634), .B1(new_n635), .B2(new_n624), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(G232gat), .A2(G233gat), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n539), .A2(new_n586), .B1(KEYINPUT41), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G190gat), .B(G218gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT99), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n587), .A2(new_n538), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n638), .A2(KEYINPUT41), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n639), .A2(new_n642), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(new_n641), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n645), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT103), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n643), .B(KEYINPUT100), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n645), .A2(KEYINPUT101), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n656), .A3(new_n650), .ZN(new_n657));
  INV_X1    g456(.A(new_n648), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT102), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(new_n661), .A3(new_n658), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n652), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n511), .A2(new_n609), .A3(new_n637), .A4(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n293), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  INV_X1    g467(.A(new_n485), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n513), .A2(new_n516), .ZN(new_n670));
  NAND2_X1  g469(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n666), .A2(new_n669), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n666), .ZN(new_n675));
  OAI21_X1  g474(.A(G8gat), .B1(new_n675), .B2(new_n485), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n672), .A2(KEYINPUT107), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT107), .B1(new_n672), .B2(new_n677), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n674), .B(new_n676), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT108), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n672), .A2(new_n677), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n678), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n686), .A2(new_n687), .A3(new_n674), .A4(new_n676), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n682), .A2(new_n688), .ZN(G1325gat));
  AOI21_X1  g488(.A(G15gat), .B1(new_n666), .B2(new_n455), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n461), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n691), .B2(G15gat), .ZN(G1326gat));
  OAI21_X1  g491(.A(KEYINPUT109), .B1(new_n675), .B2(new_n425), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n422), .A2(new_n424), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n666), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT43), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n693), .A2(new_n699), .A3(new_n696), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n698), .A2(G22gat), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(G22gat), .B1(new_n698), .B2(new_n700), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(G1327gat));
  XOR2_X1   g502(.A(new_n651), .B(KEYINPUT103), .Z(new_n704));
  AND3_X1   g503(.A1(new_n657), .A2(new_n661), .A3(new_n658), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n661), .B1(new_n657), .B2(new_n658), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n291), .A2(new_n292), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n485), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n695), .A3(KEYINPUT110), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n392), .B2(new_n425), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n459), .B1(new_n509), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n471), .B(new_n463), .C1(new_n469), .C2(new_n468), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n710), .B1(new_n719), .B2(new_n462), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n720), .A2(new_n389), .A3(new_n482), .A4(new_n478), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n506), .A2(new_n281), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n503), .A2(new_n504), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT82), .B1(new_n723), .B2(new_n486), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n725), .A2(new_n391), .A3(new_n390), .A4(new_n505), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n721), .A2(new_n425), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n727), .A2(new_n461), .A3(new_n714), .A4(new_n712), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(KEYINPUT111), .A3(new_n459), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n709), .B1(new_n718), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n708), .B1(new_n511), .B2(new_n707), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n637), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n609), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(KEYINPUT112), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(KEYINPUT112), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n710), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n511), .A2(new_n707), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n734), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n521), .A3(new_n293), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT45), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n739), .A2(new_n743), .ZN(G1328gat));
  OAI21_X1  g543(.A(G36gat), .B1(new_n738), .B2(new_n485), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n741), .A2(new_n522), .A3(new_n669), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT46), .Z(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1329gat));
  INV_X1    g547(.A(G43gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n741), .A2(new_n749), .A3(new_n455), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n732), .A2(new_n461), .A3(new_n734), .ZN(new_n751));
  OAI211_X1 g550(.A(KEYINPUT47), .B(new_n750), .C1(new_n751), .C2(new_n749), .ZN(new_n752));
  INV_X1    g551(.A(new_n750), .ZN(new_n753));
  INV_X1    g552(.A(new_n461), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n736), .B2(new_n737), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n753), .B1(new_n755), .B2(G43gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n752), .B1(new_n756), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n395), .A3(new_n695), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n732), .A2(new_n425), .A3(new_n734), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT48), .B(new_n758), .C1(new_n759), .C2(new_n395), .ZN(new_n760));
  INV_X1    g559(.A(new_n758), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n695), .B1(new_n736), .B2(new_n737), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(G50gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n760), .B1(new_n763), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g563(.A(new_n608), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n718), .B2(new_n729), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n707), .A2(new_n733), .A3(new_n562), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n293), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g570(.A1(new_n768), .A2(new_n485), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  AND2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n772), .B2(new_n773), .ZN(G1333gat));
  OAI21_X1  g575(.A(G71gat), .B1(new_n768), .B2(new_n461), .ZN(new_n777));
  INV_X1    g576(.A(new_n455), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n778), .A2(G71gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n768), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g580(.A1(new_n769), .A2(new_n695), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  INV_X1    g582(.A(new_n709), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n728), .A2(KEYINPUT111), .A3(new_n459), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT111), .B1(new_n728), .B2(new_n459), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n740), .A2(KEYINPUT44), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n637), .A2(new_n562), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n608), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT113), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  AOI211_X1 g593(.A(new_n794), .B(new_n791), .C1(new_n787), .C2(new_n788), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(KEYINPUT114), .A3(new_n293), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n796), .B2(new_n710), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(G85gat), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n716), .A2(new_n707), .A3(new_n790), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT115), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n802), .A2(new_n803), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n608), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n293), .A2(new_n206), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n801), .B1(new_n808), .B2(new_n809), .ZN(G1336gat));
  NOR3_X1   g609(.A1(new_n765), .A2(G92gat), .A3(new_n485), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n792), .B1(new_n730), .B2(new_n731), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n582), .B1(new_n814), .B2(new_n485), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n669), .B1(new_n793), .B2(new_n795), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT116), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n716), .A2(new_n819), .A3(new_n707), .A4(new_n790), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n803), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n818), .A2(KEYINPUT117), .A3(new_n803), .A4(new_n820), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n806), .A3(new_n824), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n817), .A2(new_n582), .B1(new_n811), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(KEYINPUT118), .A3(new_n813), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n811), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n794), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n789), .A2(KEYINPUT113), .A3(new_n792), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n485), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n582), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n828), .B1(new_n834), .B2(KEYINPUT52), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n816), .B1(new_n827), .B2(new_n835), .ZN(G1337gat));
  OAI21_X1  g635(.A(G99gat), .B1(new_n796), .B2(new_n461), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n455), .A2(new_n440), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n808), .B2(new_n838), .ZN(G1338gat));
  AOI21_X1  g638(.A(new_n580), .B1(new_n797), .B2(new_n695), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n425), .A2(G106gat), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n825), .A2(new_n608), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT53), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G106gat), .B1(new_n814), .B2(new_n425), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n845));
  INV_X1    g644(.A(new_n841), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n844), .B(new_n845), .C1(new_n808), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n843), .A2(new_n847), .ZN(G1339gat));
  NAND3_X1  g647(.A1(new_n588), .A2(new_n594), .A3(new_n591), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n596), .A2(KEYINPUT54), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n594), .B1(new_n588), .B2(new_n591), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n601), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n603), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n855), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n540), .A2(new_n541), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n545), .A2(new_n547), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n554), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n558), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n707), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n857), .A2(new_n562), .A3(new_n858), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n605), .A2(new_n607), .A3(new_n863), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n605), .A2(new_n607), .A3(KEYINPUT119), .A4(new_n863), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n663), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n637), .B1(new_n864), .B2(new_n871), .ZN(new_n872));
  NOR4_X1   g671(.A1(new_n707), .A2(new_n733), .A3(new_n608), .A4(new_n562), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(new_n710), .A3(new_n669), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n695), .A2(new_n778), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G113gat), .B1(new_n877), .B2(new_n563), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n695), .A2(new_n457), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n562), .A2(new_n213), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(G1340gat));
  OAI21_X1  g681(.A(G120gat), .B1(new_n877), .B2(new_n765), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT120), .ZN(new_n884));
  INV_X1    g683(.A(new_n880), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n211), .A3(new_n608), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1341gat));
  NOR3_X1   g686(.A1(new_n877), .A2(new_n216), .A3(new_n733), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n637), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n216), .B2(new_n889), .ZN(G1342gat));
  NOR3_X1   g689(.A1(new_n880), .A2(G134gat), .A3(new_n663), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n891), .A2(KEYINPUT121), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT121), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n892), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n877), .B2(new_n663), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(G1343gat));
  OR2_X1    g696(.A1(new_n872), .A2(new_n873), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n754), .A2(new_n710), .A3(new_n669), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n695), .A3(new_n899), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(G141gat), .A3(new_n563), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT124), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT55), .B1(new_n854), .B2(KEYINPUT122), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n903), .B1(KEYINPUT122), .B2(new_n854), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n562), .A3(new_n857), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n866), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n663), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n864), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n873), .B1(new_n908), .B2(new_n733), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n425), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n911), .B(new_n695), .C1(new_n872), .C2(new_n873), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n910), .A2(new_n562), .A3(new_n912), .A4(new_n899), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G141gat), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT58), .B1(new_n902), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n908), .A2(new_n733), .ZN(new_n917));
  INV_X1    g716(.A(new_n873), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n911), .B1(new_n919), .B2(new_n695), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n912), .A2(new_n899), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n910), .A2(KEYINPUT123), .A3(new_n912), .A4(new_n899), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n562), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(KEYINPUT58), .A3(G141gat), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT58), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n901), .B1(KEYINPUT124), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n915), .B1(new_n926), .B2(new_n928), .ZN(G1344gat));
  NOR3_X1   g728(.A1(new_n900), .A2(G148gat), .A3(new_n765), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT125), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT59), .B(new_n223), .C1(new_n924), .C2(new_n608), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT59), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n898), .A2(KEYINPUT57), .A3(new_n695), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n911), .B1(new_n909), .B2(new_n425), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n608), .A3(new_n899), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n933), .B1(new_n937), .B2(G148gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n931), .B1(new_n932), .B2(new_n938), .ZN(G1345gat));
  INV_X1    g738(.A(new_n900), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n245), .A3(new_n637), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n733), .B1(new_n922), .B2(new_n923), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n245), .ZN(G1346gat));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n244), .A3(new_n707), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n663), .B1(new_n922), .B2(new_n923), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n244), .ZN(G1347gat));
  NOR2_X1   g745(.A1(new_n874), .A2(new_n293), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n669), .A3(new_n876), .ZN(new_n948));
  OAI21_X1  g747(.A(G169gat), .B1(new_n948), .B2(new_n563), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n898), .A2(KEYINPUT126), .A3(new_n710), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n951), .B1(new_n874), .B2(new_n293), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n669), .A3(new_n879), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n562), .A2(new_n321), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n949), .B1(new_n954), .B2(new_n955), .ZN(G1348gat));
  NAND2_X1  g755(.A1(new_n947), .A2(new_n876), .ZN(new_n957));
  NOR4_X1   g756(.A1(new_n957), .A2(new_n322), .A3(new_n765), .A4(new_n485), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n954), .A2(new_n765), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n322), .ZN(G1349gat));
  OAI21_X1  g759(.A(G183gat), .B1(new_n948), .B2(new_n733), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n637), .A2(new_n309), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n954), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g763(.A1(new_n947), .A2(new_n669), .A3(new_n876), .A4(new_n707), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n965), .A2(new_n966), .A3(G190gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n965), .B2(G190gat), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n707), .A2(new_n305), .ZN(new_n969));
  OAI22_X1  g768(.A1(new_n967), .A2(new_n968), .B1(new_n954), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT127), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n972));
  OAI221_X1 g771(.A(new_n972), .B1(new_n954), .B2(new_n969), .C1(new_n967), .C2(new_n968), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1351gat));
  NOR2_X1   g773(.A1(new_n754), .A2(new_n485), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n953), .A2(new_n695), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n976), .A2(new_n345), .A3(new_n562), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n710), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n978), .B1(new_n934), .B2(new_n935), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n979), .A2(new_n562), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n345), .B2(new_n980), .ZN(G1352gat));
  NAND3_X1  g780(.A1(new_n976), .A2(new_n346), .A3(new_n608), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT62), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n976), .A2(new_n984), .A3(new_n346), .A4(new_n608), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n936), .A2(new_n608), .ZN(new_n986));
  OAI21_X1  g785(.A(G204gat), .B1(new_n986), .B2(new_n978), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n983), .A2(new_n985), .A3(new_n987), .ZN(G1353gat));
  OAI211_X1 g787(.A(new_n976), .B(new_n637), .C1(new_n360), .C2(new_n359), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n979), .A2(new_n637), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT63), .B1(new_n990), .B2(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  AOI21_X1  g792(.A(G218gat), .B1(new_n976), .B2(new_n707), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n663), .A2(new_n344), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n994), .B1(new_n979), .B2(new_n995), .ZN(G1355gat));
endmodule


