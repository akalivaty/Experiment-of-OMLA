//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935;
  INV_X1    g000(.A(G141gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G148gat), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n203), .A2(new_n205), .B1(KEYINPUT2), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT75), .ZN(new_n208));
  INV_X1    g007(.A(new_n206), .ZN(new_n209));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT75), .A3(new_n206), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n207), .A2(new_n211), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G155gat), .B(G162gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(G141gat), .B(G148gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(G155gat), .B2(G162gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n208), .B(new_n217), .C1(new_n218), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G113gat), .B(G120gat), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n224), .A2(KEYINPUT1), .A3(G134gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n226));
  INV_X1    g025(.A(G120gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G113gat), .ZN(new_n228));
  INV_X1    g027(.A(G113gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G120gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n226), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(G127gat), .B1(new_n225), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n226), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n236));
  INV_X1    g035(.A(G134gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n231), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G127gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n234), .A3(new_n240), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n239), .B1(new_n236), .B2(new_n238), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n222), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT78), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n241), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n242), .A2(new_n243), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(KEYINPUT78), .A3(new_n223), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n246), .A2(G225gat), .A3(G233gat), .A4(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n244), .A2(KEYINPUT4), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n240), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n222), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n252), .A2(KEYINPUT77), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT77), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n253), .A2(new_n257), .A3(new_n254), .A4(new_n222), .ZN(new_n258));
  NAND2_X1  g057(.A1(G225gat), .A2(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT76), .B1(new_n222), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT76), .ZN(new_n262));
  AOI211_X1 g061(.A(new_n262), .B(KEYINPUT3), .C1(new_n216), .C2(new_n221), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n234), .B(new_n240), .C1(new_n222), .C2(new_n260), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n258), .B(new_n259), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n249), .B(new_n251), .C1(new_n256), .C2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT0), .ZN(new_n269));
  XOR2_X1   g068(.A(G57gat), .B(G85gat), .Z(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  OAI221_X1 g070(.A(new_n247), .B1(new_n260), .B2(new_n222), .C1(new_n261), .C2(new_n263), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n252), .A2(new_n255), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n259), .A4(new_n250), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n267), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n271), .B1(new_n267), .B2(new_n274), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI211_X1 g078(.A(new_n276), .B(new_n271), .C1(new_n267), .C2(new_n274), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G8gat), .B(G36gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  XNOR2_X1  g083(.A(G211gat), .B(G218gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G197gat), .B(G204gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT22), .ZN(new_n287));
  INV_X1    g086(.A(G211gat), .ZN(new_n288));
  INV_X1    g087(.A(G218gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n285), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n285), .B1(new_n290), .B2(new_n286), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G226gat), .ZN(new_n295));
  INV_X1    g094(.A(G233gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT26), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G169gat), .ZN(new_n302));
  INV_X1    g101(.A(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT66), .B1(new_n306), .B2(new_n300), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n305), .A2(new_n307), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  INV_X1    g107(.A(G183gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT27), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT27), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G183gat), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  INV_X1    g113(.A(G190gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT66), .A3(new_n304), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n310), .A2(new_n312), .A3(new_n315), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT28), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n308), .A2(new_n316), .A3(new_n317), .A4(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n321), .B1(G183gat), .B2(G190gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT65), .B(KEYINPUT24), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n299), .A2(KEYINPUT23), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n304), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n325), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT23), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n332), .B1(new_n304), .B2(new_n326), .ZN(new_n333));
  NOR2_X1   g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n323), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT64), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT25), .B1(new_n333), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n320), .B1(new_n331), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n320), .B(KEYINPUT73), .C1(new_n331), .C2(new_n341), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n298), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n297), .A2(KEYINPUT29), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n294), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n333), .A2(new_n340), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n333), .A2(KEYINPUT25), .ZN(new_n353));
  OAI22_X1  g152(.A1(new_n352), .A2(KEYINPUT25), .B1(new_n325), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(new_n297), .A3(new_n320), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n355), .A3(new_n293), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n284), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT37), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n284), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n358), .B1(new_n350), .B2(new_n356), .ZN(new_n361));
  OAI211_X1 g160(.A(KEYINPUT85), .B(KEYINPUT38), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n363));
  INV_X1    g162(.A(new_n284), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n345), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n297), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n293), .B1(new_n366), .B2(new_n348), .ZN(new_n367));
  INV_X1    g166(.A(new_n356), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n359), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n361), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT38), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n363), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n350), .A2(new_n356), .A3(new_n284), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n369), .A2(new_n370), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n351), .A2(new_n355), .A3(new_n294), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n377), .A2(KEYINPUT37), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n293), .B1(new_n346), .B2(new_n349), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT38), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n375), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n281), .A2(new_n362), .A3(new_n373), .A4(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n259), .B1(new_n272), .B2(new_n273), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT39), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n246), .A2(new_n248), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n386), .A2(new_n387), .A3(new_n259), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n386), .B2(new_n259), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n383), .A2(new_n384), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n271), .B(new_n385), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT40), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n278), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT30), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n357), .B1(new_n374), .B2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n350), .A2(KEYINPUT30), .A3(new_n356), .A4(new_n284), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT74), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n397), .A2(new_n398), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n394), .B(new_n401), .C1(new_n393), .C2(new_n392), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n261), .B2(new_n263), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n293), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n403), .B1(new_n291), .B2(new_n292), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n222), .B1(new_n406), .B2(new_n260), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G22gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n410), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n405), .A2(new_n413), .A3(new_n408), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT80), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n405), .B2(new_n408), .ZN(new_n417));
  AOI211_X1 g216(.A(new_n410), .B(new_n407), .C1(new_n404), .C2(new_n293), .ZN(new_n418));
  OAI21_X1  g217(.A(G22gat), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT81), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT81), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n421), .B(G22gat), .C1(new_n417), .C2(new_n418), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n411), .A2(new_n423), .A3(new_n412), .A4(new_n414), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n416), .A2(new_n420), .A3(new_n422), .A4(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G78gat), .B(G106gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT31), .B(G50gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430));
  INV_X1    g229(.A(new_n428), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n419), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT82), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n415), .A2(new_n419), .A3(new_n434), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n429), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n430), .B1(new_n429), .B2(new_n436), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n382), .B(new_n402), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(G227gat), .A2(G233gat), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT68), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n342), .A2(new_n442), .A3(new_n247), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n354), .A2(new_n320), .A3(new_n253), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n342), .B2(new_n247), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT69), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n342), .A2(new_n247), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT68), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(new_n444), .A3(new_n443), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT69), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n455), .A2(KEYINPUT32), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G15gat), .B(G43gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT70), .ZN(new_n459));
  XNOR2_X1  g258(.A(G71gat), .B(G99gat), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n459), .B(new_n460), .Z(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n450), .A2(new_n440), .A3(new_n444), .A4(new_n443), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT71), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT34), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT72), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n467), .A2(KEYINPUT72), .A3(new_n469), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT32), .B1(new_n461), .B2(new_n455), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n448), .B2(new_n453), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n463), .A2(new_n472), .A3(new_n473), .A4(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n461), .B1(new_n454), .B2(new_n456), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n470), .B(new_n471), .C1(new_n478), .C2(new_n475), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT36), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT36), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n429), .A2(new_n436), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT83), .ZN(new_n484));
  INV_X1    g283(.A(new_n401), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n280), .B2(new_n279), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n429), .A2(new_n430), .A3(new_n436), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n439), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n477), .A2(new_n479), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n484), .B2(new_n487), .ZN(new_n492));
  INV_X1    g291(.A(new_n486), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(new_n490), .C1(new_n437), .C2(new_n438), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n492), .A2(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n490), .B1(new_n437), .B2(new_n438), .ZN(new_n498));
  NOR4_X1   g297(.A1(new_n498), .A2(new_n494), .A3(KEYINPUT35), .A4(new_n486), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n489), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT16), .ZN(new_n502));
  AOI21_X1  g301(.A(G1gat), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(KEYINPUT91), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n501), .B(KEYINPUT91), .C1(new_n502), .C2(G1gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(G8gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT93), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(G8gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n510), .B(KEYINPUT92), .Z(new_n511));
  AND2_X1   g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT87), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(KEYINPUT87), .A2(KEYINPUT14), .ZN(new_n516));
  OAI22_X1  g315(.A1(new_n515), .A2(new_n516), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  INV_X1    g316(.A(G29gat), .ZN(new_n518));
  INV_X1    g317(.A(G36gat), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n518), .B(new_n519), .C1(new_n513), .C2(new_n514), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G29gat), .A2(G36gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G43gat), .B(G50gat), .Z(new_n524));
  INV_X1    g323(.A(KEYINPUT15), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n521), .B(KEYINPUT89), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(KEYINPUT88), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT88), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n524), .B2(new_n525), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n525), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n522), .B(KEYINPUT90), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n529), .A2(new_n531), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n527), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT17), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n512), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n509), .A2(new_n511), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n535), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(KEYINPUT18), .A3(new_n541), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n538), .B(new_n535), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n541), .B(KEYINPUT13), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G197gat), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT11), .B(G169gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT12), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n544), .A2(new_n556), .A3(new_n545), .A4(new_n548), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(KEYINPUT94), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n549), .A2(new_n559), .A3(new_n554), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n500), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G64gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(G57gat), .ZN(new_n567));
  INV_X1    g366(.A(G57gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(G64gat), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT9), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  OR2_X1    g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n566), .B2(G57gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(new_n568), .B2(G64gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n568), .A2(KEYINPUT95), .A3(G64gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n566), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n575), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n571), .B1(new_n572), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n573), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT21), .ZN(new_n585));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT97), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n591), .B(new_n592), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n538), .B1(KEYINPUT21), .B2(new_n584), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n591), .B(new_n592), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n589), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n595), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n565), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n594), .A2(new_n595), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n599), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n603), .A3(new_n564), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G85gat), .A2(G92gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(KEYINPUT8), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G99gat), .B(G106gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n536), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n535), .A2(new_n615), .B1(KEYINPUT41), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT100), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n622), .B(new_n626), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n605), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT102), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n615), .A2(KEYINPUT10), .A3(new_n584), .ZN(new_n630));
  INV_X1    g429(.A(new_n613), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n584), .B1(new_n631), .B2(KEYINPUT103), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n615), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT10), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT104), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(KEYINPUT104), .A3(new_n634), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n630), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(G230gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(new_n296), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n633), .A2(new_n640), .A3(new_n296), .ZN(new_n643));
  XOR2_X1   g442(.A(G120gat), .B(G148gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT105), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n642), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n643), .B1(new_n639), .B2(new_n641), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n649), .A2(KEYINPUT106), .A3(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n563), .A2(new_n629), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n281), .B(KEYINPUT107), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n401), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT108), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G8gat), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(G8gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(G1325gat));
  AOI21_X1  g468(.A(G15gat), .B1(new_n657), .B2(new_n490), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n482), .B(KEYINPUT109), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(G15gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT110), .Z(new_n673));
  AOI21_X1  g472(.A(new_n670), .B1(new_n657), .B2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n437), .A2(new_n438), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n657), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  INV_X1    g477(.A(KEYINPUT111), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n654), .A2(new_n655), .ZN(new_n680));
  INV_X1    g479(.A(new_n605), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n679), .B1(new_n682), .B2(new_n627), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n656), .A2(new_n605), .ZN(new_n684));
  INV_X1    g483(.A(new_n627), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(KEYINPUT111), .A3(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n500), .A2(new_n562), .A3(new_n683), .A4(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n658), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n687), .A2(G29gat), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT45), .Z(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n439), .A2(new_n482), .A3(new_n488), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n495), .A2(new_n496), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n493), .B(new_n490), .C1(new_n438), .C2(new_n437), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n492), .A2(KEYINPUT86), .A3(new_n496), .A4(new_n493), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n691), .B1(new_n697), .B2(new_n627), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n500), .A2(KEYINPUT44), .A3(new_n685), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT112), .B1(new_n562), .B2(new_n684), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT112), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n682), .A2(new_n702), .A3(new_n561), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n705), .A2(new_n658), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n690), .B1(new_n706), .B2(new_n518), .ZN(G1328gat));
  NOR3_X1   g506(.A1(new_n687), .A2(G36gat), .A3(new_n485), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT46), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n401), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT113), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G36gat), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n710), .A2(KEYINPUT113), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(G1329gat));
  INV_X1    g513(.A(new_n482), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n715), .A3(new_n704), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G43gat), .ZN(new_n717));
  INV_X1    g516(.A(G43gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n490), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n687), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n717), .A2(KEYINPUT47), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n698), .A2(new_n699), .A3(new_n671), .A4(new_n704), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G43gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n721), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT114), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n720), .B1(new_n723), .B2(G43gat), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT114), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT47), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n722), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT115), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT115), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n722), .B(new_n733), .C1(new_n727), .C2(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1330gat));
  NAND4_X1  g534(.A1(new_n698), .A2(new_n699), .A3(new_n675), .A4(new_n704), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G50gat), .ZN(new_n737));
  INV_X1    g536(.A(new_n675), .ZN(new_n738));
  OR3_X1    g537(.A1(new_n687), .A2(G50gat), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(KEYINPUT116), .A3(KEYINPUT48), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT117), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n741), .B2(KEYINPUT48), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n740), .A2(KEYINPUT117), .A3(new_n744), .ZN(new_n748));
  OAI22_X1  g547(.A1(new_n742), .A2(new_n745), .B1(new_n747), .B2(new_n748), .ZN(G1331gat));
  XOR2_X1   g548(.A(new_n628), .B(KEYINPUT102), .Z(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(new_n561), .A3(new_n656), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n751), .A2(KEYINPUT118), .A3(new_n697), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT118), .B1(new_n751), .B2(new_n697), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n688), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(new_n568), .ZN(G1332gat));
  AND2_X1   g555(.A1(new_n752), .A2(new_n753), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n485), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT119), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT119), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n757), .A2(new_n762), .A3(new_n758), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n761), .B1(new_n760), .B2(new_n763), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n757), .A2(new_n767), .A3(new_n490), .ZN(new_n768));
  INV_X1    g567(.A(new_n671), .ZN(new_n769));
  OAI21_X1  g568(.A(G71gat), .B1(new_n754), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1334gat));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n675), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g574(.A1(new_n562), .A2(new_n605), .A3(new_n680), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n700), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(G85gat), .B1(new_n777), .B2(new_n688), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n697), .A2(new_n627), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n562), .A2(new_n605), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT51), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n783), .A3(new_n780), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n656), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n658), .A2(new_n610), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n778), .B1(new_n785), .B2(new_n786), .ZN(G1336gat));
  INV_X1    g586(.A(new_n785), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(new_n611), .A3(new_n401), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT120), .ZN(new_n790));
  OAI21_X1  g589(.A(G92gat), .B1(new_n777), .B2(new_n485), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n792), .A3(KEYINPUT52), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n789), .B(new_n791), .C1(KEYINPUT120), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1337gat));
  XOR2_X1   g595(.A(KEYINPUT121), .B(G99gat), .Z(new_n797));
  NAND3_X1  g596(.A1(new_n788), .A2(new_n490), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n777), .A2(new_n769), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n797), .ZN(G1338gat));
  NAND4_X1  g599(.A1(new_n782), .A2(new_n675), .A3(new_n656), .A4(new_n784), .ZN(new_n801));
  INV_X1    g600(.A(G106gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n700), .A2(G106gat), .A3(new_n675), .A4(new_n776), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT122), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(G1339gat));
  NOR2_X1   g606(.A1(new_n629), .A2(new_n656), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n561), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n540), .A2(new_n541), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n546), .A2(new_n547), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n553), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n557), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n627), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n557), .A2(new_n812), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT123), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n639), .A2(new_n641), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n648), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n642), .A2(KEYINPUT54), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n639), .A2(new_n641), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n649), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n818), .A2(new_n828), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n828), .A2(new_n561), .B1(new_n680), .B2(new_n816), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n627), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n809), .B1(new_n831), .B2(new_n605), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n688), .A2(new_n401), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n832), .A2(new_n738), .A3(new_n490), .A4(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n834), .A2(new_n229), .A3(new_n561), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n832), .A2(new_n485), .A3(new_n492), .A4(new_n658), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n562), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n835), .B1(new_n838), .B2(new_n229), .ZN(G1340gat));
  NOR3_X1   g638(.A1(new_n834), .A2(new_n227), .A3(new_n680), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n656), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n227), .ZN(G1341gat));
  XOR2_X1   g641(.A(KEYINPUT67), .B(G127gat), .Z(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n836), .B2(new_n681), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n681), .A2(new_n843), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n834), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT124), .ZN(G1342gat));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n627), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n826), .A2(new_n649), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n849), .A2(new_n827), .A3(new_n817), .A4(new_n815), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n851), .A2(new_n681), .B1(new_n561), .B2(new_n808), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n688), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n685), .A2(new_n485), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n853), .A2(new_n237), .A3(new_n492), .A4(new_n855), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n834), .B2(new_n627), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(G1343gat));
  NOR2_X1   g659(.A1(new_n671), .A2(new_n738), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n832), .A2(new_n485), .A3(new_n658), .A4(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n202), .B1(new_n862), .B2(new_n561), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT57), .B1(new_n852), .B2(new_n738), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n832), .A2(new_n865), .A3(new_n675), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n688), .A2(new_n715), .A3(new_n401), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n561), .A2(new_n202), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n864), .A2(new_n866), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n870), .B(new_n871), .ZN(G1344gat));
  INV_X1    g671(.A(new_n862), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n204), .A3(new_n656), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n864), .A2(new_n866), .A3(new_n656), .A4(new_n867), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n875), .A2(new_n876), .A3(G148gat), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n875), .B2(G148gat), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(G1345gat));
  NAND3_X1  g678(.A1(new_n873), .A2(new_n212), .A3(new_n605), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n864), .A2(new_n866), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n881), .A2(new_n605), .A3(new_n867), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n880), .B1(new_n882), .B2(new_n212), .ZN(G1346gat));
  NAND4_X1  g682(.A1(new_n853), .A2(new_n213), .A3(new_n855), .A4(new_n861), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n881), .A2(new_n685), .A3(new_n867), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n213), .ZN(G1347gat));
  NOR4_X1   g685(.A1(new_n852), .A2(new_n485), .A3(new_n498), .A4(new_n658), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n302), .A3(new_n562), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(KEYINPUT125), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(KEYINPUT125), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n688), .A2(new_n401), .A3(new_n490), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n852), .A2(new_n675), .A3(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(new_n562), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n889), .A2(new_n890), .B1(new_n302), .B2(new_n893), .ZN(G1348gat));
  NAND3_X1  g693(.A1(new_n887), .A2(new_n303), .A3(new_n656), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n892), .A2(new_n656), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n303), .ZN(G1349gat));
  NAND2_X1  g696(.A1(new_n892), .A2(new_n605), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G183gat), .ZN(new_n899));
  AND2_X1   g698(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n887), .A2(new_n313), .A3(new_n605), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n899), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n887), .A2(new_n315), .A3(new_n685), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n892), .A2(new_n685), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G190gat), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(G1351gat));
  NOR3_X1   g709(.A1(new_n671), .A2(new_n485), .A3(new_n658), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n864), .A2(new_n866), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G197gat), .B1(new_n912), .B2(new_n561), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n852), .A2(new_n658), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n671), .A2(new_n738), .A3(new_n485), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(G197gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n917), .A3(new_n562), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n913), .A2(new_n918), .ZN(G1352gat));
  NOR2_X1   g718(.A1(new_n680), .A2(G204gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n914), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT62), .Z(new_n922));
  OAI21_X1  g721(.A(G204gat), .B1(new_n912), .B2(new_n680), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1353gat));
  NAND3_X1  g723(.A1(new_n916), .A2(new_n288), .A3(new_n605), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n864), .A2(new_n866), .A3(new_n605), .A4(new_n911), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT63), .B1(new_n926), .B2(G211gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(G1354gat));
  NAND2_X1  g728(.A1(new_n912), .A2(KEYINPUT127), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n864), .A2(new_n866), .A3(new_n931), .A4(new_n911), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n930), .A2(new_n685), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G218gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n916), .A2(new_n289), .A3(new_n685), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1355gat));
endmodule


