//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(new_n197), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n195), .A2(KEYINPUT65), .A3(G146), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT65), .B1(new_n195), .B2(G146), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n194), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n198), .B1(new_n201), .B2(new_n189), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n193), .B2(G143), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n195), .A2(KEYINPUT65), .A3(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G128), .A4(new_n194), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n194), .A2(new_n196), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT66), .A2(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n208), .B1(G143), .B2(new_n193), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n209), .A2(new_n210), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n203), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G224), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(G953), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n220), .B(new_n222), .ZN(new_n223));
  XOR2_X1   g037(.A(G110), .B(G122), .Z(new_n224));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n225));
  INV_X1    g039(.A(G119), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G116), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n228));
  INV_X1    g042(.A(G116), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G119), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(KEYINPUT70), .A3(G119), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n226), .A2(KEYINPUT69), .A3(G116), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n227), .A2(new_n230), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT2), .ZN(new_n236));
  INV_X1    g050(.A(G113), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT67), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT2), .A3(G113), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n238), .A2(new_n240), .B1(new_n236), .B2(new_n237), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G104), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT3), .B1(new_n244), .B2(G107), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n246));
  INV_X1    g060(.A(G107), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(G104), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(G107), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n245), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G101), .ZN(new_n251));
  INV_X1    g065(.A(G101), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n245), .A2(new_n248), .A3(new_n252), .A4(new_n249), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(KEYINPUT4), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n250), .A2(new_n255), .A3(G101), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n241), .A2(new_n233), .A3(new_n234), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n243), .A2(new_n254), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n230), .A2(new_n232), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n241), .A2(new_n227), .A3(new_n259), .A4(new_n231), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n247), .A2(G104), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n244), .A2(G107), .ZN(new_n262));
  OAI21_X1  g076(.A(G101), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n253), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n226), .A2(G116), .ZN(new_n265));
  OAI21_X1  g079(.A(G113), .B1(new_n265), .B2(KEYINPUT5), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n233), .A2(new_n267), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n260), .B(new_n264), .C1(new_n266), .C2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT85), .B1(new_n258), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n224), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n258), .A2(new_n271), .A3(new_n269), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n224), .A2(new_n270), .B1(new_n272), .B2(KEYINPUT6), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT85), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n258), .A2(new_n269), .ZN(new_n275));
  AND4_X1   g089(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT6), .A4(new_n224), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n223), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT86), .ZN(new_n278));
  INV_X1    g092(.A(new_n222), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n203), .A2(KEYINPUT7), .A3(new_n279), .A4(new_n219), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n260), .B1(new_n266), .B2(new_n268), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(new_n264), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n229), .A2(KEYINPUT5), .A3(G119), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT87), .B1(new_n284), .B2(new_n237), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT87), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n286), .B(G113), .C1(new_n265), .C2(KEYINPUT5), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n285), .B(new_n287), .C1(new_n233), .C2(new_n267), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n288), .A2(new_n260), .A3(KEYINPUT88), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT88), .B1(new_n288), .B2(new_n260), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n283), .B1(new_n291), .B2(new_n264), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n224), .B(KEYINPUT8), .Z(new_n293));
  AOI21_X1  g107(.A(new_n281), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n203), .A2(new_n219), .B1(KEYINPUT7), .B2(new_n279), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(KEYINPUT89), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n298), .B(new_n223), .C1(new_n273), .C2(new_n276), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n278), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G210), .B1(G237), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n278), .A2(new_n297), .A3(new_n301), .A4(new_n299), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n188), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G953), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G952), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(G234), .B2(G237), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT21), .B(G898), .Z(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(G234), .A2(G237), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(G902), .A3(G953), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n308), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n305), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G113), .B(G122), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(new_n244), .ZN(new_n318));
  INV_X1    g132(.A(G237), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n306), .A3(G214), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n195), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n319), .A2(new_n306), .A3(G143), .A4(G214), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT90), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT18), .B(G131), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n324), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n210), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(G125), .A2(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT80), .B1(new_n329), .B2(new_n330), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n193), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n329), .A2(G146), .A3(new_n330), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT18), .A4(G131), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n327), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT91), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT91), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n327), .A2(new_n337), .A3(new_n341), .A4(new_n338), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT92), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT16), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(new_n329), .B2(new_n330), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n328), .A3(G125), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n193), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n350));
  INV_X1    g164(.A(new_n330), .ZN(new_n351));
  NOR2_X1   g165(.A1(G125), .A2(G140), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT16), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(G146), .A3(new_n347), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n353), .A2(KEYINPUT79), .A3(G146), .A4(new_n347), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT17), .ZN(new_n358));
  INV_X1    g172(.A(G131), .ZN(new_n359));
  AOI211_X1 g173(.A(new_n358), .B(new_n359), .C1(new_n321), .C2(new_n322), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n344), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  AOI211_X1 g176(.A(KEYINPUT92), .B(new_n360), .C1(new_n355), .C2(new_n356), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n323), .B(G131), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(KEYINPUT17), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n318), .B1(new_n343), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G475), .ZN(new_n368));
  INV_X1    g182(.A(G902), .ZN(new_n369));
  INV_X1    g183(.A(new_n354), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n333), .A2(new_n334), .ZN(new_n371));
  MUX2_X1   g185(.A(new_n371), .B(new_n331), .S(KEYINPUT19), .Z(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n372), .B2(new_n193), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n318), .B1(new_n373), .B2(new_n364), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n340), .A2(new_n342), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n367), .A2(new_n368), .A3(new_n369), .A4(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n357), .A2(new_n361), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT92), .ZN(new_n381));
  INV_X1    g195(.A(new_n365), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n357), .A2(new_n344), .A3(new_n361), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n375), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n385), .A2(new_n318), .B1(new_n375), .B2(new_n374), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n386), .A2(KEYINPUT20), .A3(new_n368), .A4(new_n369), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT9), .B(G234), .Z(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(G217), .A3(new_n306), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT95), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n391), .B1(new_n213), .B2(G143), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n195), .A2(KEYINPUT95), .A3(G128), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(G143), .B2(new_n216), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(G134), .ZN(new_n396));
  XNOR2_X1  g210(.A(G116), .B(G122), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT14), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n229), .A2(KEYINPUT14), .A3(G122), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(G107), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT96), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n397), .A2(new_n247), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n399), .A2(KEYINPUT96), .A3(G107), .A4(new_n400), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n396), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G134), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n216), .A2(G143), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT13), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n411), .A2(new_n395), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n395), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n397), .A2(new_n247), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n412), .A2(new_n413), .B1(new_n414), .B2(new_n404), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n390), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n404), .ZN(new_n417));
  INV_X1    g231(.A(new_n413), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n411), .A2(new_n395), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n390), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n420), .B(new_n421), .C1(new_n406), .C2(new_n396), .ZN(new_n422));
  AOI21_X1  g236(.A(G902), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G478), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(KEYINPUT15), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n423), .B(new_n425), .ZN(new_n426));
  OAI22_X1  g240(.A1(new_n343), .A2(new_n366), .B1(KEYINPUT93), .B2(new_n318), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n318), .A2(KEYINPUT93), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n384), .A2(new_n375), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n369), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT94), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n427), .A2(KEYINPUT94), .A3(new_n369), .A4(new_n429), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(G475), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n388), .A2(new_n426), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n316), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n389), .ZN(new_n437));
  OAI21_X1  g251(.A(G221), .B1(new_n437), .B2(G902), .ZN(new_n438));
  XOR2_X1   g252(.A(new_n438), .B(KEYINPUT83), .Z(new_n439));
  INV_X1    g253(.A(G469), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G140), .ZN(new_n441));
  INV_X1    g255(.A(G227), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G953), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n441), .B(new_n443), .Z(new_n444));
  OAI211_X1 g258(.A(G128), .B(new_n194), .C1(new_n199), .C2(new_n200), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n205), .A2(new_n206), .B1(G143), .B2(new_n193), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n217), .A2(new_n213), .ZN(new_n447));
  OAI22_X1  g261(.A1(new_n445), .A2(KEYINPUT1), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n264), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT10), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT11), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n408), .B2(G137), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n408), .A2(G137), .ZN(new_n454));
  INV_X1    g268(.A(G137), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(KEYINPUT11), .A3(G134), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G131), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n453), .A2(new_n456), .A3(new_n359), .A4(new_n454), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n189), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n446), .A2(new_n461), .B1(new_n191), .B2(new_n197), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n254), .A2(new_n462), .A3(new_n256), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n209), .A2(new_n218), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT10), .A3(new_n264), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n451), .A2(new_n460), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n458), .A2(new_n459), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n253), .A2(new_n263), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n468), .A2(new_n209), .A3(new_n218), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G128), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n201), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n468), .B1(new_n472), .B2(new_n209), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n467), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT12), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT12), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n476), .B(new_n467), .C1(new_n469), .C2(new_n473), .ZN(new_n477));
  AND4_X1   g291(.A1(new_n444), .A2(new_n466), .A3(new_n475), .A4(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n460), .A2(KEYINPUT84), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n463), .A2(new_n465), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n473), .A2(KEYINPUT10), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n460), .A2(KEYINPUT84), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n451), .A2(new_n483), .A3(new_n463), .A4(new_n465), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n444), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n440), .B(new_n369), .C1(new_n478), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(G469), .A2(G902), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n466), .A2(new_n475), .A3(new_n477), .ZN(new_n489));
  INV_X1    g303(.A(new_n444), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n482), .A2(new_n484), .A3(new_n444), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(G469), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n439), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  XOR2_X1   g308(.A(KEYINPUT24), .B(G110), .Z(new_n495));
  INV_X1    g309(.A(KEYINPUT75), .ZN(new_n496));
  AND2_X1   g310(.A1(KEYINPUT66), .A2(G128), .ZN(new_n497));
  NOR2_X1   g311(.A1(KEYINPUT66), .A2(G128), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n496), .B(G119), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n226), .B1(new_n214), .B2(new_n215), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT75), .B1(new_n213), .B2(G119), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT76), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT76), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n499), .B(new_n504), .C1(new_n500), .C2(new_n501), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n495), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT23), .B1(new_n213), .B2(G119), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT77), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n226), .B2(G128), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n213), .A2(KEYINPUT77), .A3(G119), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(KEYINPUT23), .B(G119), .C1(new_n497), .C2(new_n498), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(G110), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n354), .B(new_n335), .C1(new_n506), .C2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT78), .B1(new_n513), .B2(G110), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT78), .ZN(new_n517));
  INV_X1    g331(.A(G110), .ZN(new_n518));
  AOI211_X1 g332(.A(new_n517), .B(new_n518), .C1(new_n511), .C2(new_n512), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n503), .A2(new_n495), .A3(new_n505), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n520), .A2(new_n521), .A3(new_n356), .A4(new_n355), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n306), .A2(G221), .A3(G234), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT22), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(G137), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n515), .A2(new_n522), .A3(new_n526), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n369), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT25), .ZN(new_n531));
  INV_X1    g345(.A(G234), .ZN(new_n532));
  OAI21_X1  g346(.A(G217), .B1(new_n532), .B2(G902), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT74), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT25), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n528), .A2(new_n535), .A3(new_n369), .A4(new_n529), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT81), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n531), .A2(KEYINPUT81), .A3(new_n534), .A4(new_n536), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n528), .A2(new_n529), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n534), .A2(G902), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT82), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n539), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n243), .A2(new_n257), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n462), .A2(new_n467), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n455), .A2(G134), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n408), .A2(G137), .ZN(new_n549));
  OAI21_X1  g363(.A(G131), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n459), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n464), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n546), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT28), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n547), .A2(new_n552), .ZN(new_n556));
  INV_X1    g370(.A(new_n546), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n546), .A2(new_n547), .A3(new_n552), .A4(KEYINPUT28), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT26), .B(G101), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n319), .A2(new_n306), .A3(G210), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT72), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n561), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n561), .A3(new_n567), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n560), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n553), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n556), .A2(KEYINPUT30), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT30), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n547), .A2(new_n552), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n574), .B1(new_n578), .B2(new_n557), .ZN(new_n579));
  INV_X1    g393(.A(new_n570), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n568), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT31), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n547), .A2(new_n552), .A3(new_n576), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n576), .B1(new_n547), .B2(new_n552), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n557), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n585), .A2(new_n581), .A3(KEYINPUT31), .A4(new_n553), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n573), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(G472), .A2(G902), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(KEYINPUT32), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT32), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n585), .A2(new_n553), .A3(new_n581), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT31), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n572), .B1(new_n594), .B2(new_n586), .ZN(new_n595));
  INV_X1    g409(.A(new_n589), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT73), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n558), .A2(new_n598), .A3(new_n553), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT73), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(KEYINPUT28), .A3(new_n600), .ZN(new_n601));
  AND4_X1   g415(.A1(KEYINPUT29), .A2(new_n601), .A3(new_n555), .A4(new_n581), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT29), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n560), .B2(new_n571), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n581), .B1(new_n585), .B2(new_n553), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n369), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G472), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n590), .A2(new_n597), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n436), .A2(new_n494), .A3(new_n545), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n494), .A2(new_n539), .A3(new_n540), .A4(new_n544), .ZN(new_n612));
  NAND2_X1  g426(.A1(KEYINPUT97), .A2(G472), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n588), .B2(new_n369), .ZN(new_n614));
  INV_X1    g428(.A(new_n613), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n595), .A2(G902), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n611), .B1(new_n612), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n545), .A2(KEYINPUT98), .A3(new_n494), .A4(new_n617), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n416), .A2(new_n422), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n369), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n424), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT100), .B1(new_n423), .B2(G478), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n390), .B2(KEYINPUT99), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n416), .A2(new_n422), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n628), .B1(new_n416), .B2(new_n422), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n424), .A2(G902), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n625), .A2(new_n626), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n432), .A2(G475), .A3(new_n433), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n379), .A2(new_n387), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n316), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n621), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n316), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n388), .A2(new_n434), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n426), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n621), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT35), .B(G107), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT101), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n645), .B(new_n647), .ZN(G9));
  INV_X1    g462(.A(new_n435), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n523), .A2(KEYINPUT102), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n527), .A2(KEYINPUT36), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n515), .A2(new_n522), .A3(new_n652), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n651), .B1(new_n650), .B2(new_n653), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n543), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n539), .A2(new_n656), .A3(new_n540), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n657), .A2(new_n494), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n642), .A2(new_n649), .A3(new_n658), .A4(new_n617), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT37), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n518), .ZN(G12));
  NAND4_X1  g475(.A1(new_n305), .A2(new_n608), .A3(new_n657), .A4(new_n494), .ZN(new_n662));
  INV_X1    g476(.A(new_n426), .ZN(new_n663));
  INV_X1    g477(.A(new_n308), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(G900), .B2(new_n312), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT103), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n388), .A2(new_n663), .A3(new_n434), .A4(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n213), .ZN(G30));
  XNOR2_X1  g484(.A(new_n666), .B(KEYINPUT39), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n494), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT40), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n303), .A2(new_n304), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT38), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n303), .A2(KEYINPUT38), .A3(new_n304), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n599), .A2(new_n571), .A3(new_n600), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n592), .A2(new_n680), .A3(G472), .ZN(new_n681));
  NAND2_X1  g495(.A1(G472), .A2(G902), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT104), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n597), .A3(new_n590), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n539), .A2(new_n540), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n685), .A2(new_n686), .A3(new_n656), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n635), .A2(new_n636), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n688), .A2(new_n426), .A3(new_n188), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n674), .A2(new_n679), .A3(new_n687), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT105), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  NAND3_X1  g506(.A1(new_n643), .A2(new_n634), .A3(new_n667), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n662), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n193), .ZN(G48));
  INV_X1    g509(.A(new_n608), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n539), .A2(new_n540), .A3(new_n544), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n369), .B1(new_n478), .B2(new_n485), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G469), .ZN(new_n699));
  INV_X1    g513(.A(new_n439), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n700), .A3(new_n486), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n696), .A2(new_n697), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n638), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n642), .A3(new_n644), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  INV_X1    g521(.A(new_n701), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n436), .A2(new_n608), .A3(new_n657), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  NAND2_X1  g524(.A1(new_n594), .A2(new_n586), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n601), .A2(new_n555), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n571), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n596), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n588), .A2(new_n369), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT106), .B(G472), .Z(new_n716));
  AOI21_X1  g530(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n545), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n426), .B1(new_n388), .B2(new_n434), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n188), .B(new_n701), .C1(new_n303), .C2(new_n304), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n718), .A2(new_n315), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  AOI211_X1 g536(.A(new_n633), .B(new_n666), .C1(new_n388), .C2(new_n434), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n657), .A2(new_n717), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n724), .A3(new_n720), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n492), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n491), .A2(new_n492), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n728), .B1(new_n729), .B2(KEYINPUT107), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n439), .B1(new_n731), .B2(new_n488), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n187), .A3(new_n303), .A4(new_n304), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n693), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n545), .A2(new_n608), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n545), .A2(KEYINPUT108), .A3(new_n608), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n734), .A2(KEYINPUT42), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n675), .A2(new_n188), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n545), .A3(new_n608), .A4(new_n732), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n740), .B1(new_n742), .B2(new_n693), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NOR2_X1   g559(.A1(new_n742), .A2(new_n668), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT109), .B(G134), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G36));
  NAND3_X1  g562(.A1(new_n688), .A2(KEYINPUT43), .A3(new_n634), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n634), .A2(new_n388), .A3(new_n434), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n617), .B1(new_n686), .B2(new_n656), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n754), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n741), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT110), .ZN(new_n760));
  INV_X1    g574(.A(new_n486), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n730), .A2(KEYINPUT45), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n729), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(G469), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n487), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n761), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n487), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n700), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n671), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n757), .A2(new_n773), .A3(new_n741), .A4(new_n758), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n760), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  AOI21_X1  g590(.A(new_n439), .B1(new_n768), .B2(new_n769), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT47), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n693), .A2(new_n545), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n696), .A3(new_n741), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  NAND2_X1  g595(.A1(new_n699), .A2(new_n486), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n750), .B1(KEYINPUT49), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(KEYINPUT49), .B2(new_n782), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n439), .A3(new_n679), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n685), .A2(new_n697), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n187), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n187), .B1(new_n677), .B2(new_n678), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n545), .A2(new_n308), .A3(new_n717), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n753), .A2(new_n788), .A3(new_n789), .A4(new_n708), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT50), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n657), .A2(new_n717), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n741), .A2(KEYINPUT115), .A3(new_n708), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n708), .A2(new_n303), .A3(new_n187), .A4(new_n304), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n664), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(KEYINPUT116), .A3(new_n753), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n800));
  INV_X1    g614(.A(new_n753), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n801), .B2(new_n797), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n792), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n688), .A2(new_n798), .A3(new_n633), .A4(new_n786), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n791), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n777), .B(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n808), .B(new_n809), .C1(new_n700), .C2(new_n782), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n782), .A2(new_n700), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT117), .B1(new_n778), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n753), .A2(new_n741), .A3(new_n789), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT113), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n810), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n307), .B1(new_n806), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n814), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n811), .B1(new_n808), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n803), .A2(new_n804), .ZN(new_n822));
  INV_X1    g636(.A(new_n791), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n805), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n737), .A2(new_n738), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n799), .B2(new_n802), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT48), .Z(new_n828));
  AOI21_X1  g642(.A(new_n633), .B1(new_n388), .B2(new_n434), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n798), .A2(new_n829), .A3(new_n786), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n816), .A2(new_n825), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n608), .A2(new_n675), .A3(new_n187), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n663), .A2(new_n388), .A3(new_n434), .A4(new_n667), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n658), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n719), .A2(new_n187), .A3(new_n675), .A4(new_n667), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n685), .A2(new_n686), .A3(new_n656), .A4(new_n732), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n836), .B(new_n725), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n833), .B1(new_n839), .B2(new_n694), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n305), .A2(new_n708), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n693), .A2(new_n841), .A3(new_n792), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n669), .ZN(new_n843));
  INV_X1    g657(.A(new_n694), .ZN(new_n844));
  INV_X1    g658(.A(new_n837), .ZN(new_n845));
  INV_X1    g659(.A(new_n838), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(KEYINPUT52), .A3(new_n844), .A4(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n637), .B1(new_n426), .B2(new_n643), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n619), .A2(new_n850), .A3(new_n642), .A4(new_n620), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n851), .A2(new_n609), .A3(new_n709), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n746), .B1(new_n739), .B2(new_n743), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n702), .A2(new_n850), .A3(new_n642), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n854), .A2(new_n721), .A3(new_n659), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n658), .A2(new_n649), .A3(new_n608), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n724), .A2(new_n829), .A3(new_n732), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n667), .A3(new_n741), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n852), .A2(new_n853), .A3(new_n855), .A4(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n832), .B1(new_n849), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT111), .B1(new_n842), .B2(new_n669), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n833), .B1(new_n845), .B2(new_n846), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n836), .A2(new_n725), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n862), .A2(new_n863), .A3(new_n844), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n840), .ZN(new_n867));
  INV_X1    g681(.A(new_n746), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n744), .A2(new_n859), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n851), .A2(new_n609), .A3(new_n709), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n854), .A2(new_n721), .A3(new_n659), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n867), .A2(new_n869), .A3(KEYINPUT53), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n861), .A2(KEYINPUT112), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n860), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT112), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT53), .A4(new_n867), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT54), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n879));
  OR3_X1    g693(.A1(new_n849), .A2(new_n860), .A3(new_n832), .ZN(new_n880));
  INV_X1    g694(.A(new_n867), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n832), .B1(new_n881), .B2(new_n860), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n753), .A2(new_n720), .A3(new_n789), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n831), .A2(new_n878), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(G952), .A2(G953), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n787), .B1(new_n885), .B2(new_n886), .ZN(G75));
  NAND4_X1  g701(.A1(new_n874), .A2(new_n877), .A3(G210), .A4(G902), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n273), .A2(new_n276), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT118), .ZN(new_n891));
  XOR2_X1   g705(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n892));
  XNOR2_X1  g706(.A(new_n223), .B(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n891), .B(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n888), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n888), .B2(new_n889), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n306), .A2(G952), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G51));
  XOR2_X1   g712(.A(new_n487), .B(KEYINPUT57), .Z(new_n899));
  AND3_X1   g713(.A1(new_n874), .A2(KEYINPUT54), .A3(new_n877), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n878), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n478), .A2(new_n485), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n874), .A2(new_n877), .ZN(new_n904));
  OR3_X1    g718(.A1(new_n904), .A2(new_n369), .A3(new_n765), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n897), .B1(new_n903), .B2(new_n905), .ZN(G54));
  NAND4_X1  g720(.A1(new_n874), .A2(new_n877), .A3(KEYINPUT58), .A4(G902), .ZN(new_n907));
  INV_X1    g721(.A(new_n386), .ZN(new_n908));
  OR3_X1    g722(.A1(new_n907), .A2(new_n368), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n897), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n907), .B2(new_n368), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(G60));
  XOR2_X1   g726(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n913));
  NOR2_X1   g727(.A1(new_n424), .A2(new_n369), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n878), .B2(new_n883), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n631), .B(KEYINPUT120), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n917), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n919), .B(new_n915), .C1(new_n900), .C2(new_n878), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n918), .A2(new_n910), .A3(new_n920), .ZN(G63));
  INV_X1    g735(.A(new_n541), .ZN(new_n922));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT122), .Z(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT60), .Z(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n922), .B1(new_n904), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n654), .A2(new_n655), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n874), .A2(new_n877), .A3(new_n928), .A4(new_n925), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n910), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n927), .A2(KEYINPUT61), .A3(new_n910), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(G66));
  OAI21_X1  g748(.A(G953), .B1(new_n310), .B2(new_n221), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n872), .B2(G953), .ZN(new_n936));
  INV_X1    g750(.A(new_n891), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(G898), .B2(new_n306), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n936), .B(new_n938), .ZN(G69));
  NAND2_X1  g753(.A1(new_n836), .A2(new_n725), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n694), .B1(new_n940), .B2(KEYINPUT111), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n941), .A2(new_n865), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n775), .A2(new_n780), .A3(new_n853), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n689), .A2(new_n675), .ZN(new_n944));
  NOR4_X1   g758(.A1(new_n771), .A2(new_n826), .A3(new_n944), .A4(new_n671), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n306), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n578), .B(KEYINPUT123), .Z(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n372), .ZN(new_n948));
  INV_X1    g762(.A(G900), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(G953), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n941), .A2(new_n690), .A3(new_n865), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n941), .A2(KEYINPUT62), .A3(new_n690), .A4(new_n865), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n735), .A2(new_n188), .A3(new_n675), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n957), .A2(new_n494), .A3(new_n672), .A4(new_n850), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n956), .A2(new_n775), .A3(new_n780), .A4(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n306), .A3(new_n948), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n951), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(G953), .B1(new_n442), .B2(new_n949), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT124), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n961), .B(new_n964), .ZN(G72));
  XNOR2_X1  g779(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(new_n682), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n880), .B2(new_n882), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n579), .B(new_n581), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n897), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n579), .B(KEYINPUT126), .ZN(new_n972));
  INV_X1    g786(.A(new_n872), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n943), .A2(new_n973), .A3(new_n945), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n571), .B(new_n972), .C1(new_n974), .C2(new_n968), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n967), .B1(new_n959), .B2(new_n973), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n972), .A2(new_n571), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n977), .B1(new_n976), .B2(new_n978), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n971), .B(new_n975), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(G57));
endmodule


