//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  AND2_X1   g0010(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT67), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(new_n213), .B2(KEYINPUT67), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n208), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT68), .Z(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n207), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G13), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n208), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT0), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n230), .B(new_n235), .C1(new_n222), .C2(new_n223), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n225), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(G169), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT77), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n256), .A2(KEYINPUT77), .A3(G33), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT69), .B(G1698), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n264), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G87), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n263), .A2(new_n265), .B1(new_n258), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n255), .B1(new_n267), .B2(KEYINPUT83), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(KEYINPUT83), .B2(new_n267), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n254), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n254), .A2(new_n274), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(G232), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n253), .B1(new_n269), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G179), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n269), .A2(new_n277), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT16), .ZN(new_n283));
  INV_X1    g0083(.A(G68), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n257), .A2(new_n259), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n207), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT7), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n284), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G58), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n284), .ZN(new_n292));
  OAI21_X1  g0092(.A(G20), .B1(new_n292), .B2(new_n202), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT78), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(KEYINPUT78), .B(G20), .C1(new_n292), .C2(new_n202), .ZN(new_n296));
  INV_X1    g0096(.A(G159), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n295), .B(new_n296), .C1(new_n297), .C2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n283), .B1(new_n290), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT79), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(KEYINPUT79), .B(new_n283), .C1(new_n290), .C2(new_n300), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n228), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n208), .B2(G33), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n263), .A2(new_n287), .A3(new_n207), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n261), .A2(new_n207), .A3(new_n262), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n284), .B1(new_n309), .B2(KEYINPUT7), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n300), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n307), .B1(new_n311), .B2(KEYINPUT16), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n305), .A2(KEYINPUT80), .A3(new_n312), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n231), .A2(new_n207), .A3(G1), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n206), .A2(G20), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(KEYINPUT81), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT81), .B1(new_n319), .B2(new_n320), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n322), .A2(new_n323), .B1(new_n315), .B2(new_n319), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT82), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n313), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT80), .B1(new_n305), .B2(new_n312), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n282), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT18), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n326), .A2(new_n327), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n331), .A2(KEYINPUT84), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(KEYINPUT84), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n269), .A2(new_n277), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G200), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n269), .B2(new_n277), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n330), .A2(KEYINPUT17), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n305), .A2(new_n312), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT80), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n339), .A2(new_n343), .A3(new_n313), .A4(new_n325), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT17), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT18), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n282), .B(new_n347), .C1(new_n326), .C2(new_n327), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n329), .A2(new_n340), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n307), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n298), .A2(G50), .B1(G20), .B2(new_n284), .ZN(new_n352));
  INV_X1    g0152(.A(G77), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n207), .A2(G33), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT11), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n314), .A2(new_n284), .ZN(new_n358));
  OR3_X1    g0158(.A1(new_n358), .A2(KEYINPUT74), .A3(KEYINPUT12), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT74), .B1(new_n358), .B2(KEYINPUT12), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(KEYINPUT12), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n317), .A2(G68), .A3(new_n320), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n357), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  XOR2_X1   g0164(.A(new_n364), .B(KEYINPUT76), .Z(new_n365));
  INV_X1    g0165(.A(KEYINPUT13), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G232), .A2(G1698), .ZN(new_n367));
  INV_X1    g0167(.A(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT69), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT69), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G1698), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n367), .B1(new_n372), .B2(new_n217), .ZN(new_n373));
  INV_X1    g0173(.A(new_n285), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n373), .A2(new_n374), .B1(G33), .B2(G97), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n375), .A2(new_n255), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n275), .B1(G238), .B2(new_n276), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n366), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(new_n366), .A3(new_n377), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(G179), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(KEYINPUT75), .A2(G169), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n379), .B2(new_n380), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT14), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n382), .ZN(new_n386));
  INV_X1    g0186(.A(new_n380), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n384), .B(new_n386), .C1(new_n387), .C2(new_n378), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n365), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n387), .A2(new_n378), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n364), .B1(new_n391), .B2(G190), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n337), .B2(new_n391), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n320), .A2(G50), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n316), .A2(new_n395), .B1(G50), .B2(new_n315), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT70), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n396), .B(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n203), .A2(G20), .ZN(new_n399));
  INV_X1    g0199(.A(G150), .ZN(new_n400));
  OAI221_X1 g0200(.A(new_n399), .B1(new_n400), .B2(new_n299), .C1(new_n318), .C2(new_n354), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n351), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT9), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT72), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT72), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n398), .A2(new_n406), .A3(KEYINPUT9), .A4(new_n402), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n403), .A2(new_n404), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n275), .B1(G226), .B2(new_n276), .ZN(new_n410));
  INV_X1    g0210(.A(G223), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n374), .B1(new_n411), .B2(new_n368), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n264), .A2(G222), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n254), .B1(G77), .B2(new_n374), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n410), .A2(new_n414), .A3(G190), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(KEYINPUT73), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(KEYINPUT73), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n410), .A2(new_n414), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n416), .A2(new_n417), .B1(G200), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n408), .A2(new_n409), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT10), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT10), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n408), .A2(new_n422), .A3(new_n419), .A4(new_n409), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n418), .A2(G179), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n253), .B2(new_n418), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n426), .A2(new_n403), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G244), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n254), .A2(new_n274), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n374), .A2(new_n264), .A3(G232), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n374), .A2(G238), .A3(G1698), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT71), .B(G107), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n431), .B(new_n432), .C1(new_n374), .C2(new_n433), .ZN(new_n434));
  AOI211_X1 g0234(.A(new_n430), .B(new_n275), .C1(new_n434), .C2(new_n254), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n280), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n319), .A2(new_n298), .B1(G20), .B2(G77), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT15), .B(G87), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n438), .A2(new_n354), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n307), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n320), .A2(G77), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n316), .A2(new_n441), .B1(G77), .B2(new_n315), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n436), .B(new_n444), .C1(G169), .C2(new_n435), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n435), .A2(G190), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(new_n443), .C1(new_n337), .C2(new_n435), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n428), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n350), .A2(new_n394), .A3(new_n424), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n206), .A2(G33), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n307), .A2(new_n315), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G97), .ZN(new_n453));
  INV_X1    g0253(.A(G107), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(KEYINPUT6), .A3(G97), .ZN(new_n455));
  INV_X1    g0255(.A(G97), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(new_n454), .ZN(new_n457));
  NOR2_X1   g0257(.A1(G97), .A2(G107), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n455), .B1(new_n459), .B2(KEYINPUT6), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n460), .A2(G20), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n433), .B1(new_n288), .B2(new_n289), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n298), .A2(G77), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n463), .B(KEYINPUT85), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  OAI221_X1 g0265(.A(new_n453), .B1(G97), .B2(new_n315), .C1(new_n465), .C2(new_n307), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n429), .B1(new_n261), .B2(new_n262), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT4), .B1(new_n467), .B2(new_n264), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT4), .A2(G244), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n264), .A2(new_n470), .B1(G250), .B2(G1698), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n471), .B2(new_n285), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n254), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n273), .A2(G1), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n476), .A2(new_n270), .A3(new_n254), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n255), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G257), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n473), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n331), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n466), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT86), .B1(new_n482), .B2(G200), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n482), .A2(KEYINPUT86), .A3(G200), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n473), .A2(new_n481), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n280), .A3(new_n478), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n482), .A2(new_n253), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n466), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G264), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n478), .B1(new_n493), .B2(new_n479), .ZN(new_n494));
  INV_X1    g0294(.A(G257), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n261), .B2(new_n262), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n496), .A2(G1698), .B1(G33), .B2(G294), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n372), .B1(new_n261), .B2(new_n262), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G250), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n254), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n494), .B1(new_n501), .B2(KEYINPUT99), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n255), .B1(new_n497), .B2(new_n499), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT99), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(new_n331), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n337), .B1(new_n503), .B2(new_n494), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT97), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n509), .B(KEYINPUT25), .C1(new_n315), .C2(G107), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT25), .ZN(new_n511));
  AOI21_X1  g0311(.A(G107), .B1(new_n511), .B2(KEYINPUT97), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n314), .B(new_n512), .C1(KEYINPUT97), .C2(new_n511), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n510), .B(new_n513), .C1(new_n451), .C2(new_n454), .ZN(new_n514));
  XOR2_X1   g0314(.A(new_n514), .B(KEYINPUT98), .Z(new_n515));
  AOI21_X1  g0315(.A(G20), .B1(new_n261), .B2(new_n262), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(KEYINPUT22), .A3(G87), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT23), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(new_n454), .A3(G20), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT95), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n525), .A2(KEYINPUT94), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(KEYINPUT94), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n454), .A2(KEYINPUT71), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G107), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT23), .B1(new_n532), .B2(new_n207), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n257), .A2(new_n259), .A3(new_n207), .A4(G87), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT22), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n524), .A2(new_n528), .A3(new_n533), .A4(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT96), .B1(new_n518), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n524), .A2(new_n533), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n528), .A2(new_n536), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT96), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .A4(new_n517), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n542), .A3(KEYINPUT24), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT24), .ZN(new_n544));
  OAI211_X1 g0344(.A(KEYINPUT96), .B(new_n544), .C1(new_n518), .C2(new_n537), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n351), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n508), .A2(new_n515), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n505), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n477), .B1(G264), .B2(new_n480), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n503), .B2(new_n504), .ZN(new_n550));
  OAI21_X1  g0350(.A(G169), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n503), .A2(new_n494), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G179), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n546), .A2(new_n515), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n547), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n478), .B1(new_n219), .B2(new_n479), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n496), .A2(new_n264), .B1(G303), .B2(new_n285), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n261), .A2(new_n262), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n493), .A2(new_n368), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n560), .A2(KEYINPUT93), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT93), .B1(new_n560), .B2(new_n561), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n558), .B1(new_n564), .B2(new_n254), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n208), .A2(G33), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(new_n228), .B1(G20), .B2(new_n218), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n469), .B(new_n207), .C1(G33), .C2(new_n456), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT20), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(KEYINPUT20), .A3(new_n569), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n315), .A2(G116), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n451), .B2(new_n218), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n253), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n566), .A2(KEYINPUT21), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  INV_X1    g0380(.A(new_n572), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n581), .A2(new_n570), .ZN(new_n582));
  OAI21_X1  g0382(.A(G169), .B1(new_n582), .B2(new_n576), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n580), .B1(new_n583), .B2(new_n565), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n565), .B(G179), .C1(new_n582), .C2(new_n576), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n579), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n565), .A2(new_n335), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n582), .A2(new_n576), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n587), .B(new_n588), .C1(new_n337), .C2(new_n565), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n492), .A2(new_n557), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT92), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n438), .B(KEYINPUT91), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n594), .A2(new_n451), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT90), .ZN(new_n597));
  INV_X1    g0397(.A(new_n438), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(new_n315), .ZN(new_n599));
  AND2_X1   g0399(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n600));
  NOR2_X1   g0400(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n601));
  OAI211_X1 g0401(.A(G33), .B(G97), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n207), .ZN(new_n603));
  NOR2_X1   g0403(.A1(G87), .A2(G97), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT88), .B1(new_n433), .B2(new_n604), .ZN(new_n605));
  AND4_X1   g0405(.A1(KEYINPUT88), .A2(new_n529), .A3(new_n531), .A4(new_n604), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n560), .A2(new_n207), .A3(G68), .ZN(new_n608));
  INV_X1    g0408(.A(new_n600), .ZN(new_n609));
  INV_X1    g0409(.A(new_n601), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n607), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n307), .B1(new_n614), .B2(KEYINPUT89), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n612), .B1(new_n516), .B2(G68), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT89), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n607), .ZN(new_n618));
  AOI211_X1 g0418(.A(new_n597), .B(new_n599), .C1(new_n615), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n608), .A2(new_n613), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT88), .ZN(new_n621));
  INV_X1    g0421(.A(new_n604), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n532), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n433), .A2(KEYINPUT88), .A3(new_n604), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n623), .A2(new_n624), .B1(new_n207), .B2(new_n602), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT89), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n351), .A3(new_n618), .ZN(new_n627));
  INV_X1    g0427(.A(new_n599), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT90), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n596), .B1(new_n619), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n255), .B(G250), .C1(G1), .C2(new_n273), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n271), .A2(new_n475), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n498), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n467), .A2(G1698), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n637), .B2(new_n255), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n253), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n255), .B1(new_n635), .B2(new_n636), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n633), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n280), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n630), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n452), .A2(G87), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n337), .B1(new_n640), .B2(new_n633), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n638), .B2(G190), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n646), .B(new_n648), .C1(new_n619), .C2(new_n629), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n592), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n616), .A2(new_n617), .A3(new_n607), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n617), .B1(new_n616), .B2(new_n607), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n651), .A2(new_n652), .A3(new_n307), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n597), .B1(new_n653), .B2(new_n599), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n627), .A2(KEYINPUT90), .A3(new_n628), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n595), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n592), .B(new_n649), .C1(new_n656), .C2(new_n643), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n591), .B1(new_n650), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n449), .A2(new_n659), .ZN(G372));
  INV_X1    g0460(.A(new_n445), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n393), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n390), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n346), .B(new_n340), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n329), .A2(new_n348), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n424), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT102), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n427), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n491), .ZN(new_n672));
  XNOR2_X1  g0472(.A(KEYINPUT101), .B(KEYINPUT26), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n672), .B(new_n674), .C1(new_n658), .C2(new_n650), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n649), .B1(new_n656), .B2(new_n643), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n491), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n645), .ZN(new_n680));
  INV_X1    g0480(.A(new_n547), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n492), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n586), .A2(new_n556), .A3(KEYINPUT100), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT100), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n551), .A2(new_n553), .B1(new_n546), .B2(new_n515), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n579), .A2(new_n584), .A3(new_n585), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n680), .B1(new_n682), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n679), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n671), .B1(new_n690), .B2(new_n449), .ZN(G369));
  NOR3_X1   g0491(.A1(new_n231), .A2(G1), .A3(G20), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT103), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n588), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n686), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n590), .B2(new_n699), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G330), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n698), .B1(new_n546), .B2(new_n515), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n557), .A2(new_n705), .B1(new_n556), .B2(new_n698), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n686), .A2(new_n698), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n556), .A3(new_n547), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n685), .A2(new_n698), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n712), .ZN(G399));
  NOR2_X1   g0513(.A1(new_n232), .A2(G41), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n227), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n605), .A2(new_n606), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n218), .ZN(new_n717));
  INV_X1    g0517(.A(new_n714), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G1), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n715), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n591), .B(new_n698), .C1(new_n650), .C2(new_n658), .ZN(new_n722));
  INV_X1    g0522(.A(new_n698), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n488), .A2(new_n641), .A3(new_n552), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n565), .A2(G179), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n552), .A2(G179), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(new_n566), .A3(new_n638), .A4(new_n482), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n725), .A2(new_n726), .A3(new_n724), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n723), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT31), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n703), .B1(new_n722), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n723), .B1(new_n679), .B2(new_n689), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n677), .A2(new_n676), .A3(new_n491), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n677), .A2(KEYINPUT92), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n491), .B1(new_n739), .B2(new_n657), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n738), .B1(new_n740), .B2(new_n674), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n685), .A2(new_n686), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n680), .B1(new_n682), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n723), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT29), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n734), .B1(new_n736), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n721), .B1(new_n747), .B2(G1), .ZN(G364));
  NOR2_X1   g0548(.A1(new_n231), .A2(G20), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT104), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n273), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n719), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n704), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G330), .B2(new_n701), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n233), .A2(new_n374), .ZN(new_n755));
  INV_X1    g0555(.A(G355), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n756), .B1(G116), .B2(new_n233), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n263), .A2(new_n233), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n227), .B2(new_n273), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n248), .A2(G45), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n228), .B1(G20), .B2(new_n253), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT105), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT105), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n752), .B1(new_n761), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n207), .A2(G179), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(G190), .A3(G200), .ZN(new_n773));
  INV_X1    g0573(.A(G303), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n772), .A2(new_n331), .A3(new_n337), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n374), .B(new_n775), .C1(G329), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n207), .A2(new_n280), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n337), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G190), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n772), .A2(new_n331), .A3(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n781), .A2(G311), .B1(new_n783), .B2(G283), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n334), .A2(new_n780), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n331), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n207), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n785), .A2(G322), .B1(new_n788), .B2(G294), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n779), .A2(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n334), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(G190), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT33), .B(G317), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n791), .A2(G326), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n778), .A2(new_n784), .A3(new_n789), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n782), .A2(new_n454), .ZN(new_n796));
  XOR2_X1   g0596(.A(KEYINPUT106), .B(G159), .Z(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n776), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n796), .B1(new_n799), .B2(KEYINPUT32), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n787), .A2(new_n456), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G50), .B2(new_n791), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n785), .A2(G58), .B1(new_n792), .B2(G68), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT32), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n798), .A2(new_n804), .B1(new_n781), .B2(G77), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n800), .A2(new_n802), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n773), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n285), .B1(new_n807), .B2(G87), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT107), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n795), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n771), .B1(new_n765), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n768), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n701), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n754), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NAND2_X1  g0615(.A1(new_n723), .A2(new_n444), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n445), .A2(new_n447), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT108), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT108), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n445), .A2(new_n447), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n661), .A2(KEYINPUT109), .A3(new_n723), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT109), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n445), .B2(new_n698), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n735), .B(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n734), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n752), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n765), .A2(new_n766), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n752), .B1(new_n832), .B2(G77), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n374), .B(new_n801), .C1(G311), .C2(new_n777), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n785), .A2(G294), .B1(G107), .B2(new_n807), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n781), .A2(G116), .B1(new_n783), .B2(G87), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n791), .A2(G303), .B1(new_n792), .B2(G283), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n263), .B1(G132), .B2(new_n777), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n787), .A2(new_n291), .B1(new_n782), .B2(new_n284), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G50), .B2(new_n807), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n785), .A2(G143), .B1(new_n792), .B2(G150), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  INV_X1    g0643(.A(new_n791), .ZN(new_n844));
  INV_X1    g0644(.A(new_n781), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n842), .B1(new_n843), .B2(new_n844), .C1(new_n797), .C2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT34), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n839), .B(new_n841), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n838), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n833), .B1(new_n850), .B2(new_n765), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n826), .B2(new_n767), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n830), .A2(new_n852), .ZN(G384));
  OR2_X1    g0653(.A1(new_n460), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n460), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n229), .A4(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT36), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n227), .B(G77), .C1(new_n291), .C2(new_n284), .ZN(new_n858));
  INV_X1    g0658(.A(new_n201), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n284), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(G1), .A3(new_n231), .ZN(new_n861));
  INV_X1    g0661(.A(new_n449), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n736), .A2(new_n862), .A3(new_n746), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n671), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT112), .Z(new_n865));
  NOR2_X1   g0665(.A1(new_n445), .A2(new_n723), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n735), .B2(new_n826), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n311), .A2(KEYINPUT16), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n324), .B1(new_n869), .B2(new_n312), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n870), .A2(new_n696), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n349), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n344), .ZN(new_n873));
  INV_X1    g0673(.A(new_n281), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n278), .B1(new_n874), .B2(G179), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n870), .B1(new_n875), .B2(new_n696), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT37), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n697), .B1(new_n326), .B2(new_n327), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n328), .A2(new_n878), .A3(new_n344), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n872), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n365), .A2(new_n723), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n390), .A2(new_n393), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(new_n390), .B2(new_n393), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n868), .A2(new_n886), .A3(new_n891), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n665), .A2(new_n697), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n663), .A2(new_n698), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT110), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n897));
  XOR2_X1   g0697(.A(KEYINPUT111), .B(KEYINPUT38), .Z(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n878), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n349), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n328), .A2(new_n878), .A3(new_n344), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT37), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n880), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n899), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n897), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n894), .B(new_n896), .C1(new_n906), .C2(KEYINPUT39), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n892), .A2(new_n893), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n865), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n826), .B1(new_n888), .B2(new_n889), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n722), .B2(new_n733), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n901), .A2(new_n904), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n898), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n914), .B2(new_n885), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n872), .B2(new_n881), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n911), .B1(new_n897), .B2(new_n916), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n911), .A2(new_n915), .B1(new_n917), .B2(new_n912), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n449), .B1(new_n722), .B2(new_n733), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n920), .A2(new_n921), .A3(new_n703), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n909), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n750), .A2(G1), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n909), .B2(new_n922), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n857), .B(new_n861), .C1(new_n923), .C2(new_n925), .ZN(G367));
  AND2_X1   g0726(.A1(new_n487), .A2(new_n491), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n466), .A2(new_n723), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n672), .A2(new_n723), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n932), .A2(new_n710), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n927), .A2(new_n685), .A3(new_n928), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n723), .B1(new_n935), .B2(new_n491), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n933), .B2(KEYINPUT42), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n654), .A2(new_n655), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n698), .B1(new_n938), .B2(new_n646), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n680), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n677), .B2(new_n939), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n934), .A2(new_n937), .B1(KEYINPUT43), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n942), .B(new_n943), .Z(new_n944));
  NOR2_X1   g0744(.A1(new_n707), .A2(new_n932), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n714), .B(KEYINPUT41), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n712), .A2(new_n931), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT45), .Z(new_n949));
  NOR2_X1   g0749(.A1(new_n712), .A2(new_n931), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT44), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n707), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT113), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n710), .B1(new_n706), .B2(new_n709), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n704), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n747), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n747), .A2(new_n954), .A3(new_n956), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n953), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n947), .B1(new_n960), .B2(new_n747), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n751), .A2(new_n206), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n946), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n769), .B1(new_n233), .B2(new_n438), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n244), .A2(new_n758), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n752), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n374), .B1(new_n776), .B2(new_n843), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G58), .B2(new_n807), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n785), .A2(G150), .B1(new_n781), .B2(new_n859), .ZN(new_n972));
  INV_X1    g0772(.A(new_n797), .ZN(new_n973));
  AOI22_X1  g0773(.A1(G68), .A2(new_n788), .B1(new_n792), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n782), .A2(new_n353), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n791), .B2(G143), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n971), .A2(new_n972), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n263), .B1(new_n978), .B2(new_n776), .ZN(new_n979));
  INV_X1    g0779(.A(new_n792), .ZN(new_n980));
  INV_X1    g0780(.A(G294), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n980), .A2(new_n981), .B1(new_n456), .B2(new_n782), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n773), .A2(new_n218), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n979), .B(new_n982), .C1(KEYINPUT46), .C2(new_n983), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n785), .A2(G303), .B1(new_n788), .B2(new_n532), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n791), .A2(G311), .B1(new_n781), .B2(G283), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n983), .A2(KEYINPUT46), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT114), .Z(new_n989));
  OAI21_X1  g0789(.A(new_n977), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT47), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n765), .B1(new_n990), .B2(new_n991), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n969), .B1(new_n992), .B2(new_n993), .C1(new_n941), .C2(new_n812), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n964), .A2(new_n994), .ZN(G387));
  INV_X1    g0795(.A(new_n959), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n714), .B1(new_n747), .B2(new_n956), .C1(new_n996), .C2(new_n957), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n706), .A2(new_n812), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n241), .A2(new_n273), .ZN(new_n999));
  INV_X1    g0799(.A(new_n717), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n999), .A2(new_n758), .B1(new_n1000), .B2(new_n755), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n273), .B1(new_n284), .B2(new_n353), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n319), .A2(new_n216), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1002), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1000), .B(new_n1004), .C1(KEYINPUT50), .C2(new_n1003), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1001), .A2(new_n1005), .B1(new_n454), .B2(new_n232), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n752), .B1(new_n1006), .B2(new_n770), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G68), .A2(new_n781), .B1(new_n792), .B2(new_n319), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT115), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n785), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n216), .A2(new_n1010), .B1(new_n844), .B2(new_n297), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n782), .A2(new_n456), .B1(new_n773), .B2(new_n353), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n593), .A2(new_n788), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n263), .B1(G150), .B2(new_n777), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1009), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n791), .A2(G322), .B1(new_n792), .B2(G311), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT116), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(KEYINPUT116), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n785), .A2(G317), .B1(new_n781), .B2(G303), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(G283), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n787), .A2(new_n1025), .B1(new_n773), .B2(new_n981), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(KEYINPUT49), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n560), .B1(G326), .B2(new_n777), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n218), .C2(new_n782), .ZN(new_n1030));
  AOI21_X1  g0830(.A(KEYINPUT49), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1016), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1007), .B1(new_n1032), .B2(new_n765), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n956), .A2(new_n963), .B1(new_n998), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n997), .A2(new_n1034), .ZN(G393));
  INV_X1    g0835(.A(new_n953), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n996), .B2(new_n957), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1037), .A2(new_n960), .A3(new_n714), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT117), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1037), .A2(new_n960), .A3(KEYINPUT117), .A4(new_n714), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n932), .A2(new_n768), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n765), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G311), .A2(new_n785), .B1(new_n791), .B2(G317), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT52), .Z(new_n1046));
  AOI211_X1 g0846(.A(new_n374), .B(new_n796), .C1(G322), .C2(new_n777), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n781), .A2(G294), .B1(new_n807), .B2(G283), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G116), .A2(new_n788), .B1(new_n792), .B2(G303), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G150), .A2(new_n791), .B1(new_n785), .B2(G159), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT51), .Z(new_n1052));
  NOR2_X1   g0852(.A1(new_n773), .A2(new_n284), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n787), .A2(new_n353), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(new_n859), .C2(new_n792), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n845), .A2(new_n318), .B1(new_n266), .B2(new_n782), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n263), .B(new_n1056), .C1(G143), .C2(new_n777), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1052), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1044), .B1(new_n1050), .B2(new_n1058), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n251), .A2(new_n758), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n770), .B1(G97), .B2(new_n232), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n968), .B(new_n1059), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n953), .A2(new_n963), .B1(new_n1043), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1042), .A2(new_n1063), .ZN(G390));
  NAND2_X1  g0864(.A1(new_n862), .A2(new_n734), .ZN(new_n1065));
  AND3_X1   g0865(.A1(new_n863), .A2(new_n671), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n734), .A2(new_n826), .A3(new_n891), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n891), .B1(new_n734), .B2(new_n826), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n868), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1069), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n866), .B1(new_n745), .B2(new_n826), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1071), .A2(new_n1072), .A3(new_n1067), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1066), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n896), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n867), .B2(new_n890), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n894), .B1(new_n906), .B2(KEYINPUT39), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT118), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n896), .B1(new_n914), .B2(new_n885), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n1072), .C2(new_n890), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n672), .B1(new_n658), .B2(new_n650), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n737), .B1(new_n1082), .B2(new_n673), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n677), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1084), .A2(new_n927), .A3(new_n547), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n645), .B1(new_n1085), .B2(new_n742), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n698), .B(new_n826), .C1(new_n1083), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n866), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n890), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1076), .B1(new_n897), .B2(new_n905), .ZN(new_n1090));
  OAI21_X1  g0890(.A(KEYINPUT118), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI221_X4 g0891(.A(new_n1068), .B1(new_n1077), .B2(new_n1078), .C1(new_n1081), .C2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1081), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1067), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1075), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n891), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1079), .B1(new_n1098), .B2(new_n1080), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n1089), .A2(new_n1090), .A3(KEYINPUT118), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1094), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n1068), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n863), .A2(new_n671), .A3(new_n1065), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1093), .A2(new_n1094), .A3(new_n1067), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1096), .A2(new_n1106), .A3(new_n714), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1078), .A2(new_n766), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n791), .A2(G283), .B1(new_n792), .B2(new_n532), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n456), .B2(new_n845), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT120), .Z(new_n1111));
  OAI22_X1  g0911(.A1(new_n787), .A2(new_n353), .B1(new_n782), .B2(new_n284), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n285), .B1(new_n776), .B2(new_n981), .C1(new_n773), .C2(new_n266), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(G116), .C2(new_n785), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n785), .A2(G132), .B1(new_n859), .B2(new_n783), .ZN(new_n1115));
  INV_X1    g0915(.A(G128), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n844), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n843), .A2(new_n980), .B1(new_n845), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n787), .A2(new_n297), .ZN(new_n1120));
  INV_X1    g0920(.A(G125), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n374), .B1(new_n776), .B2(new_n1121), .ZN(new_n1122));
  NOR4_X1   g0922(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .A4(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n773), .A2(new_n400), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1111), .A2(new_n1114), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n752), .B1(new_n319), .B2(new_n832), .C1(new_n1127), .C2(new_n1044), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1108), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n963), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1107), .A2(new_n1131), .A3(KEYINPUT121), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT121), .B1(new_n1107), .B2(new_n1131), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(G378));
  XOR2_X1   g0934(.A(KEYINPUT125), .B(KEYINPUT56), .Z(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n403), .A2(new_n697), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT55), .Z(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n670), .B2(new_n428), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n427), .B(new_n1138), .C1(new_n668), .C2(new_n669), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n669), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT102), .B1(new_n421), .B2(new_n423), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n428), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1138), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n670), .A2(new_n428), .A3(new_n1139), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n1135), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n918), .B2(G330), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n917), .A2(new_n912), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n911), .B(KEYINPUT40), .C1(new_n897), .C2(new_n905), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1151), .A2(new_n1149), .A3(G330), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n908), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1151), .A2(G330), .A3(new_n1152), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1149), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n907), .A2(new_n893), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n892), .A4(new_n1153), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1155), .A2(KEYINPUT57), .A3(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1092), .A2(new_n1095), .A3(new_n1075), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n1103), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n1106), .B2(new_n1066), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1163), .B(new_n714), .C1(KEYINPUT57), .C2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1149), .A2(new_n766), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n752), .B1(new_n832), .B2(new_n859), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n791), .A2(G116), .B1(new_n788), .B2(G68), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT122), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n272), .B1(new_n776), .B2(new_n1025), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n560), .B(new_n1171), .C1(new_n593), .C2(new_n781), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n792), .A2(G97), .B1(new_n807), .B2(G77), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n782), .A2(new_n291), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n785), .B2(G107), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1170), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(KEYINPUT58), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n272), .B1(new_n263), .B2(new_n258), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n216), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1118), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n785), .A2(G128), .B1(new_n807), .B2(new_n1182), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT123), .Z(new_n1184));
  AOI22_X1  g0984(.A1(G150), .A2(new_n788), .B1(new_n792), .B2(G132), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n845), .A2(new_n843), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G125), .B2(new_n791), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT124), .Z(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n973), .A2(new_n783), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G33), .B(G41), .C1(new_n777), .C2(G124), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1181), .B1(KEYINPUT58), .B2(new_n1177), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1168), .B1(new_n1196), .B2(new_n765), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1167), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1164), .B2(new_n962), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1166), .A2(new_n1200), .ZN(G375));
  NAND2_X1  g1001(.A1(new_n1074), .A2(new_n963), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n752), .B1(new_n832), .B2(G68), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n374), .B(new_n975), .C1(G303), .C2(new_n777), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n791), .A2(G294), .B1(G97), .B2(new_n807), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1014), .A3(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n785), .A2(G283), .B1(new_n792), .B2(G116), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n433), .B2(new_n845), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G50), .A2(new_n788), .B1(new_n781), .B2(G150), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n843), .B2(new_n1010), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n263), .B1(G128), .B2(new_n777), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n791), .A2(G132), .B1(G159), .B2(new_n807), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1174), .B1(new_n792), .B2(new_n1182), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1206), .A2(new_n1208), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1203), .B1(new_n1215), .B2(new_n765), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n891), .B2(new_n767), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1202), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n947), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1075), .A2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1066), .A2(new_n1074), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1219), .B1(new_n1221), .B2(new_n1222), .ZN(G381));
  INV_X1    g1023(.A(G387), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(G393), .A2(G396), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(G381), .A2(G384), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1063), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1107), .A2(new_n1131), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1164), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1162), .B2(new_n1103), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT57), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1106), .A2(new_n1066), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n718), .B1(new_n1236), .B2(new_n1161), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1199), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1227), .A2(new_n1229), .A3(new_n1231), .A4(new_n1238), .ZN(G407));
  INV_X1    g1039(.A(G213), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(G343), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1238), .A2(new_n1231), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G407), .A2(G213), .A3(new_n1242), .ZN(G409));
  NAND2_X1  g1043(.A1(new_n1224), .A2(G390), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n814), .B1(new_n997), .B2(new_n1034), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1225), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G387), .A2(new_n1229), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1244), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1246), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  INV_X1    g1052(.A(G384), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1103), .A2(KEYINPUT60), .A3(new_n1070), .A4(new_n1073), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n714), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1222), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1075), .A2(KEYINPUT60), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1253), .B1(new_n1258), .B2(new_n1218), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1222), .B1(KEYINPUT60), .B2(new_n1075), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G384), .B(new_n1219), .C1(new_n1260), .C2(new_n1255), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT126), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1241), .A2(G2897), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .A4(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1263), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1262), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1265), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1199), .B1(new_n1165), .B2(new_n1220), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(new_n1230), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G378), .B2(new_n1238), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1269), .B1(new_n1272), .B2(new_n1241), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT121), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1096), .A2(new_n1106), .A3(new_n714), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1102), .A2(new_n963), .A3(new_n1105), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1108), .B2(new_n1128), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1275), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1107), .A2(new_n1131), .A3(KEYINPUT121), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1166), .A2(new_n1279), .A3(new_n1280), .A4(new_n1200), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1270), .A2(new_n1230), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n1241), .B(new_n1274), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1252), .B(new_n1273), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1241), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1274), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1281), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1286), .B(new_n1287), .C1(new_n1288), .C2(new_n1271), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1251), .B1(new_n1285), .B2(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1273), .A2(new_n1252), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1289), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1283), .A2(KEYINPUT63), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1292), .A2(new_n1294), .A3(new_n1250), .A4(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1291), .A2(new_n1296), .ZN(G405));
  NOR2_X1   g1097(.A1(new_n1238), .A2(new_n1230), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1288), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(KEYINPUT127), .A3(new_n1287), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1287), .A2(KEYINPUT127), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1287), .A2(KEYINPUT127), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1301), .B(new_n1302), .C1(new_n1288), .C2(new_n1298), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1250), .A2(new_n1300), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1250), .B1(new_n1300), .B2(new_n1303), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(G402));
endmodule


