//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT27), .B(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(KEYINPUT28), .A3(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT27), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n209));
  AOI21_X1  g008(.A(G190gat), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n205), .B1(new_n210), .B2(KEYINPUT28), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT26), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n212), .A2(KEYINPUT26), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT25), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n212), .B1(KEYINPUT23), .B2(new_n216), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n204), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n228), .A2(KEYINPUT68), .A3(new_n204), .A4(new_n229), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n225), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT24), .ZN(new_n237));
  NAND3_X1  g036(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT24), .B1(new_n214), .B2(new_n235), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT66), .A3(new_n238), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n223), .B1(new_n234), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n220), .B(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(G183gat), .A2(G190gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(new_n237), .B2(new_n214), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n222), .B1(new_n224), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT25), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n219), .B1(new_n245), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  INV_X1    g052(.A(G127gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(G134gat), .ZN(new_n255));
  INV_X1    g054(.A(G134gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(G127gat), .ZN(new_n257));
  OAI22_X1  g056(.A1(new_n253), .A2(KEYINPUT1), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G120gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G113gat), .ZN(new_n260));
  INV_X1    g059(.A(G113gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G120gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G227gat), .A2(G233gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n267), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n270), .B(new_n219), .C1(new_n245), .C2(new_n251), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT34), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT34), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n268), .A2(new_n274), .A3(new_n269), .A4(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n269), .B1(new_n268), .B2(new_n271), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT32), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G15gat), .B(G43gat), .Z(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT70), .ZN(new_n281));
  XOR2_X1   g080(.A(G71gat), .B(G99gat), .Z(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n283), .A2(KEYINPUT71), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(KEYINPUT71), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(KEYINPUT33), .A3(new_n285), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n276), .A2(KEYINPUT72), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n271), .ZN(new_n288));
  INV_X1    g087(.A(new_n269), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n283), .B1(new_n290), .B2(KEYINPUT32), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT69), .B1(new_n277), .B2(KEYINPUT33), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n273), .A2(new_n297), .A3(new_n275), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n287), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n287), .B2(new_n296), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n202), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n287), .A2(new_n296), .ZN(new_n302));
  INV_X1    g101(.A(new_n298), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n296), .A3(new_n298), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(KEYINPUT90), .A3(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(KEYINPUT76), .A2(G155gat), .A3(G162gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(G141gat), .B(G148gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT76), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT2), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n310), .B(new_n311), .C1(new_n312), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n317));
  INV_X1    g116(.A(G141gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(G148gat), .ZN(new_n319));
  INV_X1    g118(.A(G148gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(G148gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  INV_X1    g123(.A(G155gat), .ZN(new_n325));
  INV_X1    g124(.A(G162gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n324), .B1(new_n327), .B2(KEYINPUT2), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n316), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT4), .B1(new_n330), .B2(new_n267), .ZN(new_n331));
  INV_X1    g130(.A(new_n311), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n332), .A2(new_n308), .A3(new_n309), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n318), .A2(G148gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n320), .A2(G141gat), .ZN(new_n335));
  OAI22_X1  g134(.A1(new_n334), .A2(new_n335), .B1(new_n313), .B2(new_n314), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n333), .A2(new_n336), .B1(new_n323), .B2(new_n328), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n266), .A4(new_n258), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n316), .A2(new_n329), .A3(KEYINPUT78), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT78), .B1(new_n316), .B2(new_n329), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n316), .A2(new_n329), .A3(new_n344), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n267), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n340), .B(new_n341), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT78), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n267), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n270), .A2(new_n337), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n341), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT5), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n350), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n348), .B(new_n349), .C1(new_n357), .C2(new_n356), .ZN(new_n360));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT0), .ZN(new_n362));
  XNOR2_X1  g161(.A(G57gat), .B(G85gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n359), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n364), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n359), .A2(new_n360), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT88), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT88), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n359), .A2(new_n372), .A3(new_n360), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT6), .B1(new_n370), .B2(new_n369), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n368), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT35), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n223), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n206), .A2(new_n207), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT68), .B1(new_n382), .B2(new_n204), .ZN(new_n383));
  INV_X1    g182(.A(new_n233), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n224), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n242), .A2(KEYINPUT66), .A3(new_n238), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT66), .B1(new_n242), .B2(new_n238), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n381), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n247), .A2(new_n250), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT25), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n389), .A2(new_n392), .B1(new_n211), .B2(new_n218), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n380), .B1(new_n393), .B2(KEYINPUT29), .ZN(new_n394));
  NAND2_X1  g193(.A1(G211gat), .A2(G218gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT22), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(G197gat), .A2(G204gat), .ZN(new_n398));
  AND2_X1   g197(.A1(G197gat), .A2(G204gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(G211gat), .B(G218gat), .Z(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G211gat), .B(G218gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(G197gat), .B(G204gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n397), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT74), .ZN(new_n407));
  INV_X1    g206(.A(new_n380), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n252), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n252), .B2(new_n408), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n394), .B(new_n406), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n406), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT29), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n408), .B1(new_n252), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n389), .A2(new_n392), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n380), .B1(new_n415), .B2(new_n219), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n412), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n411), .A2(KEYINPUT75), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT74), .B1(new_n393), .B2(new_n380), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n252), .A2(new_n407), .A3(new_n408), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT75), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n421), .A2(new_n422), .A3(new_n406), .A4(new_n394), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND2_X1  g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT30), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n427), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n418), .A2(new_n431), .A3(new_n423), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n424), .A2(KEYINPUT30), .A3(new_n427), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n379), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G228gat), .A2(G233gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n346), .A2(new_n413), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(new_n412), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT29), .B1(new_n402), .B2(new_n405), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n352), .B(new_n353), .C1(KEYINPUT3), .C2(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n438), .A2(new_n440), .A3(KEYINPUT83), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT83), .B1(new_n438), .B2(new_n440), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n406), .B1(new_n346), .B2(new_n413), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n400), .A2(new_n401), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n403), .B1(new_n397), .B2(new_n404), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n413), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n439), .A2(KEYINPUT82), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n344), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n443), .B1(new_n450), .B2(new_n330), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n436), .B(KEYINPUT81), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  OAI22_X1  g252(.A1(new_n441), .A2(new_n442), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT84), .B1(new_n454), .B2(G22gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(G78gat), .B(G106gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT31), .B(G50gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT85), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(G22gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n438), .A2(new_n440), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n438), .A2(new_n440), .A3(KEYINPUT83), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G22gat), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n446), .A2(new_n447), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n344), .B1(new_n439), .B2(KEYINPUT82), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n330), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n443), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n452), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n466), .A2(new_n467), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n461), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n467), .B1(new_n466), .B2(new_n473), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n477), .B(new_n458), .C1(new_n478), .C2(KEYINPUT84), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n460), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n476), .B1(new_n460), .B2(new_n479), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n307), .A2(new_n435), .A3(KEYINPUT91), .A4(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT91), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT30), .B1(new_n424), .B2(new_n427), .ZN(new_n485));
  AOI211_X1 g284(.A(new_n429), .B(new_n431), .C1(new_n418), .C2(new_n423), .ZN(new_n486));
  INV_X1    g285(.A(new_n432), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n359), .A2(new_n372), .A3(new_n360), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n372), .B1(new_n359), .B2(new_n360), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n364), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n375), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT35), .B1(new_n492), .B2(new_n368), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n482), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n301), .A2(new_n306), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n484), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n365), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT80), .B1(new_n376), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT80), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n375), .A2(new_n499), .A3(new_n365), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n500), .A3(new_n368), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n488), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n460), .A2(new_n479), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n475), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n460), .A2(new_n476), .A3(new_n479), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n504), .B(new_n505), .C1(new_n300), .C2(new_n299), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT35), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n483), .A2(new_n496), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n368), .B(new_n428), .C1(new_n374), .C2(new_n376), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT37), .B1(new_n418), .B2(new_n423), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT38), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n394), .B(new_n412), .C1(new_n409), .C2(new_n410), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n406), .B1(new_n414), .B2(new_n416), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT37), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n511), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n510), .A2(new_n516), .A3(new_n427), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT89), .B1(new_n509), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n510), .ZN(new_n519));
  INV_X1    g318(.A(new_n516), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(new_n431), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n367), .B1(new_n491), .B2(new_n375), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .A4(new_n428), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n519), .A2(new_n431), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n418), .A2(KEYINPUT37), .A3(new_n423), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT38), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n518), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n504), .A2(new_n505), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT3), .ZN(new_n530));
  INV_X1    g329(.A(new_n347), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n530), .A2(new_n531), .B1(new_n331), .B2(new_n339), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n532), .A2(KEYINPUT39), .A3(new_n341), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n533), .A2(new_n364), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n354), .A2(new_n341), .A3(new_n355), .ZN(new_n535));
  OAI211_X1 g334(.A(KEYINPUT39), .B(new_n535), .C1(new_n532), .C2(new_n341), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT87), .B1(new_n537), .B2(KEYINPUT86), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT40), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT86), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT87), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(new_n539), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n538), .A2(new_n539), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n543), .A2(new_n374), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n529), .B1(new_n544), .B2(new_n434), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n547), .A2(KEYINPUT36), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(KEYINPUT36), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n304), .B(new_n305), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  OAI22_X1  g349(.A1(new_n299), .A2(new_n300), .B1(new_n547), .B2(KEYINPUT36), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n502), .A2(new_n529), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n508), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555));
  INV_X1    g354(.A(G29gat), .ZN(new_n556));
  INV_X1    g355(.A(G36gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT14), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT14), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(G29gat), .B2(G36gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n560), .A3(KEYINPUT92), .ZN(new_n564));
  NAND2_X1  g363(.A1(G29gat), .A2(G36gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G43gat), .B(G50gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT15), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n568), .A2(new_n565), .ZN(new_n570));
  INV_X1    g369(.A(new_n567), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT15), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n561), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n566), .A2(new_n569), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n555), .B1(new_n574), .B2(KEYINPUT17), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n566), .A2(new_n569), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n573), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(KEYINPUT93), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G15gat), .B(G22gat), .ZN(new_n582));
  INV_X1    g381(.A(G1gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT16), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n582), .A2(G1gat), .ZN(new_n586));
  OAI21_X1  g385(.A(G8gat), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n582), .A2(new_n584), .ZN(new_n588));
  INV_X1    g387(.A(G8gat), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n588), .B(new_n589), .C1(G1gat), .C2(new_n582), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT94), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT17), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n587), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n591), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n598), .A2(new_n574), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G229gat), .A2(G233gat), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n597), .A2(KEYINPUT18), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n578), .B(new_n591), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n601), .B(KEYINPUT13), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n599), .B1(new_n581), .B2(new_n596), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(new_n609), .B2(new_n601), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n612));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G197gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT11), .B(G169gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n606), .B(new_n611), .C1(new_n612), .C2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n612), .A3(new_n605), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n620), .B(new_n617), .C1(new_n621), .C2(new_n610), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(G64gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(G57gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(G57gat), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(KEYINPUT97), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(KEYINPUT97), .B2(new_n626), .ZN(new_n628));
  NAND2_X1  g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  OR2_X1    g428(.A1(G71gat), .A2(G78gat), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT9), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n626), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT9), .B1(new_n634), .B2(new_n625), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n629), .A3(new_n630), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT21), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n598), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT99), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  XNOR2_X1  g440(.A(G127gat), .B(G155gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n640), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G231gat), .A2(G233gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT98), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G183gat), .B(G211gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n644), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G99gat), .A2(G106gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT8), .ZN(new_n654));
  INV_X1    g453(.A(G85gat), .ZN(new_n655));
  INV_X1    g454(.A(G92gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n654), .A2(KEYINPUT102), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT102), .B1(new_n654), .B2(new_n657), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(KEYINPUT101), .A2(G85gat), .A3(G92gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT7), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT101), .B1(G85gat), .B2(G92gat), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n667));
  XOR2_X1   g466(.A(G99gat), .B(G106gat), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n660), .A2(new_n666), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n660), .A2(new_n669), .A3(new_n666), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n658), .A2(new_n659), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n662), .B(new_n663), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n671), .A2(new_n674), .A3(KEYINPUT103), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n581), .A2(new_n593), .A3(new_n670), .A4(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n670), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n678), .B2(new_n578), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G190gat), .B(G218gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n681), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n676), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G134gat), .B(G162gat), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n685), .B(new_n686), .Z(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n682), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n684), .A2(KEYINPUT104), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n676), .A2(new_n679), .A3(new_n692), .A4(new_n683), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(new_n693), .A3(new_n682), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n687), .B(KEYINPUT100), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n690), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n694), .A2(new_n690), .A3(new_n695), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n652), .B(new_n689), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n675), .A2(new_n637), .A3(new_n670), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT10), .ZN(new_n700));
  INV_X1    g499(.A(new_n637), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n671), .A3(new_n674), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n678), .A2(KEYINPUT10), .A3(new_n701), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(G230gat), .A2(G233gat), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT106), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n703), .B2(new_n704), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n699), .A2(new_n702), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n707), .ZN(new_n714));
  XNOR2_X1  g513(.A(G120gat), .B(G148gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(G176gat), .B(G204gat), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n715), .B(new_n716), .Z(new_n717));
  NAND2_X1  g516(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n717), .ZN(new_n721));
  INV_X1    g520(.A(new_n714), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(new_n709), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n698), .A2(new_n724), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n554), .A2(new_n623), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n501), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g528(.A1(new_n726), .A2(new_n434), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT16), .B(G8gat), .Z(new_n731));
  AND2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n730), .A2(new_n589), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT42), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(KEYINPUT42), .B2(new_n732), .ZN(G1325gat));
  AOI21_X1  g534(.A(G15gat), .B1(new_n726), .B2(new_n307), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n550), .A2(new_n551), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G15gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT107), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n736), .B1(new_n726), .B2(new_n740), .ZN(G1326gat));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n529), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT43), .B(G22gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1327gat));
  OAI21_X1  g543(.A(new_n689), .B1(new_n697), .B2(new_n696), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n554), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n554), .A2(new_n745), .A3(new_n750), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n623), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n724), .A2(new_n652), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G29gat), .B1(new_n755), .B2(new_n501), .ZN(new_n756));
  INV_X1    g555(.A(new_n745), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n508), .B2(new_n553), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n758), .A2(new_n754), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(new_n556), .A3(new_n727), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n756), .A2(new_n761), .ZN(G1328gat));
  NAND3_X1  g561(.A1(new_n759), .A2(new_n557), .A3(new_n434), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT46), .Z(new_n764));
  OAI21_X1  g563(.A(G36gat), .B1(new_n755), .B2(new_n488), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1329gat));
  AND2_X1   g565(.A1(new_n759), .A2(new_n307), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n767), .A2(G43gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n738), .A2(G43gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n755), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n768), .B(new_n772), .C1(new_n755), .C2(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1330gat));
  NAND2_X1  g573(.A1(new_n529), .A2(G50gat), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n759), .A2(new_n529), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n755), .A2(new_n775), .B1(G50gat), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1331gat));
  NAND2_X1  g578(.A1(new_n724), .A2(new_n753), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n698), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n554), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n727), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g584(.A1(new_n434), .A2(KEYINPUT110), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n434), .A2(KEYINPUT110), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  AND2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n789), .B2(new_n790), .ZN(G1333gat));
  OR3_X1    g592(.A1(new_n782), .A2(G71gat), .A3(new_n495), .ZN(new_n794));
  OAI21_X1  g593(.A(G71gat), .B1(new_n782), .B2(new_n737), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g596(.A1(new_n783), .A2(new_n529), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g598(.A1(new_n780), .A2(new_n652), .ZN(new_n800));
  INV_X1    g599(.A(new_n748), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n751), .B(new_n800), .C1(new_n758), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT111), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n749), .A2(new_n804), .A3(new_n751), .A4(new_n800), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n803), .A2(new_n727), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n554), .A2(new_n808), .A3(new_n745), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n652), .A2(new_n623), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n758), .A2(new_n808), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n807), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n746), .A2(KEYINPUT112), .ZN(new_n814));
  INV_X1    g613(.A(new_n810), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n758), .B2(new_n808), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n816), .A3(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n727), .A2(new_n655), .A3(new_n724), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n806), .A2(new_n655), .B1(new_n819), .B2(new_n820), .ZN(G1336gat));
  INV_X1    g620(.A(new_n724), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n788), .A2(G92gat), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825));
  OAI21_X1  g624(.A(G92gat), .B1(new_n802), .B2(new_n788), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n814), .A2(new_n816), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT51), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI211_X1 g629(.A(KEYINPUT113), .B(new_n807), .C1(new_n814), .C2(new_n816), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n803), .A2(new_n434), .A3(new_n805), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n832), .A2(new_n823), .B1(G92gat), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n827), .B1(new_n834), .B2(new_n825), .ZN(G1337gat));
  AND3_X1   g634(.A1(new_n803), .A2(new_n738), .A3(new_n805), .ZN(new_n836));
  INV_X1    g635(.A(G99gat), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n307), .A2(new_n837), .A3(new_n724), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n836), .A2(new_n837), .B1(new_n819), .B2(new_n838), .ZN(G1338gat));
  NAND3_X1  g638(.A1(new_n803), .A2(new_n529), .A3(new_n805), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G106gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n829), .B1(new_n811), .B2(new_n812), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n807), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n829), .A3(KEYINPUT51), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n822), .A2(new_n482), .A3(G106gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849));
  OAI21_X1  g648(.A(G106gat), .B1(new_n802), .B2(new_n482), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n845), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n853), .B1(new_n813), .B2(new_n817), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n849), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n811), .A2(new_n807), .A3(new_n812), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT51), .B1(new_n814), .B2(new_n816), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n845), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n858), .A2(KEYINPUT114), .A3(new_n851), .A4(new_n850), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n848), .A2(new_n860), .ZN(G1339gat));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n709), .A2(new_n710), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT106), .B(new_n707), .C1(new_n703), .C2(new_n704), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n703), .A2(new_n707), .A3(new_n704), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT54), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n717), .B1(new_n709), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT55), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n862), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n865), .A2(KEYINPUT54), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n708), .A2(new_n872), .A3(new_n711), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n873), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n869), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n719), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n606), .A2(new_n618), .A3(new_n611), .ZN(new_n876));
  OAI22_X1  g675(.A1(new_n609), .A2(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n616), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT55), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n873), .A2(new_n869), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n745), .A2(new_n875), .A3(new_n882), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n881), .A2(new_n880), .B1(new_n619), .B2(new_n622), .ZN(new_n884));
  INV_X1    g683(.A(new_n879), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n875), .A2(new_n884), .B1(new_n724), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n883), .B1(new_n886), .B2(new_n745), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n651), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n698), .A2(new_n623), .A3(new_n724), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n482), .ZN(new_n892));
  INV_X1    g691(.A(new_n788), .ZN(new_n893));
  NOR4_X1   g692(.A1(new_n892), .A2(new_n501), .A3(new_n495), .A4(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(new_n261), .A3(new_n753), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n891), .A2(new_n727), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n506), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n623), .A3(new_n788), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n896), .B1(new_n899), .B2(new_n261), .ZN(G1340gat));
  OAI21_X1  g699(.A(G120gat), .B1(new_n895), .B2(new_n822), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n788), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n724), .A2(new_n259), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT116), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n901), .B1(new_n902), .B2(new_n904), .ZN(G1341gat));
  NOR3_X1   g704(.A1(new_n895), .A2(new_n254), .A3(new_n651), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n902), .A2(KEYINPUT117), .A3(new_n651), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(G127gat), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT117), .B1(new_n902), .B2(new_n651), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(G1342gat));
  OAI21_X1  g709(.A(G134gat), .B1(new_n895), .B2(new_n757), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n757), .A2(new_n434), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n898), .A2(new_n256), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n911), .A2(new_n915), .A3(new_n916), .ZN(G1343gat));
  NAND3_X1  g716(.A1(new_n788), .A2(new_n727), .A3(new_n737), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n891), .A2(KEYINPUT57), .A3(new_n529), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n889), .B1(new_n887), .B2(new_n651), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n482), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n918), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n318), .B1(new_n923), .B2(new_n623), .ZN(new_n924));
  NAND2_X1  g723(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n925));
  NOR4_X1   g724(.A1(new_n921), .A2(new_n501), .A3(new_n482), .A4(new_n738), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n788), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n753), .A2(G141gat), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n925), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT120), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n931), .B(new_n933), .Z(G1344gat));
  NOR2_X1   g733(.A1(new_n320), .A2(KEYINPUT59), .ZN(new_n935));
  INV_X1    g734(.A(new_n923), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n822), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n871), .A2(new_n874), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n884), .A2(new_n938), .A3(new_n720), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n724), .A2(new_n885), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n745), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n883), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT122), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n944), .B(new_n883), .C1(new_n886), .C2(new_n745), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(new_n651), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n482), .B1(new_n946), .B2(new_n890), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n919), .B1(new_n947), .B2(KEYINPUT57), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n918), .A2(new_n822), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G148gat), .ZN(new_n951));
  XNOR2_X1  g750(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT123), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n320), .B1(new_n948), .B2(new_n949), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n955), .A2(new_n956), .A3(new_n952), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n937), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n926), .A2(new_n320), .A3(new_n724), .A4(new_n788), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1345gat));
  OAI21_X1  g759(.A(G155gat), .B1(new_n936), .B2(new_n651), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n652), .A2(new_n325), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n927), .B2(new_n962), .ZN(G1346gat));
  OAI21_X1  g762(.A(G162gat), .B1(new_n936), .B2(new_n757), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n926), .A2(new_n326), .A3(new_n912), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1347gat));
  NOR4_X1   g765(.A1(new_n921), .A2(new_n727), .A3(new_n506), .A4(new_n788), .ZN(new_n967));
  AOI21_X1  g766(.A(G169gat), .B1(new_n967), .B2(new_n623), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n727), .A2(new_n488), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(new_n307), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n892), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n623), .A2(G169gat), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1348gat));
  INV_X1    g772(.A(G176gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n967), .A2(new_n974), .A3(new_n724), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n892), .A2(new_n822), .A3(new_n970), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n974), .ZN(G1349gat));
  NAND3_X1  g776(.A1(new_n967), .A2(new_n203), .A3(new_n652), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n892), .A2(new_n651), .A3(new_n970), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n979), .B2(new_n382), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g780(.A1(new_n967), .A2(new_n204), .A3(new_n745), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n971), .A2(new_n745), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n984), .B2(G190gat), .ZN(new_n985));
  AOI211_X1 g784(.A(KEYINPUT61), .B(new_n204), .C1(new_n971), .C2(new_n745), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n987), .B(new_n988), .ZN(G1351gat));
  NOR2_X1   g788(.A1(new_n921), .A2(new_n727), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n893), .A2(new_n529), .A3(new_n737), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g793(.A(G197gat), .B1(new_n994), .B2(new_n623), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n969), .A2(new_n737), .ZN(new_n996));
  XNOR2_X1  g795(.A(new_n996), .B(KEYINPUT125), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n948), .A2(new_n997), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n623), .A2(G197gat), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(G1352gat));
  XOR2_X1   g799(.A(KEYINPUT126), .B(G204gat), .Z(new_n1001));
  NAND3_X1  g800(.A1(new_n994), .A2(new_n724), .A3(new_n1001), .ZN(new_n1002));
  XOR2_X1   g801(.A(new_n1002), .B(KEYINPUT62), .Z(new_n1003));
  AND2_X1   g802(.A1(new_n998), .A2(new_n724), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1003), .B1(new_n1001), .B2(new_n1004), .ZN(G1353gat));
  INV_X1    g804(.A(G211gat), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n996), .A2(new_n651), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1006), .B1(new_n948), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(KEYINPUT63), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n1006), .A3(new_n652), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(G1354gat));
  INV_X1    g810(.A(G218gat), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1012), .B1(new_n993), .B2(new_n757), .ZN(new_n1013));
  XOR2_X1   g812(.A(new_n1013), .B(KEYINPUT127), .Z(new_n1014));
  NOR2_X1   g813(.A1(new_n757), .A2(new_n1012), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n1014), .B1(new_n998), .B2(new_n1015), .ZN(G1355gat));
endmodule


