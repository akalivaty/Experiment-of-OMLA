

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  NOR2_X1 U323 ( .A1(n408), .A2(n521), .ZN(n409) );
  XNOR2_X1 U324 ( .A(n529), .B(n530), .ZN(n408) );
  XNOR2_X1 U325 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U326 ( .A(KEYINPUT99), .B(n478), .Z(n571) );
  XOR2_X1 U327 ( .A(n294), .B(KEYINPUT86), .Z(n291) );
  AND2_X1 U328 ( .A1(n506), .A2(n575), .ZN(n361) );
  INV_X1 U329 ( .A(KEYINPUT104), .ZN(n469) );
  XNOR2_X1 U330 ( .A(n327), .B(n326), .ZN(n329) );
  XNOR2_X1 U331 ( .A(n329), .B(n328), .ZN(n331) );
  AND2_X1 U332 ( .A1(n572), .A2(n451), .ZN(n452) );
  XNOR2_X1 U333 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U334 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U335 ( .A(n351), .B(n350), .ZN(n352) );
  NOR2_X1 U336 ( .A1(n582), .A2(n492), .ZN(n493) );
  XNOR2_X1 U337 ( .A(n339), .B(n338), .ZN(n388) );
  NOR2_X1 U338 ( .A1(n532), .A2(n453), .ZN(n454) );
  XOR2_X1 U339 ( .A(KEYINPUT123), .B(n454), .Z(n568) );
  XNOR2_X1 U340 ( .A(n360), .B(n359), .ZN(n553) );
  XNOR2_X1 U341 ( .A(n407), .B(n406), .ZN(n521) );
  XNOR2_X1 U342 ( .A(n495), .B(KEYINPUT38), .ZN(n504) );
  XNOR2_X1 U343 ( .A(n455), .B(G190GAT), .ZN(n456) );
  XNOR2_X1 U344 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n293) );
  XNOR2_X1 U346 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n292) );
  XNOR2_X1 U347 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(G176GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n291), .B(n295), .ZN(n393) );
  XOR2_X1 U350 ( .A(G113GAT), .B(KEYINPUT0), .Z(n436) );
  XOR2_X1 U351 ( .A(n436), .B(G127GAT), .Z(n297) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U354 ( .A(G43GAT), .B(G134GAT), .Z(n374) );
  XOR2_X1 U355 ( .A(n298), .B(n374), .Z(n306) );
  XOR2_X1 U356 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n300) );
  XNOR2_X1 U357 ( .A(G99GAT), .B(G120GAT), .ZN(n299) );
  XNOR2_X1 U358 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U359 ( .A(G183GAT), .B(KEYINPUT85), .Z(n302) );
  XNOR2_X1 U360 ( .A(G15GAT), .B(G71GAT), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n393), .B(n307), .ZN(n532) );
  XNOR2_X1 U365 ( .A(G15GAT), .B(G64GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(G22GAT), .B(G78GAT), .ZN(n413) );
  INV_X1 U367 ( .A(n413), .ZN(n308) );
  XOR2_X1 U368 ( .A(n309), .B(n308), .Z(n323) );
  XNOR2_X1 U369 ( .A(G1GAT), .B(G127GAT), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n310), .B(G155GAT), .ZN(n430) );
  XOR2_X1 U371 ( .A(KEYINPUT83), .B(n430), .Z(n312) );
  NAND2_X1 U372 ( .A1(G231GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U374 ( .A(KEYINPUT82), .B(KEYINPUT15), .Z(n314) );
  XNOR2_X1 U375 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n313) );
  XNOR2_X1 U376 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U377 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U378 ( .A(KEYINPUT81), .B(G211GAT), .Z(n318) );
  XNOR2_X1 U379 ( .A(G8GAT), .B(G183GAT), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n404) );
  XNOR2_X1 U381 ( .A(G71GAT), .B(G57GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n319), .B(KEYINPUT13), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n404), .B(n333), .ZN(n320) );
  XNOR2_X1 U384 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U385 ( .A(n323), .B(n322), .Z(n582) );
  XOR2_X1 U386 ( .A(n582), .B(KEYINPUT113), .Z(n569) );
  XOR2_X1 U387 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n325) );
  NAND2_X1 U388 ( .A1(G230GAT), .A2(G233GAT), .ZN(n324) );
  XOR2_X1 U389 ( .A(n325), .B(n324), .Z(n327) );
  XNOR2_X1 U390 ( .A(G176GAT), .B(G78GAT), .ZN(n326) );
  XOR2_X1 U391 ( .A(G99GAT), .B(G85GAT), .Z(n377) );
  XOR2_X1 U392 ( .A(G92GAT), .B(G64GAT), .Z(n402) );
  XOR2_X1 U393 ( .A(n377), .B(n402), .Z(n328) );
  XOR2_X1 U394 ( .A(G120GAT), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U395 ( .A(n431), .B(KEYINPUT32), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n339) );
  XNOR2_X1 U397 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n332), .B(G204GAT), .ZN(n421) );
  XOR2_X1 U399 ( .A(n421), .B(n333), .Z(n337) );
  XOR2_X1 U400 ( .A(KEYINPUT72), .B(KEYINPUT75), .Z(n335) );
  XNOR2_X1 U401 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n334) );
  XNOR2_X1 U402 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U403 ( .A(n388), .B(KEYINPUT64), .ZN(n341) );
  INV_X1 U404 ( .A(KEYINPUT41), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n506) );
  XOR2_X1 U406 ( .A(G15GAT), .B(G113GAT), .Z(n343) );
  XNOR2_X1 U407 ( .A(G169GAT), .B(G43GAT), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n345) );
  XOR2_X1 U409 ( .A(G36GAT), .B(G50GAT), .Z(n344) );
  XNOR2_X1 U410 ( .A(n345), .B(n344), .ZN(n351) );
  XOR2_X1 U411 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n347) );
  XNOR2_X1 U412 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n346) );
  XNOR2_X1 U413 ( .A(n347), .B(n346), .ZN(n349) );
  NAND2_X1 U414 ( .A1(G229GAT), .A2(G233GAT), .ZN(n348) );
  XOR2_X1 U415 ( .A(n352), .B(KEYINPUT69), .Z(n360) );
  XOR2_X1 U416 ( .A(G29GAT), .B(KEYINPUT7), .Z(n354) );
  XNOR2_X1 U417 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n379) );
  XNOR2_X1 U419 ( .A(n379), .B(KEYINPUT68), .ZN(n358) );
  XOR2_X1 U420 ( .A(G1GAT), .B(G197GAT), .Z(n356) );
  XNOR2_X1 U421 ( .A(G141GAT), .B(G22GAT), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n357) );
  INV_X1 U423 ( .A(n553), .ZN(n575) );
  XNOR2_X1 U424 ( .A(n361), .B(KEYINPUT46), .ZN(n362) );
  NOR2_X1 U425 ( .A1(n569), .A2(n362), .ZN(n363) );
  XNOR2_X1 U426 ( .A(KEYINPUT114), .B(n363), .ZN(n384) );
  XOR2_X1 U427 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n365) );
  XNOR2_X1 U428 ( .A(G190GAT), .B(KEYINPUT65), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n370) );
  XNOR2_X1 U430 ( .A(G50GAT), .B(KEYINPUT77), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n366), .B(G162GAT), .ZN(n425) );
  XOR2_X1 U432 ( .A(n425), .B(KEYINPUT79), .Z(n368) );
  NAND2_X1 U433 ( .A1(G232GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n383) );
  XOR2_X1 U436 ( .A(KEYINPUT78), .B(KEYINPUT10), .Z(n372) );
  XNOR2_X1 U437 ( .A(G92GAT), .B(KEYINPUT67), .ZN(n371) );
  XNOR2_X1 U438 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U439 ( .A(n373), .B(G218GAT), .Z(n376) );
  XNOR2_X1 U440 ( .A(n374), .B(G106GAT), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n378) );
  XOR2_X1 U442 ( .A(n378), .B(n377), .Z(n381) );
  XOR2_X1 U443 ( .A(G36GAT), .B(KEYINPUT80), .Z(n405) );
  XNOR2_X1 U444 ( .A(n379), .B(n405), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U446 ( .A(n383), .B(n382), .Z(n565) );
  AND2_X1 U447 ( .A1(n384), .A2(n565), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n385), .B(KEYINPUT47), .ZN(n392) );
  XOR2_X1 U449 ( .A(KEYINPUT45), .B(KEYINPUT66), .Z(n387) );
  XOR2_X1 U450 ( .A(KEYINPUT36), .B(n565), .Z(n584) );
  NAND2_X1 U451 ( .A1(n582), .A2(n584), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n390) );
  NOR2_X1 U453 ( .A1(n575), .A2(n388), .ZN(n389) );
  NAND2_X1 U454 ( .A1(n390), .A2(n389), .ZN(n391) );
  NAND2_X1 U455 ( .A1(n392), .A2(n391), .ZN(n529) );
  XNOR2_X1 U456 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n530) );
  XNOR2_X1 U457 ( .A(n393), .B(G204GAT), .ZN(n401) );
  XOR2_X1 U458 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n395) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U460 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U461 ( .A(KEYINPUT91), .B(G218GAT), .Z(n397) );
  XNOR2_X1 U462 ( .A(KEYINPUT92), .B(KEYINPUT21), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U464 ( .A(G197GAT), .B(n398), .Z(n418) );
  XOR2_X1 U465 ( .A(n399), .B(n418), .Z(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U467 ( .A(n403), .B(n402), .Z(n407) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U469 ( .A(n409), .B(KEYINPUT54), .ZN(n572) );
  XOR2_X1 U470 ( .A(G148GAT), .B(KEYINPUT93), .Z(n411) );
  XNOR2_X1 U471 ( .A(G155GAT), .B(KEYINPUT22), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n415) );
  NAND2_X1 U474 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n429) );
  XOR2_X1 U476 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n417) );
  XNOR2_X1 U477 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U479 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U480 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n420), .B(KEYINPUT3), .ZN(n432) );
  XNOR2_X1 U482 ( .A(n432), .B(n421), .ZN(n422) );
  XNOR2_X1 U483 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U484 ( .A(n424), .B(G211GAT), .Z(n427) );
  XNOR2_X1 U485 ( .A(n425), .B(KEYINPUT94), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U487 ( .A(n429), .B(n428), .Z(n472) );
  XOR2_X1 U488 ( .A(n431), .B(n430), .Z(n438) );
  XOR2_X1 U489 ( .A(KEYINPUT96), .B(n432), .Z(n434) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U494 ( .A(G85GAT), .B(G162GAT), .Z(n440) );
  XNOR2_X1 U495 ( .A(G29GAT), .B(G134GAT), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U497 ( .A(n442), .B(n441), .Z(n450) );
  XOR2_X1 U498 ( .A(KEYINPUT97), .B(G57GAT), .Z(n444) );
  XNOR2_X1 U499 ( .A(KEYINPUT95), .B(KEYINPUT98), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U501 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n446) );
  XNOR2_X1 U502 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U505 ( .A(n450), .B(n449), .Z(n478) );
  INV_X1 U506 ( .A(n571), .ZN(n464) );
  NOR2_X1 U507 ( .A1(n472), .A2(n464), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n452), .B(KEYINPUT55), .ZN(n453) );
  INV_X1 U509 ( .A(n565), .ZN(n545) );
  NAND2_X1 U510 ( .A1(n568), .A2(n545), .ZN(n457) );
  XOR2_X1 U511 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n455) );
  NAND2_X1 U512 ( .A1(n568), .A2(n506), .ZN(n461) );
  XOR2_X1 U513 ( .A(G176GAT), .B(KEYINPUT56), .Z(n459) );
  XNOR2_X1 U514 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  NOR2_X1 U517 ( .A1(n388), .A2(n553), .ZN(n494) );
  XOR2_X1 U518 ( .A(KEYINPUT16), .B(KEYINPUT84), .Z(n463) );
  NAND2_X1 U519 ( .A1(n582), .A2(n565), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n463), .B(n462), .ZN(n482) );
  XNOR2_X1 U521 ( .A(n532), .B(KEYINPUT88), .ZN(n466) );
  XOR2_X1 U522 ( .A(n521), .B(KEYINPUT27), .Z(n475) );
  NAND2_X1 U523 ( .A1(n464), .A2(n475), .ZN(n550) );
  XOR2_X1 U524 ( .A(n472), .B(KEYINPUT28), .Z(n525) );
  INV_X1 U525 ( .A(n525), .ZN(n465) );
  NOR2_X1 U526 ( .A1(n550), .A2(n465), .ZN(n534) );
  NAND2_X1 U527 ( .A1(n466), .A2(n534), .ZN(n481) );
  NOR2_X1 U528 ( .A1(n521), .A2(n532), .ZN(n467) );
  XOR2_X1 U529 ( .A(KEYINPUT103), .B(n467), .Z(n468) );
  NOR2_X1 U530 ( .A1(n472), .A2(n468), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U532 ( .A(KEYINPUT25), .B(n471), .Z(n477) );
  NAND2_X1 U533 ( .A1(n532), .A2(n472), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n473), .B(KEYINPUT102), .ZN(n474) );
  XOR2_X1 U535 ( .A(KEYINPUT26), .B(n474), .Z(n549) );
  NAND2_X1 U536 ( .A1(n549), .A2(n475), .ZN(n476) );
  NAND2_X1 U537 ( .A1(n477), .A2(n476), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n479), .A2(n478), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n481), .A2(n480), .ZN(n491) );
  AND2_X1 U540 ( .A1(n482), .A2(n491), .ZN(n507) );
  NAND2_X1 U541 ( .A1(n494), .A2(n507), .ZN(n489) );
  NOR2_X1 U542 ( .A1(n571), .A2(n489), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT34), .B(KEYINPUT105), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NOR2_X1 U546 ( .A1(n521), .A2(n489), .ZN(n486) );
  XOR2_X1 U547 ( .A(G8GAT), .B(n486), .Z(G1325GAT) );
  NOR2_X1 U548 ( .A1(n532), .A2(n489), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n525), .A2(n489), .ZN(n490) );
  XOR2_X1 U552 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  NAND2_X1 U553 ( .A1(n584), .A2(n491), .ZN(n492) );
  XOR2_X1 U554 ( .A(KEYINPUT37), .B(n493), .Z(n519) );
  NAND2_X1 U555 ( .A1(n494), .A2(n519), .ZN(n495) );
  NOR2_X1 U556 ( .A1(n571), .A2(n504), .ZN(n499) );
  XOR2_X1 U557 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n497) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U561 ( .A1(n521), .A2(n504), .ZN(n500) );
  XOR2_X1 U562 ( .A(KEYINPUT108), .B(n500), .Z(n501) );
  XNOR2_X1 U563 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  NOR2_X1 U564 ( .A1(n504), .A2(n532), .ZN(n502) );
  XOR2_X1 U565 ( .A(KEYINPUT40), .B(n502), .Z(n503) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NOR2_X1 U567 ( .A1(n525), .A2(n504), .ZN(n505) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n505), .Z(G1331GAT) );
  INV_X1 U569 ( .A(n506), .ZN(n557) );
  NOR2_X1 U570 ( .A1(n575), .A2(n557), .ZN(n518) );
  NAND2_X1 U571 ( .A1(n518), .A2(n507), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n571), .A2(n514), .ZN(n508) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n508), .Z(n509) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n509), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n521), .A2(n514), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1333GAT) );
  NOR2_X1 U578 ( .A1(n532), .A2(n514), .ZN(n512) );
  XOR2_X1 U579 ( .A(KEYINPUT110), .B(n512), .Z(n513) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  NOR2_X1 U581 ( .A1(n525), .A2(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U584 ( .A(G78GAT), .B(n517), .Z(G1335GAT) );
  NAND2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n524) );
  NOR2_X1 U586 ( .A1(n571), .A2(n524), .ZN(n520) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n520), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n521), .A2(n524), .ZN(n522) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n532), .A2(n524), .ZN(n523) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n523), .Z(G1338GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U595 ( .A(G106GAT), .B(n528), .Z(G1339GAT) );
  XOR2_X1 U596 ( .A(n530), .B(n529), .Z(n552) );
  INV_X1 U597 ( .A(n552), .ZN(n531) );
  NOR2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n540) );
  NOR2_X1 U600 ( .A1(n553), .A2(n540), .ZN(n535) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n535), .Z(n536) );
  XNOR2_X1 U602 ( .A(KEYINPUT116), .B(n536), .ZN(G1340GAT) );
  NOR2_X1 U603 ( .A1(n557), .A2(n540), .ZN(n538) );
  XNOR2_X1 U604 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U606 ( .A(G120GAT), .B(n539), .Z(G1341GAT) );
  INV_X1 U607 ( .A(n540), .ZN(n546) );
  NAND2_X1 U608 ( .A1(n569), .A2(n546), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XOR2_X1 U610 ( .A(n542), .B(KEYINPUT119), .Z(n544) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(KEYINPUT118), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  INV_X1 U616 ( .A(n549), .ZN(n573) );
  NOR2_X1 U617 ( .A1(n573), .A2(n550), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n564) );
  NOR2_X1 U619 ( .A1(n553), .A2(n564), .ZN(n554) );
  XOR2_X1 U620 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n556) );
  XNOR2_X1 U622 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n561) );
  NOR2_X1 U624 ( .A1(n557), .A2(n564), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  INV_X1 U628 ( .A(n582), .ZN(n562) );
  NOR2_X1 U629 ( .A1(n562), .A2(n564), .ZN(n563) );
  XOR2_X1 U630 ( .A(G155GAT), .B(n563), .Z(G1346GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(G162GAT), .B(n566), .Z(G1347GAT) );
  NAND2_X1 U633 ( .A1(n575), .A2(n568), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G169GAT), .B(n567), .ZN(G1348GAT) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT126), .ZN(n579) );
  XOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .Z(n577) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n574) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n585) );
  NAND2_X1 U641 ( .A1(n585), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  NAND2_X1 U645 ( .A1(n585), .A2(n388), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n585), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

