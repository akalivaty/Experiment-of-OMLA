//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008;
  NOR2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR3_X1   g006(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n203), .B(new_n204), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n203), .A2(KEYINPUT76), .A3(new_n204), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n211));
  INV_X1    g010(.A(new_n204), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(new_n202), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n216));
  XOR2_X1   g015(.A(G155gat), .B(G162gat), .Z(new_n217));
  AND3_X1   g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n215), .B2(new_n217), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n209), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G113gat), .B(G120gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT70), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G127gat), .B(G134gat), .Z(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n222), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n224), .B(KEYINPUT69), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n224), .B1(KEYINPUT1), .B2(new_n221), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n220), .B(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G225gat), .A2(G233gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT39), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n209), .ZN(new_n239));
  INV_X1    g038(.A(new_n219), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n232), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(KEYINPUT4), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n220), .B2(new_n232), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT78), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n232), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n251), .B(new_n209), .C1(new_n218), .C2(new_n219), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n248), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n243), .B1(new_n220), .B2(KEYINPUT3), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(KEYINPUT78), .A3(new_n252), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n247), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n238), .B1(new_n257), .B2(new_n234), .ZN(new_n258));
  XNOR2_X1  g057(.A(G1gat), .B(G29gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT0), .ZN(new_n260));
  XNOR2_X1  g059(.A(G57gat), .B(G85gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n260), .B(new_n261), .Z(new_n262));
  INV_X1    g061(.A(new_n247), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n255), .A2(KEYINPUT78), .A3(new_n252), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT78), .B1(new_n255), .B2(new_n252), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(new_n237), .A3(new_n235), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n258), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT40), .ZN(new_n269));
  INV_X1    g068(.A(new_n262), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n256), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n234), .A4(new_n263), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT79), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n234), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n272), .B1(new_n233), .B2(new_n235), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n273), .A2(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n274), .A3(new_n276), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n270), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT67), .B(G190gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n284));
  OR2_X1    g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n283), .A2(new_n284), .B1(G183gat), .B2(G190gat), .ZN(new_n286));
  OR3_X1    g085(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT23), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n294), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n295), .A3(new_n288), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT66), .ZN(new_n297));
  AND3_X1   g096(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(KEYINPUT64), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n300));
  INV_X1    g099(.A(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(G190gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(KEYINPUT64), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n299), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(KEYINPUT25), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n297), .B(new_n305), .C1(new_n296), .C2(new_n307), .ZN(new_n308));
  AOI211_X1 g107(.A(new_n298), .B(new_n300), .C1(new_n281), .C2(new_n301), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT25), .B1(new_n309), .B2(new_n296), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n291), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n311), .A2(G226gat), .A3(G233gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n311), .A2(new_n313), .B1(G226gat), .B2(G233gat), .ZN(new_n314));
  XOR2_X1   g113(.A(G211gat), .B(G218gat), .Z(new_n315));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G211gat), .B(G218gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322));
  INV_X1    g121(.A(G211gat), .ZN(new_n323));
  INV_X1    g122(.A(G218gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n317), .A2(new_n325), .A3(new_n321), .A4(new_n319), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n312), .A2(new_n314), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n312), .B2(new_n314), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G8gat), .B(G36gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(G64gat), .B(G92gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n337), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(new_n332), .B2(new_n333), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT30), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n337), .B(KEYINPUT75), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n332), .A2(new_n333), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n269), .A2(KEYINPUT83), .A3(new_n280), .A4(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT40), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n266), .A2(new_n235), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n270), .B1(new_n349), .B2(new_n238), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n348), .B1(new_n350), .B2(new_n267), .ZN(new_n351));
  AND4_X1   g150(.A1(new_n348), .A2(new_n258), .A3(new_n262), .A4(new_n267), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n280), .B(new_n346), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT83), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n347), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT38), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n332), .A2(new_n333), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT37), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT37), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n334), .A2(new_n360), .ZN(new_n361));
  AND4_X1   g160(.A1(new_n357), .A2(new_n359), .A3(new_n361), .A4(new_n344), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n337), .B1(new_n334), .B2(new_n360), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n357), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n362), .A2(new_n364), .A3(new_n342), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n274), .B1(new_n275), .B2(KEYINPUT5), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n275), .A2(new_n276), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(new_n262), .A3(new_n278), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n280), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(KEYINPUT6), .B(new_n270), .C1(new_n277), .C2(new_n279), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n372), .A2(KEYINPUT84), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(KEYINPUT84), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n365), .B(new_n371), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376));
  INV_X1    g175(.A(G50gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(G22gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n327), .A2(new_n313), .A3(new_n328), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n382), .A2(new_n251), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n381), .B1(new_n383), .B2(new_n242), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n330), .B1(new_n252), .B2(new_n313), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT3), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n327), .A2(KEYINPUT81), .A3(new_n313), .A4(new_n328), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n242), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(G228gat), .B(G233gat), .C1(new_n390), .C2(new_n385), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n386), .B2(new_n391), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n396), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n386), .A2(new_n391), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT82), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n400), .B2(new_n393), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n380), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n396), .B1(new_n394), .B2(new_n395), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(new_n393), .A3(new_n398), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n379), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n356), .A2(new_n375), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n311), .A2(new_n243), .ZN(new_n408));
  INV_X1    g207(.A(G227gat), .ZN(new_n409));
  INV_X1    g208(.A(G233gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n232), .A2(new_n291), .A3(new_n308), .A4(new_n310), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n408), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT71), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT71), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n408), .A2(new_n415), .A3(new_n411), .A4(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n408), .A2(new_n412), .ZN(new_n418));
  INV_X1    g217(.A(new_n411), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(KEYINPUT32), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT32), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n418), .B(new_n419), .C1(new_n415), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT34), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT72), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(new_n419), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT73), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n417), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G15gat), .B(G43gat), .Z(new_n432));
  XNOR2_X1  g231(.A(G71gat), .B(G99gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n429), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT33), .B1(new_n414), .B2(new_n416), .ZN(new_n436));
  INV_X1    g235(.A(new_n434), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n436), .A2(new_n428), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n424), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n431), .A2(new_n429), .A3(new_n434), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n428), .B1(new_n436), .B2(new_n437), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n423), .A4(new_n421), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT36), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n371), .A2(new_n372), .ZN(new_n446));
  INV_X1    g245(.A(new_n346), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n402), .A2(new_n405), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n407), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n446), .A2(new_n406), .A3(new_n447), .A4(new_n443), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n453));
  INV_X1    g252(.A(new_n343), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n345), .B1(new_n342), .B2(KEYINPUT30), .ZN(new_n455));
  XNOR2_X1  g254(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n402), .A3(new_n405), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n439), .A2(KEYINPUT85), .A3(new_n442), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT85), .B1(new_n439), .B2(new_n442), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n453), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n451), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G113gat), .B(G141gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(G169gat), .B(G197gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n468), .A2(new_n470), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT12), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT12), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n471), .B2(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G29gat), .ZN(new_n478));
  INV_X1    g277(.A(G36gat), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT14), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT14), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(G29gat), .B2(G36gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(G29gat), .A2(G36gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(G43gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(G50gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n377), .A2(G43gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT15), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n484), .B(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT15), .ZN(new_n490));
  OR2_X1    g289(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n492));
  AOI21_X1  g291(.A(G50gat), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT89), .B1(new_n377), .B2(G43gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(new_n485), .A3(G50gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n490), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT17), .B1(new_n489), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G1gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT16), .ZN(new_n502));
  INV_X1    g301(.A(G15gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G22gat), .ZN(new_n504));
  INV_X1    g303(.A(G22gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G15gat), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(G1gat), .B1(new_n504), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g307(.A(G8gat), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n506), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n501), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n512));
  INV_X1    g311(.A(G8gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n490), .B1(new_n485), .B2(G50gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n484), .A2(new_n487), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n488), .A2(new_n482), .A3(new_n483), .A4(new_n480), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n498), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n500), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n493), .ZN(new_n525));
  INV_X1    g324(.A(new_n497), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n527), .A2(new_n490), .B1(new_n518), .B2(new_n519), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n515), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n523), .A2(KEYINPUT18), .A3(new_n524), .A4(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n524), .B(KEYINPUT13), .Z(new_n531));
  INV_X1    g330(.A(new_n529), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n528), .A2(new_n515), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n477), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n522), .A2(new_n516), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n521), .B1(new_n520), .B2(new_n498), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n524), .B(new_n529), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT90), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT90), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n523), .A2(new_n541), .A3(new_n524), .A4(new_n529), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT92), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n535), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(new_n535), .B2(new_n543), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n534), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n543), .B2(KEYINPUT91), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT91), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n539), .A2(new_n550), .A3(new_n540), .A4(new_n542), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n477), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555));
  INV_X1    g354(.A(G57gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(G64gat), .ZN(new_n557));
  INV_X1    g356(.A(G64gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT93), .A3(G57gat), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n557), .B(new_n559), .C1(G57gat), .C2(new_n558), .ZN(new_n560));
  NAND2_X1  g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  OR2_X1    g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT9), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n556), .A2(G64gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n558), .A2(G57gat), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT9), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n562), .A2(new_n561), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G127gat), .ZN(new_n576));
  XOR2_X1   g375(.A(G183gat), .B(G211gat), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n516), .B1(new_n572), .B2(new_n571), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT94), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G155gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n583), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n579), .A2(new_n580), .A3(new_n586), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT95), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT41), .ZN(new_n593));
  OR2_X1    g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(KEYINPUT97), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n597));
  AND2_X1   g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(G92gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n595), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(KEYINPUT96), .A2(G99gat), .A3(G106gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(KEYINPUT8), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n601), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT7), .ZN(new_n614));
  INV_X1    g413(.A(G85gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(G92gat), .A3(new_n604), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT8), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n618), .B1(new_n595), .B2(new_n608), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n617), .A2(new_n603), .B1(new_n619), .B2(new_n610), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n596), .A2(new_n600), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n613), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n520), .A2(new_n498), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n593), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n500), .A2(new_n522), .A3(new_n623), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT99), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n592), .A2(KEYINPUT41), .ZN(new_n633));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  INV_X1    g434(.A(new_n631), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n625), .A2(new_n626), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n528), .A2(new_n622), .A3(new_n613), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT98), .B1(new_n638), .B2(new_n593), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n636), .B(new_n628), .C1(new_n637), .C2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n632), .A2(new_n635), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n635), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n636), .B1(new_n627), .B2(new_n628), .ZN(new_n643));
  INV_X1    g442(.A(new_n640), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n590), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n601), .B2(new_n612), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n564), .A2(new_n560), .B1(new_n568), .B2(new_n569), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n601), .A2(new_n612), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n620), .A2(new_n621), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n622), .B(new_n613), .C1(new_n571), .C2(new_n649), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT10), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n623), .A2(new_n657), .A3(new_n571), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n648), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n655), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n648), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT101), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n665), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n647), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n465), .A2(new_n554), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n446), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(new_n501), .ZN(G1324gat));
  INV_X1    g472(.A(new_n671), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n346), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n674), .A2(KEYINPUT42), .A3(new_n346), .A4(new_n675), .ZN(new_n679));
  OAI21_X1  g478(.A(G8gat), .B1(new_n671), .B2(new_n447), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n678), .A2(KEYINPUT102), .A3(new_n679), .A4(new_n680), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(G1325gat));
  XNOR2_X1  g484(.A(new_n443), .B(KEYINPUT36), .ZN(new_n686));
  OAI21_X1  g485(.A(G15gat), .B1(new_n671), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n459), .A2(new_n460), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n503), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n671), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n671), .A2(new_n406), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  AOI22_X1  g492(.A1(new_n407), .A2(new_n450), .B1(new_n453), .B2(new_n463), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n590), .A2(new_n669), .ZN(new_n695));
  INV_X1    g494(.A(new_n646), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n694), .A2(new_n553), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n446), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n478), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n694), .B2(new_n646), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n346), .B1(new_n371), .B2(new_n372), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n686), .B1(new_n704), .B2(new_n406), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n449), .B1(new_n347), .B2(new_n355), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n375), .B2(new_n706), .ZN(new_n707));
  AOI22_X1  g506(.A1(KEYINPUT35), .A2(new_n452), .B1(new_n461), .B2(new_n462), .ZN(new_n708));
  OAI211_X1 g507(.A(KEYINPUT44), .B(new_n696), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n703), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT103), .B1(new_n547), .B2(new_n552), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n543), .A2(KEYINPUT91), .ZN(new_n712));
  INV_X1    g511(.A(new_n548), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n713), .A3(new_n551), .ZN(new_n714));
  INV_X1    g513(.A(new_n477), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n535), .A2(new_n543), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT92), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n535), .A2(new_n543), .A3(new_n544), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n716), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n711), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n723), .A2(new_n590), .A3(new_n669), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n710), .A2(new_n699), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n701), .B1(new_n478), .B2(new_n725), .ZN(G1328gat));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n465), .A2(new_n554), .A3(new_n696), .A4(new_n695), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n447), .A2(G36gat), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT104), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n698), .A2(new_n732), .A3(new_n729), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n727), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n731), .A2(new_n733), .A3(new_n727), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n710), .A2(new_n346), .A3(new_n724), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G36gat), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n735), .A2(new_n736), .A3(new_n737), .A4(new_n739), .ZN(G1329gat));
  NAND2_X1  g539(.A1(new_n491), .A2(new_n492), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n698), .B2(new_n688), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(KEYINPUT47), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n710), .A2(new_n445), .A3(new_n741), .A4(new_n724), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1330gat));
  NAND4_X1  g548(.A1(new_n703), .A2(new_n449), .A3(new_n709), .A4(new_n724), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G50gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n698), .A2(new_n377), .A3(new_n449), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1331gat));
  AND2_X1   g554(.A1(new_n711), .A2(new_n722), .ZN(new_n756));
  INV_X1    g555(.A(new_n669), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n756), .A2(new_n647), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n465), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n446), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(new_n556), .ZN(G1332gat));
  XNOR2_X1  g560(.A(new_n759), .B(KEYINPUT107), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n346), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT49), .B(G64gat), .Z(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n763), .B2(new_n765), .ZN(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n686), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n688), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n759), .B2(new_n770), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n769), .A2(KEYINPUT50), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT50), .B1(new_n769), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n762), .A2(new_n449), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g575(.A1(new_n756), .A2(new_n590), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n696), .B(new_n777), .C1(new_n707), .C2(new_n708), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n465), .A2(KEYINPUT51), .A3(new_n696), .A4(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n782), .A2(new_n615), .A3(new_n699), .A4(new_n669), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n756), .A2(new_n590), .A3(new_n757), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n703), .A2(new_n699), .A3(new_n709), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G85gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT108), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n783), .A2(new_n789), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1336gat));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n780), .A2(new_n792), .A3(new_n781), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n778), .A2(KEYINPUT110), .A3(new_n779), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n447), .A2(G92gat), .A3(new_n757), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n703), .A2(new_n346), .A3(new_n709), .A4(new_n784), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(KEYINPUT109), .A3(G92gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT109), .B1(new_n797), .B2(G92gat), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT52), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(new_n797), .B2(G92gat), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n782), .A2(KEYINPUT111), .A3(new_n795), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT111), .B1(new_n782), .B2(new_n795), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n801), .A2(new_n805), .ZN(G1337gat));
  NAND3_X1  g605(.A1(new_n710), .A2(new_n445), .A3(new_n784), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G99gat), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n770), .A2(G99gat), .A3(new_n757), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT112), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n782), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(G1338gat));
  NOR3_X1   g611(.A1(new_n406), .A2(G106gat), .A3(new_n757), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n793), .A2(new_n794), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n703), .A2(new_n449), .A3(new_n709), .A4(new_n784), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G106gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT53), .B1(new_n782), .B2(new_n813), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n816), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1339gat));
  NOR3_X1   g620(.A1(new_n756), .A2(new_n647), .A3(new_n669), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT113), .ZN(new_n823));
  INV_X1    g622(.A(new_n590), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n524), .B1(new_n523), .B2(new_n529), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n532), .A2(new_n533), .A3(new_n531), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n473), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n545), .B2(new_n546), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n646), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n830), .B(new_n648), .C1(new_n656), .C2(new_n658), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n665), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(KEYINPUT114), .A3(new_n665), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n660), .A2(new_n657), .ZN(new_n837));
  INV_X1    g636(.A(new_n658), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n837), .A2(G230gat), .A3(G233gat), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(KEYINPUT54), .A3(new_n659), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n837), .A2(new_n838), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n830), .B1(new_n844), .B2(new_n648), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n842), .B1(new_n845), .B2(new_n839), .ZN(new_n846));
  AOI211_X1 g645(.A(KEYINPUT115), .B(new_n666), .C1(new_n836), .C2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n831), .A2(KEYINPUT114), .A3(new_n665), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT114), .B1(new_n831), .B2(new_n665), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT55), .B(new_n840), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n848), .B1(new_n851), .B2(new_n667), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n829), .B(new_n843), .C1(new_n847), .C2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n828), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n669), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n843), .B1(new_n847), .B2(new_n852), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n723), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n854), .B1(new_n858), .B2(new_n646), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n824), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI211_X1 g660(.A(KEYINPUT116), .B(new_n854), .C1(new_n858), .C2(new_n646), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n823), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n863), .A2(new_n699), .ZN(new_n864));
  INV_X1    g663(.A(new_n443), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n449), .A2(new_n865), .A3(new_n346), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(G113gat), .B1(new_n867), .B2(new_n756), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n863), .A2(new_n406), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n699), .A2(new_n447), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n869), .A2(new_n770), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n554), .A2(G113gat), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(G1340gat));
  AOI21_X1  g672(.A(G120gat), .B1(new_n867), .B2(new_n669), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n669), .A2(G120gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n871), .B2(new_n875), .ZN(G1341gat));
  NAND2_X1  g675(.A1(new_n867), .A2(new_n590), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(KEYINPUT117), .ZN(new_n878));
  AOI21_X1  g677(.A(G127gat), .B1(new_n877), .B2(KEYINPUT117), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n590), .A2(G127gat), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n878), .A2(new_n879), .B1(new_n871), .B2(new_n880), .ZN(G1342gat));
  INV_X1    g680(.A(G134gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n882), .A3(new_n696), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n871), .A2(new_n696), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n884), .B(new_n885), .C1(new_n882), .C2(new_n886), .ZN(G1343gat));
  NOR2_X1   g686(.A1(new_n870), .A2(new_n445), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT118), .Z(new_n889));
  AOI21_X1  g688(.A(KEYINPUT57), .B1(new_n863), .B2(new_n449), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n666), .B1(new_n836), .B2(new_n846), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n843), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n553), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n843), .A2(KEYINPUT119), .A3(new_n892), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n895), .A2(new_n896), .B1(new_n669), .B2(new_n855), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n853), .B1(new_n897), .B2(new_n696), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n824), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n891), .B(new_n406), .C1(new_n899), .C2(new_n823), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n889), .B1(new_n890), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G141gat), .B1(new_n901), .B2(new_n553), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n863), .A2(new_n699), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n686), .A2(new_n449), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n903), .A2(new_n346), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(G141gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n906), .A3(new_n554), .ZN(new_n907));
  XNOR2_X1  g706(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n902), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G141gat), .B1(new_n901), .B2(new_n723), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(new_n907), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(G1344gat));
  NAND2_X1  g712(.A1(new_n905), .A2(new_n669), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT59), .ZN(new_n915));
  INV_X1    g714(.A(G148gat), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n901), .A2(KEYINPUT59), .A3(new_n757), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n898), .A2(new_n824), .B1(new_n553), .B2(new_n670), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n449), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n919), .A2(new_n920), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n891), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n406), .A2(new_n891), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n863), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(new_n669), .A3(new_n889), .ZN(new_n928));
  NAND2_X1  g727(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n917), .B(new_n918), .C1(new_n928), .C2(new_n929), .ZN(G1345gat));
  OAI21_X1  g729(.A(G155gat), .B1(new_n901), .B2(new_n824), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n905), .A2(new_n205), .A3(new_n590), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1346gat));
  OAI21_X1  g732(.A(G162gat), .B1(new_n901), .B2(new_n646), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n905), .A2(new_n206), .A3(new_n696), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n699), .A2(new_n447), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n938), .A2(new_n770), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n863), .A2(new_n406), .A3(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(G169gat), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n940), .A2(new_n941), .A3(new_n553), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n863), .A2(new_n446), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n449), .A2(new_n865), .A3(new_n447), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n756), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n942), .B1(new_n947), .B2(new_n941), .ZN(G1348gat));
  OAI21_X1  g747(.A(G176gat), .B1(new_n940), .B2(new_n757), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n757), .A2(G176gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n945), .B2(new_n950), .ZN(G1349gat));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n863), .A2(new_n406), .A3(new_n590), .A4(new_n939), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G183gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n590), .A2(new_n282), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n863), .A2(new_n446), .A3(new_n944), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n954), .A2(KEYINPUT122), .A3(new_n957), .ZN(new_n961));
  AND4_X1   g760(.A1(new_n952), .A2(new_n960), .A3(KEYINPUT60), .A4(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT60), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n954), .A2(new_n963), .A3(new_n957), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT123), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n963), .B1(new_n958), .B2(new_n959), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n961), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n962), .A2(new_n967), .ZN(G1350gat));
  NAND3_X1  g767(.A1(new_n946), .A2(new_n281), .A3(new_n696), .ZN(new_n969));
  OAI21_X1  g768(.A(G190gat), .B1(new_n940), .B2(new_n646), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n970), .A2(KEYINPUT61), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n970), .A2(KEYINPUT61), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1351gat));
  NOR2_X1   g772(.A1(new_n938), .A2(new_n445), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n927), .A2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(G197gat), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n975), .A2(new_n976), .A3(new_n553), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n904), .A2(new_n447), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n943), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(G197gat), .B1(new_n979), .B2(new_n756), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n977), .A2(new_n980), .ZN(G1352gat));
  INV_X1    g780(.A(new_n923), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n406), .B1(new_n919), .B2(new_n920), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT57), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(new_n926), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n669), .B(new_n974), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT126), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n927), .A2(new_n988), .A3(new_n669), .A4(new_n974), .ZN(new_n989));
  XNOR2_X1  g788(.A(KEYINPUT124), .B(G204gat), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n992));
  AOI211_X1 g791(.A(new_n990), .B(new_n757), .C1(new_n992), .C2(KEYINPUT62), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n979), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n991), .A2(new_n996), .ZN(G1353gat));
  OAI211_X1 g796(.A(new_n590), .B(new_n974), .C1(new_n984), .C2(new_n985), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(G211gat), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(KEYINPUT63), .ZN(new_n1000));
  AND4_X1   g799(.A1(new_n323), .A2(new_n943), .A3(new_n590), .A4(new_n978), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT63), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n998), .A2(new_n1004), .A3(G211gat), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1000), .A2(new_n1003), .A3(new_n1005), .ZN(G1354gat));
  OAI21_X1  g805(.A(G218gat), .B1(new_n975), .B2(new_n646), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n979), .A2(new_n324), .A3(new_n696), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n1008), .ZN(G1355gat));
endmodule


