//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(G125), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n464), .A2(KEYINPUT65), .A3(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT65), .B1(new_n464), .B2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G101), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n465), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n468), .A2(G136), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT66), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G124), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n476), .A2(new_n481), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n483));
  NAND2_X1  g058(.A1(G126), .A2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n466), .B2(new_n467), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n464), .A2(G114), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n483), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(G2104), .ZN(new_n493));
  AND2_X1   g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n497), .A3(KEYINPUT67), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n464), .C1(new_n495), .C2(new_n496), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n462), .A2(new_n501), .A3(G138), .A4(new_n464), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n489), .A2(new_n498), .B1(new_n500), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n505), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G62), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n512), .A2(new_n513), .B1(G75), .B2(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n511), .A2(KEYINPUT70), .A3(G62), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n504), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  INV_X1    g092(.A(new_n506), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n505), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n519));
  AOI21_X1  g094(.A(KEYINPUT69), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n517), .B(new_n518), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G88), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n526), .B2(G50), .ZN(new_n527));
  INV_X1    g102(.A(G50), .ZN(new_n528));
  NOR3_X1   g103(.A1(new_n525), .A2(KEYINPUT68), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n523), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n516), .A2(new_n530), .ZN(G166));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n511), .B(new_n532), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n533), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  INV_X1    g111(.A(G51), .ZN(new_n537));
  INV_X1    g112(.A(G89), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n536), .B1(new_n525), .B2(new_n537), .C1(new_n521), .C2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n534), .A2(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(new_n509), .A2(new_n510), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(new_n518), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(new_n532), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n511), .A2(KEYINPUT71), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n543), .A2(G64), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n504), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n522), .A2(G90), .B1(G52), .B2(new_n526), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(G171));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n521), .A2(new_n551), .B1(new_n552), .B2(new_n525), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n533), .A2(G56), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n553), .B1(new_n556), .B2(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND3_X1  g138(.A1(new_n517), .A2(G53), .A3(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(KEYINPUT74), .B(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n542), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n565), .A2(new_n566), .B1(new_n569), .B2(G651), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n521), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n511), .A2(KEYINPUT73), .A3(new_n517), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(G91), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  OR2_X1    g151(.A1(new_n534), .A2(new_n539), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND3_X1  g153(.A1(new_n572), .A2(G87), .A3(new_n573), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n526), .A2(G49), .ZN(new_n580));
  AOI21_X1  g155(.A(G74), .B1(new_n543), .B2(new_n544), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n504), .ZN(G288));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n542), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n572), .A2(G86), .A3(new_n573), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT75), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n572), .A2(new_n589), .A3(G86), .A4(new_n573), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n526), .A2(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  NAND3_X1  g168(.A1(new_n543), .A2(G60), .A3(new_n544), .ZN(new_n594));
  AND2_X1   g169(.A1(G72), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(KEYINPUT76), .B1(new_n594), .B2(new_n596), .ZN(new_n600));
  NOR3_X1   g175(.A1(new_n599), .A2(new_n504), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n521), .A2(new_n602), .B1(new_n603), .B2(new_n525), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT77), .Z(new_n605));
  NOR2_X1   g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  OR3_X1    g183(.A1(G171), .A2(KEYINPUT78), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT78), .B1(G171), .B2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n526), .A2(G54), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n504), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n572), .A2(G92), .A3(new_n573), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n572), .A2(KEYINPUT10), .A3(G92), .A4(new_n573), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n609), .B(new_n610), .C1(G868), .C2(new_n618), .ZN(G284));
  OAI211_X1 g194(.A(new_n609), .B(new_n610), .C1(G868), .C2(new_n618), .ZN(G321));
  NAND2_X1  g195(.A1(G299), .A2(new_n608), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G168), .B2(new_n608), .ZN(G280));
  XNOR2_X1  g197(.A(G280), .B(KEYINPUT79), .ZN(G297));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n618), .B1(new_n624), .B2(G860), .ZN(G148));
  AOI21_X1  g200(.A(new_n504), .B1(new_n554), .B2(new_n555), .ZN(new_n626));
  NOR3_X1   g201(.A1(new_n626), .A2(G868), .A3(new_n553), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n618), .A2(new_n624), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT80), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n627), .B1(new_n629), .B2(G868), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g206(.A1(new_n470), .A2(new_n471), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(new_n462), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n468), .A2(G135), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n480), .A2(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n464), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n637), .A2(new_n638), .A3(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2430), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n654), .A2(KEYINPUT82), .A3(new_n655), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n652), .A2(new_n653), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n650), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  AOI211_X1 g238(.A(new_n661), .B(new_n649), .C1(new_n658), .C2(new_n659), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n648), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n659), .ZN(new_n668));
  AOI21_X1  g243(.A(KEYINPUT82), .B1(new_n654), .B2(new_n655), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n662), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(new_n649), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n660), .A2(new_n662), .A3(new_n650), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(new_n672), .A3(new_n647), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n665), .A2(new_n667), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT83), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n676));
  NAND4_X1  g251(.A1(new_n665), .A2(new_n676), .A3(new_n673), .A4(new_n667), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G14), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n665), .A2(new_n673), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n666), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(G401));
  XOR2_X1   g257(.A(KEYINPUT84), .B(KEYINPUT17), .Z(new_n683));
  XNOR2_X1  g258(.A(G2072), .B(G2078), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2067), .B(G2678), .ZN(new_n686));
  XOR2_X1   g261(.A(G2084), .B(G2090), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n685), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n686), .B2(new_n684), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n685), .B2(new_n686), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n687), .A2(new_n686), .A3(new_n684), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT18), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n689), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G2096), .B(G2100), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G227));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1956), .B(G2474), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1961), .B(G1966), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n700), .A2(new_n701), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n699), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n699), .A2(new_n706), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(G1991), .B(G1996), .Z(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n714), .A2(new_n717), .A3(new_n715), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(G229));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT87), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(KEYINPUT87), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n606), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(G24), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G1986), .ZN(new_n730));
  INV_X1    g305(.A(G1986), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n727), .A2(new_n731), .A3(new_n728), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n468), .A2(G131), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n480), .A2(G119), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n464), .A2(G107), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n734), .B(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  MUX2_X1   g313(.A(G25), .B(new_n738), .S(G29), .Z(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n739), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n733), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n723), .B1(new_n591), .B2(new_n592), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n723), .A2(G6), .ZN(new_n748));
  OR3_X1    g323(.A1(new_n747), .A2(KEYINPUT89), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT32), .B(G1981), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT89), .B1(new_n747), .B2(new_n748), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(G166), .A2(new_n726), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G22), .B2(new_n726), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G1971), .ZN(new_n755));
  INV_X1    g330(.A(G1971), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n753), .B(new_n756), .C1(G22), .C2(new_n726), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n723), .A2(G23), .ZN(new_n758));
  INV_X1    g333(.A(G288), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n723), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT33), .B(G1976), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT90), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n762), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n758), .B(new_n764), .C1(new_n759), .C2(new_n723), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n755), .A2(new_n757), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n752), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n750), .B1(new_n749), .B2(new_n751), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n746), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n768), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n770), .A2(new_n752), .A3(new_n766), .A4(new_n745), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n744), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT36), .ZN(new_n773));
  AOI21_X1  g348(.A(KEYINPUT92), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(KEYINPUT91), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(KEYINPUT36), .B1(new_n772), .B2(KEYINPUT91), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n772), .A2(KEYINPUT91), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n779), .A2(new_n775), .A3(KEYINPUT92), .A4(KEYINPUT36), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n723), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n723), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G1966), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT95), .Z(new_n784));
  NOR2_X1   g359(.A1(G171), .A2(new_n723), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G5), .B2(new_n723), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G1961), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT31), .B(G11), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n790), .A2(G28), .ZN(new_n791));
  INV_X1    g366(.A(G29), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n790), .B2(G28), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n789), .B1(new_n791), .B2(new_n793), .C1(new_n643), .C2(new_n792), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n782), .B2(G1966), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n784), .A2(new_n788), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT96), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n723), .A2(G4), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n618), .B2(new_n723), .ZN(new_n799));
  INV_X1    g374(.A(G1348), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(G29), .A2(G33), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT93), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n468), .A2(G139), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT94), .Z(new_n805));
  NAND3_X1  g380(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT25), .Z(new_n807));
  AOI22_X1  g382(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n805), .B(new_n807), .C1(new_n464), .C2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n803), .B1(new_n809), .B2(new_n792), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(G2072), .Z(new_n811));
  NAND3_X1  g386(.A1(new_n724), .A2(G20), .A3(new_n725), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT23), .Z(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G299), .B2(G16), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(G1956), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n792), .A2(G32), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n632), .A2(G105), .B1(G141), .B2(new_n468), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n480), .A2(G129), .ZN(new_n818));
  NAND3_X1  g393(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT26), .Z(new_n820));
  AND3_X1   g395(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n816), .B1(new_n821), .B2(new_n792), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT27), .B(G1996), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT24), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n792), .B1(new_n826), .B2(G34), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n826), .B2(G34), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G160), .B2(G29), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(G2084), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n822), .A2(new_n824), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(G2084), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n825), .A2(new_n830), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(G164), .A2(new_n792), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G27), .B2(new_n792), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT97), .B(G2078), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n792), .A2(G26), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT28), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n468), .A2(G140), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n480), .A2(G128), .ZN(new_n841));
  OR2_X1    g416(.A1(G104), .A2(G2105), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n842), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n839), .B1(new_n845), .B2(new_n792), .ZN(new_n846));
  INV_X1    g421(.A(G2067), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n835), .A2(new_n836), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n837), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR4_X1   g425(.A1(new_n811), .A2(new_n815), .A3(new_n833), .A4(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G19), .ZN(new_n852));
  MUX2_X1   g427(.A(new_n852), .B(new_n557), .S(new_n726), .Z(new_n853));
  INV_X1    g428(.A(G1341), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n787), .A2(G1961), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(G29), .A2(G35), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(G162), .B2(G29), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT29), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G2090), .ZN(new_n859));
  AOI211_X1 g434(.A(new_n855), .B(new_n859), .C1(new_n854), .C2(new_n853), .ZN(new_n860));
  AND4_X1   g435(.A1(new_n797), .A2(new_n801), .A3(new_n851), .A4(new_n860), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n778), .A2(new_n780), .A3(new_n861), .ZN(G311));
  NAND3_X1  g437(.A1(new_n778), .A2(new_n780), .A3(new_n861), .ZN(G150));
  NAND2_X1  g438(.A1(new_n618), .A2(G559), .ZN(new_n864));
  XOR2_X1   g439(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n543), .A2(G67), .A3(new_n544), .ZN(new_n867));
  NAND2_X1  g442(.A1(G80), .A2(G543), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n504), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G93), .ZN(new_n870));
  INV_X1    g445(.A(G55), .ZN(new_n871));
  OAI22_X1  g446(.A1(new_n521), .A2(new_n870), .B1(new_n871), .B2(new_n525), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n557), .A2(new_n873), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n626), .A2(new_n553), .B1(new_n869), .B2(new_n872), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n866), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n878));
  AOI21_X1  g453(.A(G860), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT99), .ZN(new_n881));
  INV_X1    g456(.A(new_n873), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G860), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT37), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(G145));
  NAND2_X1  g460(.A1(new_n493), .A2(new_n497), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(new_n500), .B2(new_n502), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n844), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n888), .A2(new_n821), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n809), .A2(KEYINPUT101), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n821), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n809), .A2(KEYINPUT101), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n892), .B(new_n893), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n480), .A2(G130), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n464), .A2(G118), .ZN(new_n896));
  OAI21_X1  g471(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(G142), .B2(new_n468), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n634), .B(new_n899), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n738), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n894), .B(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(G162), .B(new_n643), .Z(new_n903));
  XOR2_X1   g478(.A(G160), .B(KEYINPUT100), .Z(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n894), .A2(new_n901), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n894), .A2(new_n901), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT40), .Z(G395));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n876), .B(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(new_n629), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n618), .B2(G299), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n616), .A2(new_n617), .ZN(new_n919));
  INV_X1    g494(.A(new_n613), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G299), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT104), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n618), .A2(KEYINPUT103), .A3(G299), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT103), .B1(new_n618), .B2(G299), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n918), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n916), .A2(new_n927), .ZN(new_n928));
  XOR2_X1   g503(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n929));
  NOR2_X1   g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n923), .A2(new_n918), .ZN(new_n931));
  INV_X1    g506(.A(new_n925), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n618), .A2(KEYINPUT103), .A3(G299), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT41), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n916), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n592), .B(new_n591), .C1(new_n601), .C2(new_n605), .ZN(new_n937));
  INV_X1    g512(.A(new_n605), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n600), .A2(new_n504), .ZN(new_n939));
  OAI211_X1 g514(.A(G305), .B(new_n938), .C1(new_n599), .C2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n941));
  NOR2_X1   g516(.A1(G288), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G288), .A2(new_n941), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(G303), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(G166), .B1(new_n946), .B2(new_n942), .ZN(new_n947));
  AND4_X1   g522(.A1(new_n937), .A2(new_n940), .A3(new_n945), .A4(new_n947), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n937), .A2(new_n940), .B1(new_n947), .B2(new_n945), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n953));
  AND4_X1   g528(.A1(new_n928), .A2(new_n936), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n928), .A2(new_n936), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  OAI21_X1  g530(.A(G868), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n882), .A2(new_n608), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(G295));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n957), .ZN(G331));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  NAND2_X1  g535(.A1(G171), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT107), .B1(new_n547), .B2(new_n549), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(G286), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(G168), .A2(G171), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n876), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n963), .A2(new_n964), .A3(new_n875), .A4(new_n874), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n935), .B2(new_n930), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n874), .A2(new_n875), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n964), .A4(new_n963), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n970), .A2(new_n973), .A3(new_n926), .A4(new_n966), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n951), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n969), .A2(new_n950), .A3(new_n974), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n908), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n929), .B1(new_n931), .B2(new_n934), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n926), .A2(KEYINPUT41), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n970), .A2(new_n973), .A3(new_n966), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n966), .A2(new_n926), .A3(new_n967), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n951), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n908), .A4(new_n977), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n979), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n985), .B1(new_n982), .B2(new_n983), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n908), .B(new_n977), .C1(new_n992), .C2(new_n950), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n976), .A2(new_n987), .A3(new_n908), .A4(new_n977), .ZN(new_n995));
  AND4_X1   g570(.A1(KEYINPUT109), .A2(new_n994), .A3(KEYINPUT44), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n990), .B1(new_n993), .B2(KEYINPUT43), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT109), .B1(new_n997), .B2(new_n995), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n991), .B1(new_n996), .B2(new_n998), .ZN(G397));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(new_n887), .B2(G1384), .ZN(new_n1001));
  INV_X1    g576(.A(G125), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n466), .B2(new_n467), .ZN(new_n1003));
  OAI21_X1  g578(.A(G2105), .B1(new_n1003), .B2(new_n461), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1004), .A2(G40), .A3(new_n472), .A4(new_n469), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT110), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n844), .B(new_n847), .ZN(new_n1008));
  INV_X1    g583(.A(G1996), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n821), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1006), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(G1996), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n821), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n738), .B(new_n741), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n1007), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n606), .B(new_n731), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1018), .B1(new_n1006), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n1021));
  INV_X1    g596(.A(G1966), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1000), .A2(G1384), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT116), .B1(G164), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n500), .A2(new_n502), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n485), .A2(new_n488), .A3(new_n483), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT67), .B1(new_n493), .B2(new_n497), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n1030), .A3(new_n1023), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1005), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n886), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1026), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(KEYINPUT111), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n887), .B2(G1384), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT45), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1022), .B1(new_n1034), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1005), .A2(G2084), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1021), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1005), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT111), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n887), .A2(new_n1039), .A3(G1384), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1000), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1966), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1047), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1053), .A2(new_n1054), .A3(KEYINPUT118), .ZN(new_n1055));
  OAI21_X1  g630(.A(G168), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n1057));
  NAND2_X1  g632(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1042), .A2(new_n1021), .A3(new_n1047), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT118), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1062));
  AOI21_X1  g637(.A(G286), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT119), .B1(new_n1063), .B2(new_n1058), .ZN(new_n1064));
  OAI21_X1  g639(.A(G8), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1065), .A2(KEYINPUT120), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(KEYINPUT120), .ZN(new_n1067));
  INV_X1    g642(.A(G8), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G168), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(KEYINPUT51), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1066), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1060), .A2(new_n1064), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1061), .A2(new_n1062), .A3(new_n1069), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1044), .A2(new_n1045), .A3(new_n1033), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT121), .B(G1961), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G2078), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1049), .A2(new_n1052), .A3(KEYINPUT53), .A4(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1005), .B1(new_n1036), .B2(new_n1023), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1000), .B1(G164), .B2(G1384), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n1081), .A3(new_n1078), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1082), .A2(KEYINPUT122), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT122), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1077), .B(new_n1079), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G171), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1082), .A2(KEYINPUT122), .A3(new_n1083), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1080), .A2(KEYINPUT53), .A3(new_n1078), .A4(new_n1001), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1092), .A2(G301), .A3(new_n1077), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1087), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT123), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1095), .A2(new_n1099), .A3(new_n1096), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT55), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(G166), .B2(new_n1068), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n756), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1075), .B2(G2090), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1108), .A3(G8), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT50), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1110));
  NOR2_X1   g685(.A1(G164), .A2(G1384), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1005), .B1(new_n1111), .B2(new_n1043), .ZN(new_n1112));
  INV_X1    g687(.A(G2090), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1068), .B1(new_n1114), .B2(new_n1107), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1109), .B1(new_n1105), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1077), .B(new_n1093), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1096), .B1(new_n1117), .B2(G171), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1092), .A2(G301), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1038), .A2(new_n1040), .A3(new_n1033), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G8), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G1981), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n522), .A2(G86), .B1(G48), .B2(new_n526), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n585), .A2(G651), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1981), .B1(new_n526), .B2(G48), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n591), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1122), .B1(new_n1128), .B2(KEYINPUT49), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n588), .A2(new_n590), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1126), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(KEYINPUT49), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT113), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1128), .A2(KEYINPUT113), .A3(KEYINPUT49), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1129), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT112), .B(G1976), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT52), .B1(G288), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(G1976), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G288), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1122), .A2(new_n1139), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT52), .B1(new_n1121), .B2(new_n1141), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT115), .B1(new_n1137), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT49), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1121), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AND4_X1   g724(.A1(KEYINPUT113), .A2(new_n1131), .A3(KEYINPUT49), .A4(new_n1132), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT113), .B1(new_n1128), .B2(KEYINPUT49), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT115), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI221_X4 g730(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .C1(new_n1146), .C2(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT58), .B(G1341), .Z(new_n1157));
  NAND2_X1  g732(.A1(new_n1120), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(G1996), .B2(new_n1106), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n557), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT59), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1120), .A2(G2067), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1163), .B1(new_n800), .B2(new_n1075), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1164), .A2(KEYINPUT60), .A3(new_n921), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1159), .A2(KEYINPUT59), .A3(new_n557), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1162), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n921), .B1(new_n1164), .B2(KEYINPUT60), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(KEYINPUT60), .B2(new_n1164), .ZN(new_n1169));
  AOI21_X1  g744(.A(G1956), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1170));
  XNOR2_X1  g745(.A(KEYINPUT56), .B(G2072), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1080), .A2(new_n1081), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT57), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1174), .A2(KEYINPUT117), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(KEYINPUT117), .ZN(new_n1176));
  NAND3_X1  g751(.A1(G299), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n570), .A2(new_n574), .A3(KEYINPUT117), .A4(new_n1174), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1173), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1179), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1182), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1167), .B(new_n1169), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1183), .B1(new_n921), .B2(new_n1164), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1181), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1074), .A2(new_n1101), .A3(new_n1156), .A4(new_n1189), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n1065), .A2(G286), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1109), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1137), .A2(new_n1145), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1108), .A2(G8), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1194), .B(new_n1195), .C1(new_n1105), .C2(new_n1196), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1116), .B(new_n1191), .C1(new_n1146), .C2(new_n1155), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1197), .B1(new_n1198), .B2(KEYINPUT63), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1131), .B(KEYINPUT114), .Z(new_n1200));
  NAND2_X1  g775(.A1(new_n759), .A2(new_n1140), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1200), .B1(new_n1137), .B2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g777(.A1(new_n1202), .A2(new_n1122), .B1(new_n1195), .B2(new_n1192), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1190), .A2(new_n1199), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1116), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1205), .A2(G171), .A3(new_n1086), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1074), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1072), .A2(KEYINPUT62), .A3(new_n1073), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1206), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1020), .B1(new_n1204), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1008), .A2(new_n821), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1007), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1013), .ZN(new_n1214));
  AND2_X1   g789(.A1(new_n1214), .A2(KEYINPUT46), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1214), .A2(KEYINPUT46), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1213), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n1217), .B(KEYINPUT47), .Z(new_n1218));
  NOR2_X1   g793(.A1(G290), .A2(G1986), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1219), .ZN(new_n1220));
  XOR2_X1   g795(.A(KEYINPUT124), .B(KEYINPUT48), .Z(new_n1221));
  INV_X1    g796(.A(new_n1221), .ZN(new_n1222));
  NOR3_X1   g797(.A1(new_n1220), .A2(new_n1012), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1221), .B1(new_n1219), .B2(new_n1006), .ZN(new_n1224));
  NOR3_X1   g799(.A1(new_n1223), .A2(new_n1018), .A3(new_n1224), .ZN(new_n1225));
  OR2_X1    g800(.A1(new_n738), .A2(new_n741), .ZN(new_n1226));
  OAI22_X1  g801(.A1(new_n1015), .A2(new_n1226), .B1(G2067), .B2(new_n844), .ZN(new_n1227));
  AOI211_X1 g802(.A(new_n1218), .B(new_n1225), .C1(new_n1007), .C2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1211), .A2(new_n1228), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g804(.A1(new_n678), .A2(new_n681), .ZN(new_n1231));
  NOR2_X1   g805(.A1(G227), .A2(new_n459), .ZN(new_n1232));
  NAND3_X1  g806(.A1(new_n1231), .A2(KEYINPUT125), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n1233), .A2(new_n721), .ZN(new_n1234));
  INV_X1    g808(.A(new_n1232), .ZN(new_n1235));
  AOI21_X1  g809(.A(new_n1235), .B1(new_n678), .B2(new_n681), .ZN(new_n1236));
  NOR2_X1   g810(.A1(new_n1236), .A2(KEYINPUT125), .ZN(new_n1237));
  OAI21_X1  g811(.A(KEYINPUT126), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g812(.A(KEYINPUT125), .ZN(new_n1239));
  OAI21_X1  g813(.A(new_n1239), .B1(G401), .B2(new_n1235), .ZN(new_n1240));
  INV_X1    g814(.A(KEYINPUT126), .ZN(new_n1241));
  NAND4_X1  g815(.A1(new_n1240), .A2(new_n1241), .A3(new_n721), .A4(new_n1233), .ZN(new_n1242));
  AOI21_X1  g816(.A(new_n912), .B1(new_n1238), .B2(new_n1242), .ZN(new_n1243));
  AND2_X1   g817(.A1(new_n1243), .A2(new_n989), .ZN(G308));
  NAND2_X1  g818(.A1(new_n1243), .A2(new_n989), .ZN(G225));
endmodule


