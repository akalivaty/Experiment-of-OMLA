//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G141gat), .B(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n211), .B1(G155gat), .B2(G162gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT74), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G155gat), .B(G162gat), .Z(new_n214));
  OR2_X1    g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n214), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT29), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n217), .B(KEYINPUT76), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n208), .B2(KEYINPUT29), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(G228gat), .B2(G233gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G228gat), .A2(G233gat), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n215), .A2(new_n216), .ZN(new_n227));
  AOI211_X1 g026(.A(new_n226), .B(new_n221), .C1(new_n227), .C2(new_n223), .ZN(new_n228));
  OR3_X1    g027(.A1(new_n225), .A2(G22gat), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT79), .ZN(new_n230));
  OAI21_X1  g029(.A(G22gat), .B1(new_n225), .B2(new_n228), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G78gat), .B(G106gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT31), .B(G50gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT78), .ZN(new_n236));
  OAI211_X1 g035(.A(KEYINPUT79), .B(G22gat), .C1(new_n225), .C2(new_n228), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n229), .A2(new_n235), .A3(new_n231), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n243), .B(new_n244), .C1(G183gat), .C2(G190gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(KEYINPUT23), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n248), .B(KEYINPUT65), .ZN(new_n252));
  AOI22_X1  g051(.A1(KEYINPUT23), .A2(new_n252), .B1(new_n245), .B2(new_n246), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n245), .B(KEYINPUT64), .Z(new_n255));
  AOI211_X1 g054(.A(KEYINPUT25), .B(new_n250), .C1(KEYINPUT23), .C2(new_n248), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n254), .A2(KEYINPUT25), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT27), .B(G183gat), .ZN(new_n258));
  INV_X1    g057(.A(G190gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT26), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n252), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n252), .A2(new_n266), .A3(new_n263), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n249), .B1(new_n248), .B2(new_n263), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n241), .B(new_n262), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n257), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT72), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n273), .A3(new_n270), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n220), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n276), .B1(new_n257), .B2(new_n270), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT73), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n279), .A3(new_n209), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n271), .A2(new_n220), .A3(new_n276), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n272), .A2(new_n274), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n208), .B(new_n281), .C1(new_n282), .C2(new_n276), .ZN(new_n283));
  XNOR2_X1  g082(.A(G8gat), .B(G36gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(G64gat), .B(G92gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT30), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n280), .A2(new_n283), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n286), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G113gat), .B(G120gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(KEYINPUT1), .ZN(new_n298));
  XNOR2_X1  g097(.A(G127gat), .B(G134gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n222), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT4), .ZN(new_n302));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n300), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n217), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n227), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n217), .B2(new_n218), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n308), .A2(new_n300), .A3(new_n310), .A4(new_n219), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n302), .A2(new_n303), .A3(new_n307), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n227), .A2(new_n300), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n305), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(G225gat), .A3(G233gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(KEYINPUT5), .A3(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n305), .A2(new_n306), .ZN(new_n317));
  INV_X1    g116(.A(new_n301), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n311), .A2(KEYINPUT4), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n303), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G57gat), .B(G85gat), .Z(new_n324));
  XNOR2_X1  g123(.A(G1gat), .B(G29gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT6), .ZN(new_n330));
  INV_X1    g129(.A(new_n328), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n322), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n323), .A2(KEYINPUT6), .A3(new_n328), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n240), .B1(new_n296), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT36), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT70), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT69), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n271), .B2(new_n300), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n271), .A2(new_n300), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n257), .A2(new_n270), .A3(KEYINPUT69), .A4(new_n304), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT32), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n346), .B1(new_n343), .B2(new_n344), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G15gat), .B(G43gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(G71gat), .B(G99gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n343), .A2(new_n344), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT33), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n345), .A2(new_n347), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n349), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n358), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n356), .B1(new_n360), .B2(new_n348), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n359), .B2(new_n361), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n337), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n359), .A2(new_n361), .ZN(new_n367));
  INV_X1    g166(.A(new_n362), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(KEYINPUT36), .A3(new_n363), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n336), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n335), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT38), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT37), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n209), .B1(new_n277), .B2(new_n279), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n281), .B1(new_n282), .B2(new_n276), .ZN(new_n376));
  AOI211_X1 g175(.A(new_n374), .B(new_n375), .C1(new_n209), .C2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT37), .B1(new_n280), .B2(new_n283), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n373), .B(new_n286), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n378), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n280), .A2(new_n283), .A3(KEYINPUT37), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n373), .B1(new_n382), .B2(new_n286), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n372), .B(new_n379), .C1(KEYINPUT83), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n381), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n286), .B1(new_n385), .B2(new_n378), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT38), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n288), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n240), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n320), .A2(new_n303), .ZN(new_n391));
  NAND2_X1  g190(.A1(KEYINPUT80), .A2(KEYINPUT39), .ZN(new_n392));
  OR2_X1    g191(.A1(KEYINPUT80), .A2(KEYINPUT39), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n313), .A2(new_n303), .A3(new_n305), .ZN(new_n395));
  OAI211_X1 g194(.A(KEYINPUT39), .B(new_n395), .C1(new_n320), .C2(new_n303), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n331), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT40), .B1(new_n397), .B2(KEYINPUT81), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(KEYINPUT81), .A3(KEYINPUT40), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n401), .A2(KEYINPUT82), .A3(new_n329), .A4(new_n295), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n397), .A2(KEYINPUT81), .A3(KEYINPUT40), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n404), .A2(new_n398), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n295), .A2(new_n329), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n371), .B1(new_n390), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT35), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT84), .ZN(new_n411));
  AND4_X1   g210(.A1(new_n240), .A2(new_n369), .A3(new_n296), .A4(new_n363), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(new_n335), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n410), .A2(KEYINPUT84), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n412), .A2(new_n335), .A3(new_n411), .A4(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n409), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n418));
  INV_X1    g217(.A(G29gat), .ZN(new_n419));
  INV_X1    g218(.A(G36gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n421), .A2(new_n422), .B1(G29gat), .B2(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G43gat), .B(G50gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT15), .ZN(new_n426));
  OR3_X1    g225(.A1(new_n423), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n426), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(KEYINPUT15), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n423), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G15gat), .B(G22gat), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n434), .A2(G1gat), .ZN(new_n435));
  INV_X1    g234(.A(G8gat), .ZN(new_n436));
  INV_X1    g235(.A(G1gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT16), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n436), .B1(new_n435), .B2(new_n439), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT17), .A3(new_n430), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n433), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  OR2_X1    g243(.A1(new_n440), .A2(new_n441), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n431), .ZN(new_n446));
  NAND2_X1  g245(.A1(G229gat), .A2(G233gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT85), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT18), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n442), .B(new_n431), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT86), .B(KEYINPUT13), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(new_n447), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT18), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n448), .A2(KEYINPUT85), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(G113gat), .B(G141gat), .Z(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(G197gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT11), .B(G169gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(KEYINPUT12), .Z(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n463), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n450), .A2(new_n465), .A3(new_n455), .A4(new_n457), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT87), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n466), .A2(KEYINPUT87), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g269(.A1(G71gat), .A2(G78gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(G71gat), .A2(G78gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G57gat), .B(G64gat), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(G57gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(G64gat), .ZN(new_n478));
  INV_X1    g277(.A(G64gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G57gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G71gat), .B(G78gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n475), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n445), .B1(KEYINPUT21), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(G231gat), .A2(G233gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G183gat), .B(G211gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n485), .A2(KEYINPUT21), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT20), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT89), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n492), .B(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n490), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n498));
  XNOR2_X1  g297(.A(G127gat), .B(G155gat), .ZN(new_n499));
  XOR2_X1   g298(.A(new_n498), .B(new_n499), .Z(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n497), .B(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT41), .ZN(new_n503));
  INV_X1    g302(.A(G232gat), .ZN(new_n504));
  INV_X1    g303(.A(G233gat), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT8), .ZN(new_n508));
  NAND2_X1  g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G85gat), .ZN(new_n512));
  INV_X1    g311(.A(G92gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n508), .A2(new_n511), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n507), .ZN(new_n520));
  INV_X1    g319(.A(new_n507), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT92), .B1(new_n521), .B2(new_n517), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n521), .A2(new_n517), .ZN(new_n527));
  AOI22_X1  g326(.A1(KEYINPUT8), .A2(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .A4(new_n519), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n506), .B1(new_n431), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n532));
  XOR2_X1   g331(.A(G190gat), .B(G218gat), .Z(new_n533));
  NAND2_X1  g332(.A1(new_n433), .A2(new_n443), .ZN(new_n534));
  OAI221_X1 g333(.A(new_n531), .B1(new_n532), .B2(new_n533), .C1(new_n534), .C2(new_n530), .ZN(new_n535));
  XOR2_X1   g334(.A(G134gat), .B(G162gat), .Z(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n532), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n537), .B(new_n540), .Z(new_n541));
  NAND2_X1  g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT95), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n516), .A2(KEYINPUT94), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n527), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n518), .A2(new_n507), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n516), .A2(KEYINPUT94), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n485), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n476), .A2(new_n484), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT10), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n530), .A2(new_n485), .A3(KEYINPUT10), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n544), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT97), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n523), .A2(new_n529), .B1(new_n476), .B2(new_n484), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n516), .A2(KEYINPUT94), .A3(new_n547), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n547), .B1(new_n516), .B2(KEYINPUT94), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n558), .B1(new_n561), .B2(new_n485), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n543), .ZN(new_n563));
  OAI211_X1 g362(.A(KEYINPUT97), .B(new_n544), .C1(new_n552), .C2(new_n554), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G120gat), .B(G148gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G176gat), .B(G204gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT98), .ZN(new_n570));
  INV_X1    g369(.A(new_n568), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n571), .A3(new_n563), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT96), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n502), .A2(new_n541), .A3(new_n574), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n417), .A2(new_n470), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n372), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n295), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT16), .B(G8gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n581), .A2(KEYINPUT42), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(G8gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(KEYINPUT42), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G1325gat));
  NAND2_X1  g384(.A1(new_n369), .A2(new_n363), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(G15gat), .B1(new_n576), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n366), .A2(new_n370), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(G15gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT99), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n588), .B1(new_n576), .B2(new_n592), .ZN(G1326gat));
  INV_X1    g392(.A(new_n240), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT43), .B(G22gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(G1327gat));
  INV_X1    g398(.A(new_n541), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n289), .B1(new_n383), .B2(KEYINPUT83), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n335), .B1(new_n387), .B2(new_n388), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n602), .A3(new_n379), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n603), .A2(new_n240), .A3(new_n407), .A4(new_n402), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n413), .B1(new_n604), .B2(new_n371), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n600), .B1(new_n605), .B2(new_n416), .ZN(new_n606));
  INV_X1    g405(.A(new_n574), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n606), .A2(new_n470), .A3(new_n502), .A4(new_n607), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n608), .A2(G29gat), .A3(new_n335), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT45), .Z(new_n610));
  INV_X1    g409(.A(KEYINPUT44), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n417), .A2(new_n611), .A3(new_n541), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n417), .B2(new_n541), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n502), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n470), .A2(KEYINPUT102), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n617), .B(new_n464), .C1(new_n468), .C2(new_n469), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n615), .A2(new_n574), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(G29gat), .B1(new_n622), .B2(new_n335), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n610), .A2(new_n623), .ZN(G1328gat));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n622), .B2(new_n296), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n614), .A2(KEYINPUT103), .A3(new_n295), .A4(new_n621), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(G36gat), .A3(new_n627), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n608), .A2(G36gat), .A3(new_n296), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT46), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(G1329gat));
  INV_X1    g430(.A(G43gat), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n632), .B1(new_n608), .B2(new_n586), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n614), .A2(G43gat), .A3(new_n621), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n589), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT47), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT47), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n637), .B(new_n633), .C1(new_n634), .C2(new_n589), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(G1330gat));
  OAI211_X1 g438(.A(new_n594), .B(new_n621), .C1(new_n612), .C2(new_n613), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(G50gat), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT48), .B1(new_n641), .B2(KEYINPUT104), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n608), .A2(G50gat), .A3(new_n240), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n643), .B(new_n641), .C1(KEYINPUT104), .C2(KEYINPUT48), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(G1331gat));
  NOR2_X1   g446(.A1(new_n502), .A2(new_n541), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n335), .A2(new_n607), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n417), .A2(new_n648), .A3(new_n620), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G57gat), .ZN(G1332gat));
  NAND4_X1  g450(.A1(new_n417), .A2(new_n648), .A3(new_n574), .A4(new_n620), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n296), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT49), .B(G64gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n655), .B1(new_n653), .B2(new_n656), .ZN(G1333gat));
  INV_X1    g456(.A(G71gat), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n652), .B2(new_n586), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n652), .A2(new_n658), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(new_n590), .ZN(new_n662));
  NOR4_X1   g461(.A1(new_n652), .A2(KEYINPUT105), .A3(new_n658), .A4(new_n589), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n659), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g464(.A1(new_n652), .A2(new_n240), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(G78gat), .Z(G1335gat));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n615), .A2(new_n619), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT51), .B1(new_n606), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n417), .A2(new_n541), .A3(new_n669), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT51), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n668), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n606), .A2(KEYINPUT51), .A3(new_n669), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT106), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n674), .A2(new_n512), .A3(new_n649), .A4(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n574), .B(new_n669), .C1(new_n612), .C2(new_n613), .ZN(new_n679));
  OAI21_X1  g478(.A(G85gat), .B1(new_n679), .B2(new_n335), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(G1336gat));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n607), .B1(new_n675), .B2(new_n676), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n296), .A2(G92gat), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(G92gat), .B1(new_n679), .B2(new_n296), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT52), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT52), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n685), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1337gat));
  NOR3_X1   g490(.A1(new_n586), .A2(G99gat), .A3(new_n607), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT108), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n674), .A2(new_n677), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G99gat), .B1(new_n679), .B2(new_n589), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n694), .A2(new_n695), .A3(KEYINPUT109), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1338gat));
  INV_X1    g499(.A(G106gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n683), .A2(new_n701), .A3(new_n594), .ZN(new_n702));
  OAI21_X1  g501(.A(G106gat), .B1(new_n679), .B2(new_n240), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT53), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT53), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(G1339gat));
  NOR4_X1   g507(.A1(new_n502), .A2(new_n541), .A3(new_n619), .A4(new_n574), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT54), .B1(new_n557), .B2(new_n564), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n543), .B(new_n553), .C1(new_n562), .C2(KEYINPUT10), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n555), .A2(new_n712), .A3(KEYINPUT54), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n711), .A2(new_n571), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n710), .B1(new_n714), .B2(KEYINPUT55), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT54), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n553), .B1(new_n562), .B2(KEYINPUT10), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT97), .B1(new_n717), .B2(new_n544), .ZN(new_n718));
  INV_X1    g517(.A(new_n564), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n555), .A2(new_n712), .A3(KEYINPUT54), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n568), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT55), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(KEYINPUT111), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n715), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n720), .A2(KEYINPUT55), .A3(new_n568), .A4(new_n721), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n573), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n727), .A2(new_n726), .A3(new_n573), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n725), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n727), .A2(new_n726), .A3(new_n573), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n728), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(KEYINPUT112), .A3(new_n725), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n451), .A2(new_n454), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n444), .A2(new_n446), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(new_n447), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n462), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n468), .B2(new_n469), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT113), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n744), .B(new_n741), .C1(new_n468), .C2(new_n469), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n737), .A2(new_n541), .A3(new_n743), .A4(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n607), .A2(new_n742), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n737), .B2(new_n619), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n748), .B2(new_n541), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n709), .B1(new_n749), .B2(new_n502), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n750), .A2(new_n335), .A3(new_n295), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n586), .A2(new_n594), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OR3_X1    g552(.A1(new_n753), .A2(G113gat), .A3(new_n620), .ZN(new_n754));
  INV_X1    g553(.A(new_n753), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n470), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(KEYINPUT114), .A3(G113gat), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT114), .B1(new_n756), .B2(G113gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n754), .B1(new_n758), .B2(new_n759), .ZN(G1340gat));
  NAND2_X1  g559(.A1(new_n755), .A2(new_n574), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g561(.A1(new_n753), .A2(new_n502), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(G127gat), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n763), .B(new_n765), .ZN(G1342gat));
  NOR2_X1   g565(.A1(new_n753), .A2(new_n600), .ZN(new_n767));
  INV_X1    g566(.A(G134gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n769), .A2(KEYINPUT56), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(KEYINPUT56), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n770), .B(new_n771), .C1(new_n768), .C2(new_n767), .ZN(G1343gat));
  INV_X1    g571(.A(KEYINPUT58), .ZN(new_n773));
  AND4_X1   g572(.A1(KEYINPUT112), .A2(new_n725), .A3(new_n729), .A4(new_n730), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT112), .B1(new_n735), .B2(new_n725), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n619), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n747), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n541), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n743), .A2(new_n541), .A3(new_n745), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n733), .B2(new_n736), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n502), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n709), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n240), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT116), .B1(new_n783), .B2(KEYINPUT57), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n785), .B(new_n786), .C1(new_n750), .C2(new_n240), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n722), .A2(KEYINPUT117), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n722), .A2(KEYINPUT117), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n723), .A3(new_n789), .ZN(new_n790));
  AND4_X1   g589(.A1(new_n470), .A2(new_n790), .A3(new_n573), .A4(new_n727), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n600), .B1(new_n791), .B2(new_n747), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n615), .B1(new_n746), .B2(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(KEYINPUT57), .B(new_n594), .C1(new_n793), .C2(new_n709), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n784), .A2(new_n787), .A3(new_n794), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n590), .A2(new_n335), .A3(new_n295), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n619), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G141gat), .ZN(new_n798));
  INV_X1    g597(.A(G141gat), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n590), .A2(new_n240), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n751), .A2(new_n799), .A3(new_n470), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n773), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n773), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n795), .A2(new_n470), .A3(new_n796), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(G141gat), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT118), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(G141gat), .ZN(new_n807));
  INV_X1    g606(.A(new_n803), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810));
  INV_X1    g609(.A(new_n801), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n797), .B2(G141gat), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n809), .B(new_n810), .C1(new_n773), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n806), .A2(new_n813), .ZN(G1344gat));
  INV_X1    g613(.A(new_n800), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n607), .ZN(new_n816));
  INV_X1    g615(.A(G148gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n751), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n795), .A2(new_n796), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AOI211_X1 g619(.A(KEYINPUT59), .B(new_n817), .C1(new_n820), .C2(new_n574), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n783), .A2(KEYINPUT57), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n792), .B1(new_n731), .B2(new_n779), .ZN(new_n826));
  INV_X1    g625(.A(new_n470), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n826), .A2(new_n502), .B1(new_n575), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n786), .B1(new_n828), .B2(new_n240), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n783), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n825), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n574), .A3(new_n796), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n822), .B1(new_n832), .B2(G148gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n818), .B1(new_n821), .B2(new_n833), .ZN(G1345gat));
  NAND2_X1  g633(.A1(new_n751), .A2(new_n800), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(G155gat), .B1(new_n836), .B2(new_n615), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n615), .A2(G155gat), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n820), .B2(new_n838), .ZN(G1346gat));
  AOI21_X1  g638(.A(G162gat), .B1(new_n836), .B2(new_n541), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n541), .A2(G162gat), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n820), .B2(new_n841), .ZN(G1347gat));
  NAND2_X1  g641(.A1(new_n781), .A2(new_n782), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n372), .A2(new_n296), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n752), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G169gat), .B1(new_n845), .B2(new_n827), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT121), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n845), .B(KEYINPUT120), .ZN(new_n848));
  INV_X1    g647(.A(G169gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(new_n619), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(G1348gat));
  INV_X1    g650(.A(new_n845), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n852), .A2(G176gat), .A3(new_n574), .ZN(new_n853));
  AOI21_X1  g652(.A(G176gat), .B1(new_n848), .B2(new_n574), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(G1349gat));
  NAND3_X1  g657(.A1(new_n852), .A2(new_n258), .A3(new_n615), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n860));
  OAI21_X1  g659(.A(G183gat), .B1(new_n845), .B2(new_n502), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT125), .Z(new_n863));
  AND3_X1   g662(.A1(new_n859), .A2(KEYINPUT123), .A3(new_n861), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT123), .B1(new_n859), .B2(new_n861), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT124), .B1(new_n866), .B2(KEYINPUT60), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n868));
  NOR4_X1   g667(.A1(new_n864), .A2(new_n865), .A3(new_n868), .A4(new_n860), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n863), .B1(new_n867), .B2(new_n869), .ZN(G1350gat));
  OAI21_X1  g669(.A(G190gat), .B1(new_n845), .B2(new_n600), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT61), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n848), .A2(new_n259), .A3(new_n541), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1351gat));
  XOR2_X1   g673(.A(KEYINPUT126), .B(G197gat), .Z(new_n875));
  NAND2_X1  g674(.A1(new_n589), .A2(new_n844), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n831), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n878), .B2(new_n827), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n843), .A2(new_n800), .A3(new_n844), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n620), .A2(new_n875), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(G1352gat));
  XNOR2_X1  g681(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n883));
  INV_X1    g682(.A(new_n816), .ZN(new_n884));
  INV_X1    g683(.A(G204gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n843), .A2(new_n885), .A3(new_n844), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OR3_X1    g686(.A1(new_n884), .A2(new_n883), .A3(new_n886), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n831), .A2(new_n574), .A3(new_n877), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n887), .B(new_n888), .C1(new_n889), .C2(new_n885), .ZN(G1353gat));
  INV_X1    g689(.A(new_n880), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n203), .A3(new_n615), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n831), .A2(new_n615), .A3(new_n877), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n893), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT63), .B1(new_n893), .B2(G211gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(G1354gat));
  OAI21_X1  g695(.A(G218gat), .B1(new_n878), .B2(new_n600), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n891), .A2(new_n204), .A3(new_n541), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1355gat));
endmodule


