//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G71gat), .ZN(new_n204));
  INV_X1    g003(.A(G78gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G71gat), .A2(G78gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT9), .ZN(new_n209));
  XNOR2_X1  g008(.A(G57gat), .B(G64gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT91), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT93), .ZN(new_n213));
  INV_X1    g012(.A(G64gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT92), .ZN(new_n215));
  INV_X1    g014(.A(G57gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT92), .A2(G57gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n216), .A2(G64gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n213), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n218), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT92), .A2(G57gat), .ZN(new_n223));
  OAI21_X1  g022(.A(G64gat), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n220), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(KEYINPUT93), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n206), .B1(KEYINPUT9), .B2(new_n207), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT94), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT94), .ZN(new_n231));
  AOI211_X1 g030(.A(new_n231), .B(new_n228), .C1(new_n221), .C2(new_n226), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n212), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234));
  INV_X1    g033(.A(G85gat), .ZN(new_n235));
  INV_X1    g034(.A(G92gat), .ZN(new_n236));
  AOI22_X1  g035(.A1(KEYINPUT8), .A2(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT7), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(new_n235), .B2(new_n236), .ZN(new_n239));
  NAND3_X1  g038(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G99gat), .B(G106gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n233), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT10), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n212), .B(new_n243), .C1(new_n230), .C2(new_n232), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT10), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n203), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n202), .B1(new_n245), .B2(new_n247), .ZN(new_n252));
  XOR2_X1   g051(.A(G176gat), .B(G204gat), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT98), .ZN(new_n254));
  XNOR2_X1  g053(.A(G120gat), .B(G148gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OR3_X1    g056(.A1(new_n251), .A2(new_n252), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n251), .B2(new_n252), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT27), .B(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n271), .A2(new_n274), .B1(G183gat), .B2(G190gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n277), .A2(KEYINPUT26), .ZN(new_n278));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(KEYINPUT26), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n275), .B(new_n281), .C1(new_n274), .C2(new_n271), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT64), .B(G176gat), .Z(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(KEYINPUT23), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n279), .A2(KEYINPUT23), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n277), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(new_n273), .ZN(new_n291));
  NAND3_X1  g090(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n273), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n285), .A2(new_n286), .A3(new_n288), .A4(new_n294), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n292), .A2(KEYINPUT65), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(KEYINPUT65), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n296), .A2(new_n297), .A3(new_n293), .A4(new_n291), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n298), .A2(new_n288), .A3(new_n299), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n282), .B(new_n295), .C1(new_n300), .C2(new_n286), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G226gat), .A2(G233gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(G226gat), .A3(G233gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(KEYINPUT72), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n268), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n307), .A2(new_n267), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G8gat), .B(G36gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT30), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT73), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n322), .A3(new_n319), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n313), .A2(KEYINPUT30), .A3(new_n317), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n316), .B1(new_n311), .B2(new_n312), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(G113gat), .B(G120gat), .Z(new_n330));
  AOI21_X1  g129(.A(KEYINPUT1), .B1(new_n330), .B2(KEYINPUT69), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(KEYINPUT69), .B2(new_n330), .ZN(new_n332));
  XNOR2_X1  g131(.A(G127gat), .B(G134gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n333), .B(KEYINPUT68), .Z(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G113gat), .B(G120gat), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n336), .A2(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(KEYINPUT70), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .A4(new_n333), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G148gat), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n342), .A2(G141gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(G141gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n343), .A2(new_n344), .B1(new_n345), .B2(KEYINPUT2), .ZN(new_n346));
  NAND2_X1  g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT74), .ZN(new_n348));
  INV_X1    g147(.A(G155gat), .ZN(new_n349));
  INV_X1    g148(.A(G162gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n347), .A2(KEYINPUT74), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n346), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n347), .B1(new_n351), .B2(KEYINPUT2), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n343), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n354), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n359), .ZN(new_n360));
  OR2_X1    g159(.A1(new_n360), .A2(KEYINPUT4), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(KEYINPUT4), .ZN(new_n362));
  INV_X1    g161(.A(new_n359), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT3), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n341), .B1(new_n365), .B2(new_n359), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n361), .A2(new_n362), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n370));
  OAI21_X1  g169(.A(KEYINPUT78), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n372));
  INV_X1    g171(.A(new_n370), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n367), .A2(new_n372), .A3(new_n368), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n341), .A2(new_n359), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n360), .ZN(new_n377));
  INV_X1    g176(.A(new_n368), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n369), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(G57gat), .B(G85gat), .Z(new_n382));
  XNOR2_X1  g181(.A(G1gat), .B(G29gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  OR3_X1    g187(.A1(new_n367), .A2(KEYINPUT39), .A3(new_n368), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n376), .A2(new_n368), .A3(new_n360), .ZN(new_n390));
  OAI211_X1 g189(.A(KEYINPUT39), .B(new_n390), .C1(new_n367), .C2(new_n368), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT40), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n387), .B1(KEYINPUT81), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n392), .A2(KEYINPUT81), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n329), .A2(new_n388), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n359), .B2(new_n365), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n268), .B1(new_n398), .B2(KEYINPUT80), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(KEYINPUT80), .B2(new_n398), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n365), .B1(new_n267), .B2(KEYINPUT29), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n363), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n402), .B(new_n406), .C1(new_n268), .C2(new_n398), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(KEYINPUT31), .B(G50gat), .Z(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT79), .ZN(new_n410));
  XOR2_X1   g209(.A(G78gat), .B(G106gat), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(G22gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n410), .B(new_n412), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n408), .A2(new_n413), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n371), .A2(new_n374), .B1(new_n369), .B2(new_n379), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(new_n386), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n375), .A2(new_n386), .A3(new_n380), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT82), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n386), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n388), .A2(new_n422), .A3(new_n417), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n381), .A2(KEYINPUT6), .A3(new_n387), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT37), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n313), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n316), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(KEYINPUT38), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n309), .A2(new_n310), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n432), .B2(new_n268), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n309), .A2(new_n431), .A3(new_n268), .A4(new_n310), .ZN(new_n434));
  INV_X1    g233(.A(new_n307), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n434), .B1(new_n268), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT37), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n313), .A2(new_n427), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT38), .B1(new_n429), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n318), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n397), .B(new_n416), .C1(new_n426), .C2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n301), .B(new_n341), .ZN(new_n443));
  INV_X1    g242(.A(G227gat), .ZN(new_n444));
  INV_X1    g243(.A(G233gat), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT32), .ZN(new_n447));
  OR3_X1    g246(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT34), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT34), .B1(new_n446), .B2(new_n447), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G43gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(G71gat), .B(G99gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n452), .B(new_n453), .Z(new_n454));
  OAI211_X1 g253(.A(new_n451), .B(new_n454), .C1(new_n446), .C2(KEYINPUT33), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456));
  INV_X1    g255(.A(new_n454), .ZN(new_n457));
  OAI221_X1 g256(.A(new_n443), .B1(new_n456), .B2(new_n457), .C1(new_n444), .C2(new_n445), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n450), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n448), .A2(new_n449), .A3(new_n458), .A4(new_n455), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT36), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n425), .B1(new_n419), .B2(new_n420), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n327), .B1(new_n321), .B2(new_n323), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n416), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n462), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT35), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n426), .A2(new_n472), .A3(new_n465), .A4(new_n469), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n442), .A2(new_n468), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(G113gat), .B(G141gat), .Z(new_n475));
  XNOR2_X1  g274(.A(KEYINPUT84), .B(G197gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT11), .B(G169gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT12), .ZN(new_n480));
  INV_X1    g279(.A(G50gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G43gat), .ZN(new_n482));
  INV_X1    g281(.A(G43gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G50gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT15), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT86), .ZN(new_n487));
  NOR3_X1   g286(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n490), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT14), .ZN(new_n492));
  INV_X1    g291(.A(G29gat), .ZN(new_n493));
  INV_X1    g292(.A(G36gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(KEYINPUT86), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n489), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n496), .ZN(new_n499));
  OAI22_X1  g298(.A1(new_n499), .A2(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n484), .A3(KEYINPUT15), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT85), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n495), .A2(new_n496), .B1(G29gat), .B2(G36gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n504), .A2(new_n505), .A3(new_n501), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n498), .B(KEYINPUT17), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G8gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(G1gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G1gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT16), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n508), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n514), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n516), .A2(new_n510), .A3(G8gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n489), .A2(new_n491), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT85), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n505), .B1(new_n504), .B2(new_n501), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n519), .A2(new_n497), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n523));
  OAI211_X1 g322(.A(new_n507), .B(new_n518), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n515), .A2(new_n517), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n498), .B1(new_n503), .B2(new_n506), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n524), .A2(KEYINPUT18), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(KEYINPUT13), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n525), .A2(new_n526), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n522), .A2(new_n518), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n480), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n524), .A2(new_n528), .A3(new_n527), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(KEYINPUT89), .A3(new_n537), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n536), .A2(KEYINPUT88), .A3(new_n537), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT88), .B1(new_n536), .B2(new_n537), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n534), .ZN(new_n545));
  NOR3_X1   g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n542), .B1(new_n546), .B2(new_n480), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT90), .B1(new_n474), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n426), .A2(new_n441), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n396), .A2(new_n388), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n416), .B1(new_n465), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n468), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n473), .A2(new_n471), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT90), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(new_n547), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n260), .B1(new_n549), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n244), .B(new_n507), .C1(new_n522), .C2(new_n523), .ZN(new_n559));
  AND2_X1   g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n526), .A2(new_n243), .B1(KEYINPUT41), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n561), .A2(KEYINPUT96), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(KEYINPUT96), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n560), .A2(KEYINPUT41), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI221_X1 g365(.A(new_n559), .B1(KEYINPUT41), .B2(new_n560), .C1(new_n562), .C2(new_n563), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT97), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT97), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G190gat), .B(G218gat), .Z(new_n572));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n569), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n574), .B1(new_n569), .B2(new_n571), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(KEYINPUT21), .B(new_n212), .C1(new_n230), .C2(new_n232), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n518), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT20), .Z(new_n585));
  NOR2_X1   g384(.A1(new_n579), .A2(new_n581), .ZN(new_n586));
  OR3_X1    g385(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n583), .B2(new_n586), .ZN(new_n588));
  INV_X1    g387(.A(new_n233), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(new_n290), .ZN(new_n591));
  INV_X1    g390(.A(G211gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n589), .A2(KEYINPUT21), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT21), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n595), .B1(new_n233), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n587), .A2(new_n588), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n587), .B2(new_n588), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n577), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n558), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(new_n464), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(new_n512), .ZN(G1324gat));
  NAND3_X1  g405(.A1(new_n558), .A2(new_n603), .A3(new_n329), .ZN(new_n607));
  XOR2_X1   g406(.A(KEYINPUT16), .B(G8gat), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n607), .A2(KEYINPUT42), .A3(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n607), .A2(new_n609), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT42), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n612), .B1(new_n607), .B2(G8gat), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n610), .B1(new_n611), .B2(new_n613), .ZN(G1325gat));
  INV_X1    g413(.A(new_n604), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n615), .A2(G15gat), .A3(new_n463), .ZN(new_n616));
  INV_X1    g415(.A(new_n462), .ZN(new_n617));
  AOI21_X1  g416(.A(G15gat), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n616), .A2(new_n618), .ZN(G1326gat));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n416), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT43), .B(G22gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(G1327gat));
  INV_X1    g421(.A(KEYINPUT45), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n388), .A2(new_n417), .A3(new_n423), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n493), .A3(new_n425), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n558), .A2(new_n602), .A3(new_n577), .A4(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(KEYINPUT99), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n577), .A2(new_n602), .ZN(new_n630));
  AOI211_X1 g429(.A(new_n260), .B(new_n630), .C1(new_n549), .C2(new_n557), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n631), .B2(new_n626), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n623), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n555), .A2(KEYINPUT101), .A3(KEYINPUT44), .A4(new_n577), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n602), .ZN(new_n635));
  INV_X1    g434(.A(new_n577), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n553), .B2(new_n554), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT44), .B1(new_n637), .B2(KEYINPUT101), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n260), .B(KEYINPUT100), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(new_n548), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n635), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(G29gat), .B1(new_n644), .B2(new_n464), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n627), .A2(KEYINPUT99), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n631), .A2(new_n629), .A3(new_n626), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(KEYINPUT45), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n633), .A2(new_n645), .A3(new_n648), .ZN(G1328gat));
  NAND3_X1  g448(.A1(new_n631), .A2(new_n494), .A3(new_n329), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n650), .A2(KEYINPUT46), .ZN(new_n651));
  OAI21_X1  g450(.A(G36gat), .B1(new_n644), .B2(new_n465), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(KEYINPUT46), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(G1329gat));
  AOI21_X1  g453(.A(new_n483), .B1(new_n643), .B2(new_n463), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n462), .A2(G43gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n631), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(KEYINPUT47), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT47), .ZN(new_n660));
  INV_X1    g459(.A(new_n658), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(G1330gat));
  AOI21_X1  g462(.A(new_n481), .B1(new_n643), .B2(new_n467), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n416), .A2(G50gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n631), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(KEYINPUT48), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT48), .ZN(new_n669));
  INV_X1    g468(.A(new_n667), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n664), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(G1331gat));
  OAI211_X1 g471(.A(new_n601), .B(new_n548), .C1(new_n575), .C2(new_n576), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n474), .A2(new_n639), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n464), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n624), .A2(KEYINPUT102), .A3(new_n425), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n222), .A2(new_n223), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1332gat));
  AOI21_X1  g481(.A(new_n465), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT103), .ZN(new_n685));
  NOR2_X1   g484(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1333gat));
  AOI21_X1  g486(.A(G71gat), .B1(new_n674), .B2(new_n617), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT36), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n462), .B(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n204), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n688), .B1(new_n674), .B2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT104), .B(KEYINPUT50), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1334gat));
  NAND2_X1  g493(.A1(new_n674), .A2(new_n467), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G78gat), .ZN(G1335gat));
  INV_X1    g495(.A(KEYINPUT51), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n601), .A2(new_n547), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n637), .B2(KEYINPUT105), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n474), .A2(new_n700), .A3(new_n636), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n697), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n474), .B2(new_n636), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n637), .A2(KEYINPUT105), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT51), .A4(new_n698), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n260), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n464), .A2(G85gat), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n637), .A2(KEYINPUT101), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n707), .A2(new_n547), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n712), .A2(new_n602), .A3(new_n634), .A4(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G85gat), .B1(new_n714), .B2(new_n464), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n709), .A2(new_n715), .ZN(G1336gat));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  INV_X1    g516(.A(new_n713), .ZN(new_n718));
  NOR4_X1   g517(.A1(new_n635), .A2(new_n638), .A3(new_n465), .A4(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n719), .B2(new_n236), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n465), .A2(G92gat), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  AOI211_X1 g521(.A(new_n639), .B(new_n722), .C1(new_n702), .C2(new_n705), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT52), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n639), .B1(new_n702), .B2(new_n705), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n721), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727));
  OAI21_X1  g526(.A(G92gat), .B1(new_n714), .B2(new_n465), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n726), .A2(new_n717), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n724), .A2(new_n729), .ZN(G1337gat));
  NOR3_X1   g529(.A1(new_n462), .A2(new_n707), .A3(G99gat), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n706), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(G99gat), .B1(new_n714), .B2(new_n690), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1338gat));
  OAI21_X1  g533(.A(KEYINPUT107), .B1(new_n714), .B2(new_n416), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n635), .A2(new_n638), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n736), .A2(new_n737), .A3(new_n467), .A4(new_n713), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n735), .A2(new_n738), .A3(G106gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n416), .A2(G106gat), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT53), .B1(new_n725), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n740), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n639), .B(new_n743), .C1(new_n702), .C2(new_n705), .ZN(new_n744));
  INV_X1    g543(.A(G106gat), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n635), .A2(new_n638), .A3(new_n718), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n467), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT53), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n742), .A2(new_n748), .ZN(G1339gat));
  NAND2_X1  g548(.A1(new_n248), .A2(new_n250), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n202), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n248), .A2(new_n250), .A3(new_n203), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(KEYINPUT54), .A3(new_n752), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT108), .B(KEYINPUT54), .Z(new_n754));
  AOI21_X1  g553(.A(new_n256), .B1(new_n251), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(KEYINPUT55), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n258), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT109), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n756), .A2(new_n759), .A3(new_n258), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT55), .B1(new_n753), .B2(new_n755), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n758), .A2(new_n547), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n532), .A2(new_n533), .A3(new_n531), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n528), .B1(new_n524), .B2(new_n527), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n479), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n542), .A2(new_n767), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n260), .A2(KEYINPUT110), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT110), .B1(new_n260), .B2(new_n768), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n577), .B1(new_n763), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n761), .B1(new_n757), .B2(KEYINPUT109), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(new_n577), .A3(new_n768), .A4(new_n760), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n602), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n673), .A2(new_n260), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n470), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n678), .A2(new_n329), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT111), .Z(new_n782));
  NOR2_X1   g581(.A1(new_n548), .A2(G113gat), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT112), .Z(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n779), .A2(new_n425), .A3(new_n624), .A4(new_n465), .ZN(new_n786));
  OAI21_X1  g585(.A(G113gat), .B1(new_n786), .B2(new_n548), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1340gat));
  INV_X1    g587(.A(G120gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n782), .A2(new_n789), .A3(new_n260), .ZN(new_n790));
  OAI21_X1  g589(.A(G120gat), .B1(new_n786), .B2(new_n639), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1341gat));
  INV_X1    g591(.A(G127gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n786), .A2(new_n793), .A3(new_n602), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n601), .A3(new_n780), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n793), .B2(new_n795), .ZN(G1342gat));
  OR3_X1    g595(.A1(new_n781), .A2(G134gat), .A3(new_n636), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(KEYINPUT56), .ZN(new_n798));
  OAI21_X1  g597(.A(G134gat), .B1(new_n786), .B2(new_n636), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(KEYINPUT56), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(G1343gat));
  NOR3_X1   g600(.A1(new_n463), .A2(new_n329), .A3(new_n464), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n260), .A2(new_n768), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n547), .A2(new_n756), .A3(new_n258), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n248), .A2(new_n250), .A3(new_n203), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n806), .A2(new_n251), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n750), .A2(new_n202), .A3(new_n754), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n257), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT113), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n753), .A2(new_n813), .A3(new_n755), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n804), .B1(new_n805), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n774), .B1(new_n577), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n777), .B1(new_n817), .B2(new_n602), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n416), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n803), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n547), .A2(new_n756), .A3(new_n258), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n753), .A2(new_n755), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT55), .B1(new_n824), .B2(KEYINPUT113), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n823), .B1(new_n814), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n636), .B1(new_n826), .B2(new_n804), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n601), .B1(new_n827), .B2(new_n774), .ZN(new_n828));
  OAI211_X1 g627(.A(KEYINPUT114), .B(new_n820), .C1(new_n828), .C2(new_n777), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n822), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n776), .A2(new_n778), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT57), .B1(new_n831), .B2(new_n467), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n547), .B(new_n802), .C1(new_n830), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(G141gat), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n678), .A2(new_n329), .A3(new_n463), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n416), .B1(new_n776), .B2(new_n778), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n548), .A2(G141gat), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n834), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI211_X1 g640(.A(KEYINPUT116), .B(new_n838), .C1(new_n833), .C2(G141gat), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT58), .B(new_n841), .C1(new_n842), .C2(new_n840), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n834), .A2(new_n839), .ZN(new_n846));
  OAI211_X1 g645(.A(KEYINPUT115), .B(new_n845), .C1(new_n846), .C2(KEYINPUT116), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n844), .B1(new_n843), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(G1344gat));
  AND2_X1   g649(.A1(new_n835), .A2(new_n836), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n342), .A3(new_n260), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n773), .A2(new_n577), .A3(new_n760), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n768), .B1(new_n854), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n827), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n777), .B1(new_n858), .B2(new_n602), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n819), .B1(new_n859), .B2(new_n416), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n836), .A2(KEYINPUT57), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n802), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n862), .A2(new_n707), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n853), .B1(new_n864), .B2(G148gat), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n830), .A2(new_n832), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n863), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT59), .B(new_n342), .C1(new_n867), .C2(new_n260), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n852), .B1(new_n865), .B2(new_n868), .ZN(G1345gat));
  AOI21_X1  g668(.A(G155gat), .B1(new_n851), .B2(new_n601), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n602), .A2(new_n349), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n867), .B2(new_n871), .ZN(G1346gat));
  NAND3_X1  g671(.A1(new_n851), .A2(new_n350), .A3(new_n577), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT119), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n866), .A2(new_n636), .A3(new_n863), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n350), .B2(new_n875), .ZN(G1347gat));
  NOR2_X1   g675(.A1(new_n679), .A2(new_n465), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n779), .ZN(new_n878));
  OAI21_X1  g677(.A(G169gat), .B1(new_n878), .B2(new_n548), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n831), .A2(new_n464), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n470), .A2(new_n465), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT120), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n547), .A2(new_n284), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(G1348gat));
  OR3_X1    g685(.A1(new_n878), .A2(new_n283), .A3(new_n639), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(KEYINPUT121), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(KEYINPUT121), .ZN(new_n889));
  AOI21_X1  g688(.A(G176gat), .B1(new_n883), .B2(new_n260), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(G1349gat));
  NAND3_X1  g690(.A1(new_n883), .A2(new_n601), .A3(new_n272), .ZN(new_n892));
  OAI21_X1  g691(.A(G183gat), .B1(new_n878), .B2(new_n602), .ZN(new_n893));
  NAND2_X1  g692(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n895), .B(new_n896), .Z(G1350gat));
  OAI21_X1  g696(.A(G190gat), .B1(new_n878), .B2(new_n636), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT61), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n273), .A3(new_n577), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1351gat));
  NAND2_X1  g700(.A1(new_n877), .A2(new_n690), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n862), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G197gat), .B1(new_n904), .B2(new_n548), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n463), .A2(new_n465), .A3(new_n416), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT123), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(new_n880), .ZN(new_n908));
  INV_X1    g707(.A(G197gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n547), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n905), .A2(new_n910), .ZN(G1352gat));
  OAI21_X1  g710(.A(G204gat), .B1(new_n904), .B2(new_n639), .ZN(new_n912));
  INV_X1    g711(.A(G204gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n908), .A2(new_n913), .A3(new_n260), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915));
  OR3_X1    g714(.A1(new_n914), .A2(new_n915), .A3(KEYINPUT62), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(KEYINPUT62), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n915), .B1(new_n914), .B2(KEYINPUT62), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n912), .A2(new_n916), .A3(new_n917), .A4(new_n918), .ZN(G1353gat));
  NAND3_X1  g718(.A1(new_n908), .A2(new_n592), .A3(new_n601), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT125), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n592), .B1(new_n903), .B2(new_n601), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(KEYINPUT63), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(KEYINPUT63), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(G1354gat));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n908), .A2(new_n577), .ZN(new_n927));
  INV_X1    g726(.A(G218gat), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n903), .A2(G218gat), .A3(new_n577), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n926), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n929), .B(KEYINPUT126), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(KEYINPUT127), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1355gat));
endmodule


