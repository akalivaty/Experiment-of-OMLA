//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G219), .A3(G220), .A4(G218), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G137), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n461), .A2(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n460), .A2(new_n462), .B1(new_n463), .B2(G101), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(new_n461), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G160));
  NAND2_X1  g042(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n461), .B1(new_n468), .B2(new_n473), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  AND2_X1   g056(.A1(G126), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n460), .A2(new_n482), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(new_n469), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT68), .B(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n460), .A2(new_n494), .A3(KEYINPUT4), .A4(new_n489), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n487), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  NAND2_X1  g072(.A1(G75), .A2(G543), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G62), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT69), .B(G651), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT69), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI211_X1 g088(.A(G50), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n516), .B1(new_n512), .B2(new_n513), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n506), .B(new_n514), .C1(new_n515), .C2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NOR2_X1   g094(.A1(new_n510), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n508), .A2(KEYINPUT69), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT6), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n513), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n501), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n526), .B1(new_n522), .B2(new_n523), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n501), .A2(new_n508), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n529), .A2(G63), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n525), .A2(new_n528), .A3(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  AOI22_X1  g110(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n504), .ZN(new_n537));
  OAI211_X1 g112(.A(G52), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n538));
  OAI211_X1 g113(.A(G90), .B(new_n516), .C1(new_n512), .C2(new_n513), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n540), .B1(new_n538), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT71), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n545), .B(new_n537), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n524), .A2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n527), .A2(G43), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n504), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n523), .B1(new_n504), .B2(new_n507), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n560), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT72), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n566), .B2(new_n501), .ZN(new_n567));
  AOI22_X1  g142(.A1(G91), .A2(new_n524), .B1(new_n567), .B2(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(G299));
  AND2_X1   g144(.A1(new_n544), .A2(new_n546), .ZN(G301));
  NAND2_X1  g145(.A1(new_n524), .A2(G87), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n560), .A2(G49), .A3(G543), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n573), .B(G651), .C1(new_n516), .C2(G74), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT73), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n571), .A2(new_n572), .A3(new_n574), .A4(new_n576), .ZN(G288));
  OAI211_X1 g152(.A(G48), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n578));
  OAI211_X1 g153(.A(G86), .B(new_n516), .C1(new_n512), .C2(new_n513), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n516), .B2(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT74), .B1(new_n583), .B2(new_n504), .ZN(new_n584));
  OAI21_X1  g159(.A(G61), .B1(new_n499), .B2(new_n500), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(new_n581), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT74), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n586), .A2(new_n587), .A3(new_n505), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n580), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n524), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n527), .A2(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n592), .C1(new_n504), .C2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(new_n524), .A2(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n501), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n527), .A2(G54), .B1(G651), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g179(.A(new_n603), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G297));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G280));
  INV_X1    g184(.A(new_n602), .ZN(new_n610));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n460), .A2(new_n463), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT76), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT75), .ZN(new_n625));
  OR3_X1    g200(.A1(new_n625), .A2(new_n461), .A3(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n461), .B2(G111), .ZN(new_n627));
  AND3_X1   g202(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n623), .A2(new_n628), .B1(new_n476), .B2(G123), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n474), .A2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2096), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n620), .A2(new_n632), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT77), .B(KEYINPUT14), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT15), .B(G2435), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2438), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2430), .Z(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n637), .B2(new_n638), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n640), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(G401));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1961), .B(G1966), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT78), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  OR2_X1    g245(.A1(new_n663), .A2(new_n665), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n671), .A2(new_n668), .A3(new_n666), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n670), .B(new_n672), .C1(new_n668), .C2(new_n671), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT79), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT82), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT81), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT80), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  XOR2_X1   g255(.A(G1981), .B(G1986), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n674), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(new_n682), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(G229));
  NAND2_X1  g263(.A1(new_n610), .A2(G16), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G4), .B2(G16), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT88), .B(G1348), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G35), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G162), .B2(new_n693), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT29), .B(G2090), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(G16), .A2(G19), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n552), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT89), .B(G1341), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n693), .A2(G26), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT28), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n474), .A2(G140), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n476), .A2(G128), .ZN(new_n705));
  OR2_X1    g280(.A1(G104), .A2(G2105), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n706), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n703), .B1(new_n708), .B2(G29), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G2067), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n692), .A2(new_n697), .A3(new_n701), .A4(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G20), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT23), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n607), .B2(new_n712), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(G1956), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(G1956), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n690), .B2(new_n691), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n711), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(G303), .A2(G16), .ZN(new_n720));
  INV_X1    g295(.A(G22), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(G16), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(G1971), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G1971), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n725), .B(new_n722), .C1(G303), .C2(G16), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n712), .A2(G23), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G288), .B2(G16), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT33), .B(G1976), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n730), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n728), .B(new_n732), .C1(G288), .C2(G16), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n727), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT34), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n580), .A2(new_n589), .A3(G16), .ZN(new_n736));
  OR2_X1    g311(.A1(G6), .A2(G16), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT32), .B(G1981), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(KEYINPUT85), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT85), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n741), .A2(new_n745), .A3(new_n742), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n734), .A2(new_n735), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT35), .B(G1991), .Z(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G107), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n476), .B2(G119), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT83), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n474), .A2(G131), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n754), .B1(new_n753), .B2(new_n755), .ZN(new_n758));
  OAI21_X1  g333(.A(G29), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT84), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n693), .A2(G25), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n749), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n758), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n693), .B1(new_n766), .B2(new_n756), .ZN(new_n767));
  INV_X1    g342(.A(new_n761), .ZN(new_n768));
  OAI21_X1  g343(.A(KEYINPUT84), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n769), .A2(new_n748), .A3(new_n762), .ZN(new_n770));
  MUX2_X1   g345(.A(G24), .B(G290), .S(G16), .Z(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1986), .Z(new_n772));
  NAND4_X1  g347(.A1(new_n747), .A2(new_n765), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n734), .A2(new_n744), .A3(new_n746), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(KEYINPUT34), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT86), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n774), .A2(KEYINPUT86), .A3(KEYINPUT34), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n719), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  AND4_X1   g360(.A1(new_n747), .A2(new_n765), .A3(new_n770), .A4(new_n772), .ZN(new_n786));
  AOI21_X1  g361(.A(KEYINPUT86), .B1(new_n774), .B2(KEYINPUT34), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n774), .A2(KEYINPUT86), .A3(KEYINPUT34), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n786), .B(new_n781), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n693), .A2(G32), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n476), .A2(G129), .ZN(new_n793));
  NAND3_X1  g368(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT26), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n796), .A2(new_n797), .B1(G105), .B2(new_n463), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n474), .A2(G141), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n792), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT27), .B(G1996), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n693), .A2(G33), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n474), .A2(G139), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT25), .Z(new_n808));
  AOI22_X1  g383(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n806), .B(new_n808), .C1(new_n461), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n805), .B1(new_n810), .B2(G29), .ZN(new_n811));
  INV_X1    g386(.A(G2072), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n811), .A2(KEYINPUT90), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(KEYINPUT90), .B1(new_n811), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(G27), .A2(G29), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G164), .B2(G29), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(G2078), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT24), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(G34), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(G34), .ZN(new_n821));
  AOI21_X1  g396(.A(G29), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n466), .B2(G29), .ZN(new_n823));
  INV_X1    g398(.A(G2084), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G2078), .B2(new_n817), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n826), .B(new_n828), .C1(new_n812), .C2(new_n811), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n804), .A2(new_n815), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(G5), .A2(G16), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G171), .B2(G16), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT93), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G1961), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n712), .B1(new_n544), .B2(new_n546), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT93), .B1(new_n836), .B2(new_n831), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n830), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT94), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT91), .B1(new_n631), .B2(new_n693), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT91), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n629), .A2(new_n842), .A3(G29), .A4(new_n630), .ZN(new_n843));
  INV_X1    g418(.A(G28), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(KEYINPUT30), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(G29), .B1(new_n844), .B2(KEYINPUT30), .ZN(new_n847));
  NOR2_X1   g422(.A1(KEYINPUT31), .A2(G11), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(KEYINPUT31), .A2(G11), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n846), .A2(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n841), .A2(new_n843), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n712), .A2(G21), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G286), .B2(G16), .ZN(new_n854));
  INV_X1    g429(.A(G1966), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(KEYINPUT92), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT92), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n854), .B2(new_n855), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n852), .B(new_n856), .C1(new_n858), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n834), .A2(new_n837), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(G1961), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n839), .B1(new_n840), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n835), .B1(new_n834), .B2(new_n837), .ZN(new_n866));
  OAI21_X1  g441(.A(KEYINPUT94), .B1(new_n866), .B2(new_n861), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n862), .A2(G1961), .ZN(new_n869));
  INV_X1    g444(.A(new_n861), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n870), .A3(new_n840), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n830), .A2(new_n838), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n872), .A3(new_n867), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT95), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n791), .A2(KEYINPUT96), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT96), .B1(new_n791), .B2(new_n875), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(G311));
  NAND2_X1  g453(.A1(new_n791), .A2(new_n875), .ZN(G150));
  NAND2_X1  g454(.A1(new_n610), .A2(G559), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n527), .A2(G55), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n524), .A2(G93), .ZN(new_n883));
  NAND2_X1  g458(.A1(G80), .A2(G543), .ZN(new_n884));
  INV_X1    g459(.A(G67), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n501), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n886), .A2(KEYINPUT97), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n505), .B1(new_n886), .B2(KEYINPUT97), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n882), .B(new_n883), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n552), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n881), .B(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n891), .A2(KEYINPUT39), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(KEYINPUT39), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n892), .A2(new_n893), .A3(G860), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n889), .A2(G860), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT37), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n894), .A2(new_n896), .ZN(G145));
  XNOR2_X1  g472(.A(new_n801), .B(new_n496), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n753), .A2(new_n755), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n708), .B(KEYINPUT98), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n810), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n474), .A2(G142), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n476), .A2(G130), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n461), .A2(G118), .ZN(new_n906));
  OAI21_X1  g481(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n904), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n618), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n903), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n903), .A2(new_n910), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n901), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n913), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n900), .A3(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n631), .B(new_n466), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n480), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n919), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n914), .A2(new_n916), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g500(.A(G868), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n889), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(G290), .B(G166), .ZN(new_n928));
  XNOR2_X1  g503(.A(G305), .B(G288), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n928), .B(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n932), .B2(KEYINPUT42), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(KEYINPUT42), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n610), .A2(new_n607), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n602), .A2(G299), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(KEYINPUT41), .B2(new_n938), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n938), .B(KEYINPUT99), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n552), .B(new_n889), .Z(new_n944));
  XNOR2_X1  g519(.A(new_n613), .B(new_n944), .ZN(new_n945));
  MUX2_X1   g520(.A(new_n942), .B(new_n943), .S(new_n945), .Z(new_n946));
  XNOR2_X1  g521(.A(new_n935), .B(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n927), .B1(new_n947), .B2(new_n926), .ZN(G295));
  OAI21_X1  g523(.A(new_n927), .B1(new_n947), .B2(new_n926), .ZN(G331));
  AND3_X1   g524(.A1(new_n544), .A2(G168), .A3(new_n546), .ZN(new_n950));
  AOI21_X1  g525(.A(G168), .B1(new_n544), .B2(new_n546), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n950), .A2(new_n951), .A3(new_n890), .ZN(new_n952));
  NAND2_X1  g527(.A1(G171), .A2(G286), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n544), .A2(G168), .A3(new_n546), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n944), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n952), .A2(new_n955), .A3(new_n938), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n952), .B2(new_n955), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(new_n944), .A3(new_n954), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT102), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n956), .B1(new_n961), .B2(new_n942), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n962), .B2(new_n931), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n890), .B1(new_n950), .B2(new_n951), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT102), .B1(new_n964), .B2(new_n959), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n952), .A2(new_n957), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n942), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n956), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n930), .B(KEYINPUT103), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT43), .B1(new_n963), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n967), .A2(new_n931), .A3(new_n968), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n923), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n938), .A2(KEYINPUT41), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n964), .A2(new_n959), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n979), .B(new_n980), .C1(new_n977), .C2(new_n978), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n943), .A2(new_n958), .A3(new_n960), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n970), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n975), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT44), .B1(new_n973), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n984), .B1(new_n963), .B2(new_n972), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n975), .A2(new_n983), .A3(KEYINPUT43), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n986), .A2(new_n990), .ZN(G397));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT45), .B1(new_n496), .B2(new_n992), .ZN(new_n994));
  OAI211_X1 g569(.A(G40), .B(new_n464), .C1(new_n465), .C2(new_n461), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT114), .B1(new_n996), .B2(G1966), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n496), .A2(new_n998), .A3(new_n992), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n496), .B2(new_n992), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n999), .A2(new_n1000), .A3(new_n995), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n824), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n496), .A2(new_n992), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n995), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n855), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n997), .A2(G168), .A3(new_n1002), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n995), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1966), .B1(new_n1013), .B2(new_n1007), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1014), .A2(new_n1009), .B1(new_n1001), .B2(new_n824), .ZN(new_n1015));
  AOI21_X1  g590(.A(G168), .B1(new_n1015), .B2(new_n997), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT51), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT62), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1011), .A2(new_n1019), .A3(G8), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n583), .A2(KEYINPUT74), .A3(new_n504), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n587), .B1(new_n586), .B2(new_n505), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n578), .A2(new_n579), .ZN(new_n1025));
  OAI21_X1  g600(.A(G1981), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT111), .B(G1981), .Z(new_n1027));
  NAND3_X1  g602(.A1(new_n580), .A2(new_n589), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(KEYINPUT112), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n1030));
  NAND3_X1  g605(.A1(G305), .A2(new_n1030), .A3(G1981), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT49), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1006), .A2(new_n992), .A3(new_n496), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G8), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1029), .A2(new_n1037), .A3(new_n1031), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1007), .A2(KEYINPUT107), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT107), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n496), .A2(new_n1041), .A3(KEYINPUT45), .A4(new_n992), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1013), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT108), .B(G1971), .Z(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT109), .B(G2090), .Z(new_n1046));
  NAND2_X1  g621(.A1(new_n1001), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  NOR3_X1   g625(.A1(G166), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1048), .A2(new_n1054), .A3(G8), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(KEYINPUT110), .ZN(new_n1057));
  INV_X1    g632(.A(G1976), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1036), .B(new_n1057), .C1(new_n1058), .C2(G288), .ZN(new_n1059));
  NAND3_X1  g634(.A1(G288), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1060));
  NOR2_X1   g635(.A1(G288), .A2(new_n1058), .ZN(new_n1061));
  OAI22_X1  g636(.A1(new_n1035), .A2(new_n1061), .B1(KEYINPUT110), .B2(new_n1056), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1039), .A2(new_n1055), .A3(new_n1063), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1043), .A2(new_n1044), .B1(new_n1001), .B2(new_n1046), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1050), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1048), .A2(KEYINPUT113), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1053), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n1071));
  INV_X1    g646(.A(G2078), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1013), .A2(new_n1040), .A3(new_n1072), .A4(new_n1042), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1074), .A2(G2078), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1013), .A2(new_n1007), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n995), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n496), .A2(new_n998), .A3(new_n992), .ZN(new_n1084));
  AOI21_X1  g659(.A(G1961), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1079), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n835), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(KEYINPUT123), .A3(new_n1081), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(G301), .B1(new_n1078), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1064), .A2(new_n1070), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT126), .B1(new_n1021), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1039), .A2(new_n1055), .A3(new_n1063), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1054), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1094), .A2(new_n1095), .A3(new_n1098), .A4(new_n1091), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT62), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1093), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1028), .ZN(new_n1103));
  NOR2_X1   g678(.A1(G288), .A2(G1976), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1039), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1039), .A2(new_n1063), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1105), .A2(new_n1035), .B1(new_n1106), .B2(new_n1055), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1050), .B(G286), .C1(new_n1015), .C2(new_n997), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1098), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1053), .B1(new_n1065), .B2(new_n1050), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1064), .A2(new_n1112), .A3(KEYINPUT63), .A4(new_n1108), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1107), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G1956), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1087), .A2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1013), .A2(new_n1040), .A3(new_n1042), .A4(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n563), .A2(new_n568), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n563), .B2(new_n568), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1116), .B(new_n1118), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT117), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1119), .ZN(new_n1125));
  NAND2_X1  g700(.A1(G299), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n563), .A2(new_n568), .A3(new_n1119), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1130), .A2(KEYINPUT118), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT118), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G2067), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1006), .A2(new_n992), .A3(new_n1135), .A4(new_n496), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT116), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1348), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1087), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n610), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1123), .B1(new_n1134), .B2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1122), .A2(KEYINPUT61), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1131), .A2(new_n1128), .A3(new_n1126), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT61), .B1(new_n1148), .B2(new_n1122), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT60), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1138), .A2(KEYINPUT60), .A3(new_n1140), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n610), .A2(KEYINPUT122), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n602), .B(KEYINPUT122), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1154), .A2(KEYINPUT60), .A3(new_n1140), .A4(new_n1138), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1149), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1144), .B(KEYINPUT121), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1147), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(G1996), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1013), .A2(new_n1040), .A3(new_n1159), .A4(new_n1042), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT58), .B(G1341), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n1034), .A2(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1161), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n552), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT59), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1143), .B1(new_n1158), .B2(new_n1170), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1082), .A2(new_n1079), .A3(new_n1085), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT123), .B1(new_n1088), .B2(new_n1081), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1077), .ZN(new_n1174));
  OAI22_X1  g749(.A1(new_n1172), .A2(new_n1173), .B1(new_n1174), .B2(new_n1075), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT54), .ZN(new_n1176));
  XNOR2_X1  g751(.A(G171), .B(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1080), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1088), .B1(new_n1043), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(G301), .A2(new_n1176), .ZN(new_n1181));
  NAND2_X1  g756(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1078), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1064), .A2(new_n1070), .A3(new_n1178), .A4(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1020), .ZN(new_n1186));
  INV_X1    g761(.A(new_n997), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1002), .A2(new_n1010), .ZN(new_n1188));
  OAI21_X1  g763(.A(G286), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1189), .A2(G8), .A3(new_n1011), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1186), .B1(new_n1190), .B2(KEYINPUT51), .ZN(new_n1191));
  OAI21_X1  g766(.A(KEYINPUT125), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1175), .A2(new_n1177), .B1(new_n1183), .B2(new_n1078), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1100), .A2(new_n1098), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1102), .B(new_n1114), .C1(new_n1171), .C2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n994), .A2(new_n1006), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1159), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1200), .A2(new_n801), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n708), .B(new_n1135), .ZN(new_n1202));
  INV_X1    g777(.A(new_n801), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1202), .B1(new_n1159), .B2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g779(.A(new_n1198), .B(KEYINPUT105), .Z(new_n1205));
  AOI21_X1  g780(.A(new_n1201), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1205), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n899), .B(new_n748), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g784(.A(G290), .B(G1986), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1209), .B1(new_n1199), .B2(new_n1210), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT106), .Z(new_n1212));
  NAND2_X1  g787(.A1(new_n1197), .A2(new_n1212), .ZN(new_n1213));
  XOR2_X1   g788(.A(new_n1200), .B(KEYINPUT46), .Z(new_n1214));
  NAND2_X1  g789(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1214), .B1(new_n1205), .B2(new_n1215), .ZN(new_n1216));
  XOR2_X1   g791(.A(new_n1216), .B(KEYINPUT47), .Z(new_n1217));
  NOR3_X1   g792(.A1(new_n1198), .A2(G290), .A3(G1986), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1218), .B(KEYINPUT48), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1217), .B1(new_n1209), .B2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1206), .A2(new_n748), .A3(new_n766), .A4(new_n756), .ZN(new_n1221));
  OR2_X1    g796(.A1(new_n708), .A2(G2067), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1207), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n1224));
  AND2_X1   g799(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1226));
  NOR3_X1   g801(.A1(new_n1220), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1213), .A2(new_n1227), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g803(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1230));
  AND3_X1   g804(.A1(new_n684), .A2(new_n687), .A3(new_n1230), .ZN(new_n1231));
  OAI211_X1 g805(.A(new_n1231), .B(new_n924), .C1(new_n988), .C2(new_n989), .ZN(G225));
  INV_X1    g806(.A(G225), .ZN(G308));
endmodule


