//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n196), .B(KEYINPUT77), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT24), .B(G110), .Z(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n194), .A2(G128), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n200), .B(new_n195), .C1(new_n201), .C2(KEYINPUT23), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G110), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT78), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT78), .A2(G125), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n205), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT16), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n209), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(new_n205), .ZN(new_n216));
  AOI21_X1  g030(.A(G146), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT79), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n213), .A2(G146), .A3(new_n216), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n213), .A2(KEYINPUT79), .A3(G146), .A4(new_n216), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n204), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(KEYINPUT80), .B(G110), .Z(new_n223));
  OAI22_X1  g037(.A1(new_n197), .A2(new_n198), .B1(new_n202), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(G125), .A2(G140), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n211), .A2(KEYINPUT81), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT81), .B1(new_n211), .B2(new_n226), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n224), .A2(new_n219), .A3(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT82), .B1(new_n222), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n218), .ZN(new_n232));
  INV_X1    g046(.A(new_n217), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(new_n221), .ZN(new_n234));
  INV_X1    g048(.A(new_n204), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n224), .A2(new_n219), .A3(new_n229), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT22), .B(G137), .ZN(new_n240));
  INV_X1    g054(.A(G953), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n241), .A2(G221), .A3(G234), .ZN(new_n242));
  XOR2_X1   g056(.A(new_n240), .B(new_n242), .Z(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n231), .A2(new_n239), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT83), .B1(new_n246), .B2(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n231), .A2(KEYINPUT83), .A3(new_n239), .A4(new_n244), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n191), .B1(new_n250), .B2(new_n188), .ZN(new_n251));
  AOI211_X1 g065(.A(G902), .B(new_n190), .C1(new_n248), .C2(new_n249), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n189), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n189), .A2(G902), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G472), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G146), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n225), .A2(KEYINPUT65), .A3(G143), .ZN(new_n262));
  AND2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(G146), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n261), .A2(new_n262), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n225), .A2(KEYINPUT64), .A3(G143), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n260), .B2(G146), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n260), .A2(G146), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT0), .B(G128), .ZN(new_n275));
  OAI22_X1  g089(.A1(new_n267), .A2(new_n268), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G137), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT11), .A3(G134), .ZN(new_n278));
  INV_X1    g092(.A(G134), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G137), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n282));
  INV_X1    g096(.A(G131), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT11), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n279), .B2(G137), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n281), .A2(new_n282), .A3(new_n283), .A4(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n285), .A2(new_n278), .A3(new_n283), .A4(new_n280), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n278), .A3(new_n280), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n286), .A2(new_n288), .B1(G131), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(new_n288), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n277), .A2(G134), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n280), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G131), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n225), .A2(G143), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n192), .B1(new_n296), .B2(KEYINPUT1), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT64), .B1(new_n225), .B2(G143), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n296), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n269), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n261), .A2(new_n262), .A3(new_n301), .A4(new_n264), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n295), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  OAI22_X1  g118(.A1(new_n276), .A2(new_n290), .B1(new_n292), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n194), .A2(G116), .ZN(new_n306));
  INV_X1    g120(.A(G116), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G119), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G116), .B(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT68), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT2), .B(G113), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n309), .A2(new_n314), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n258), .B1(new_n305), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G101), .ZN(new_n320));
  NOR2_X1   g134(.A1(G237), .A2(G953), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G210), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n320), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n319), .A2(KEYINPUT29), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT69), .B1(new_n276), .B2(new_n290), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n275), .B1(new_n299), .B2(new_n269), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n261), .A2(new_n262), .A3(new_n264), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT66), .A3(new_n263), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n265), .A2(new_n266), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n289), .A2(G131), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT69), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT1), .ZN(new_n340));
  OAI21_X1  g154(.A(G128), .B1(new_n272), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n273), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n342), .A2(new_n302), .B1(G131), .B2(new_n294), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n318), .B1(new_n343), .B2(new_n291), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n328), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT70), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n328), .A2(new_n339), .A3(new_n344), .A4(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n347), .B1(new_n346), .B2(new_n349), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n343), .A2(new_n291), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n328), .A2(new_n339), .A3(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n353), .A2(new_n318), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n355), .A2(new_n356), .A3(new_n258), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n346), .A2(new_n349), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n358), .B2(KEYINPUT74), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT75), .B1(new_n361), .B2(KEYINPUT28), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n327), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT73), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n325), .B(KEYINPUT72), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n319), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n305), .A2(new_n318), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n358), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n369), .B2(KEYINPUT28), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT30), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n305), .A2(new_n372), .B1(new_n315), .B2(new_n317), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n328), .A2(new_n339), .A3(KEYINPUT30), .A4(new_n352), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n346), .A2(new_n349), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n371), .B1(new_n375), .B2(new_n325), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n364), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n374), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n358), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n325), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n367), .B1(new_n346), .B2(new_n349), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n319), .B(new_n365), .C1(new_n382), .C2(new_n258), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(KEYINPUT73), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(G902), .B1(new_n377), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n257), .B1(new_n363), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT32), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n358), .A2(new_n325), .A3(new_n378), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT31), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n375), .A2(KEYINPUT31), .A3(new_n325), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n319), .B1(new_n382), .B2(new_n258), .ZN(new_n393));
  INV_X1    g207(.A(new_n365), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(G472), .A2(G902), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n387), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n397), .ZN(new_n399));
  AOI211_X1 g213(.A(KEYINPUT32), .B(new_n399), .C1(new_n392), .C2(new_n395), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT76), .B1(new_n386), .B2(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n370), .A2(new_n376), .A3(new_n364), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT73), .B1(new_n381), .B2(new_n383), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n188), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n356), .B1(new_n355), .B2(new_n258), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n361), .A2(KEYINPUT75), .A3(KEYINPUT28), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n326), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G472), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT76), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n390), .A2(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT32), .B1(new_n411), .B2(new_n399), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n396), .A2(new_n387), .A3(new_n397), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n256), .B1(new_n402), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G214), .B1(G237), .B2(G902), .ZN(new_n417));
  OAI21_X1  g231(.A(G210), .B1(G237), .B2(G902), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G122), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OR2_X1    g234(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n421));
  NAND2_X1  g235(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n422));
  INV_X1    g236(.A(G107), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n421), .A2(new_n422), .B1(G104), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(G104), .A3(new_n423), .ZN(new_n425));
  INV_X1    g239(.A(G104), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G107), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G101), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(G104), .ZN(new_n430));
  AND2_X1   g244(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n431));
  NOR2_X1   g245(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G101), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n425), .A4(new_n427), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n429), .A2(KEYINPUT4), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(G101), .C1(new_n424), .C2(new_n428), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n436), .A2(new_n318), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT88), .B(KEYINPUT5), .ZN(new_n440));
  OAI21_X1  g254(.A(G113), .B1(new_n440), .B2(new_n306), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n311), .A2(new_n313), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(new_n440), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n430), .A2(new_n427), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G101), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n435), .A2(new_n445), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n443), .A2(new_n316), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n420), .B1(new_n439), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n442), .A2(new_n440), .ZN(new_n449));
  INV_X1    g263(.A(new_n441), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n435), .A2(new_n445), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n317), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n436), .A2(new_n318), .A3(new_n438), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n419), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n448), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n457), .B(new_n420), .C1(new_n439), .C2(new_n447), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n333), .A2(new_n214), .ZN(new_n459));
  INV_X1    g273(.A(G224), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G953), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n342), .A2(new_n302), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n208), .A3(new_n209), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n459), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n462), .B1(new_n459), .B2(new_n464), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n456), .A2(new_n458), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT89), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n456), .A2(new_n467), .A3(new_n470), .A4(new_n458), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n459), .A2(new_n464), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(KEYINPUT7), .A3(new_n462), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n451), .A2(new_n317), .A3(new_n446), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n441), .B1(KEYINPUT5), .B2(new_n312), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n452), .B1(new_n476), .B2(new_n316), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n419), .B(KEYINPUT8), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n462), .A2(KEYINPUT7), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n459), .A2(new_n464), .A3(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n474), .A2(new_n479), .A3(new_n455), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n188), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n418), .B1(new_n472), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n418), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n486), .B(new_n483), .C1(new_n469), .C2(new_n471), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n417), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G475), .ZN(new_n489));
  INV_X1    g303(.A(G237), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n241), .A3(G214), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n260), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n321), .A2(G143), .A3(G214), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(KEYINPUT90), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(KEYINPUT18), .A2(G131), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n212), .B1(new_n214), .B2(G140), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G146), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n229), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n492), .A2(new_n493), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(KEYINPUT17), .A3(G131), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(G131), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n492), .A2(new_n283), .A3(new_n493), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n502), .B1(new_n505), .B2(KEYINPUT17), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n500), .B1(new_n234), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G113), .B(G122), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT92), .B(G104), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n508), .B(new_n509), .Z(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(new_n500), .C1(new_n234), .C2(new_n506), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n489), .B1(new_n514), .B2(new_n188), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n497), .A2(KEYINPUT19), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n227), .B2(new_n228), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n219), .B(new_n505), .C1(new_n519), .C2(G146), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n500), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT91), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n500), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n511), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n513), .ZN(new_n526));
  NOR2_X1   g340(.A1(G475), .A2(G902), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT20), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT20), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n526), .A2(new_n530), .A3(new_n527), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n515), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n307), .A2(KEYINPUT14), .A3(G122), .ZN(new_n533));
  XNOR2_X1  g347(.A(G116), .B(G122), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(G107), .B(new_n533), .C1(new_n535), .C2(KEYINPUT14), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n423), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n260), .A2(G128), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n260), .A2(G128), .ZN(new_n540));
  OAI21_X1  g354(.A(G134), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n192), .A2(G143), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n538), .A2(new_n542), .A3(new_n279), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n536), .A2(new_n537), .A3(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(KEYINPUT93), .A2(KEYINPUT13), .ZN(new_n546));
  NOR2_X1   g360(.A1(KEYINPUT93), .A2(KEYINPUT13), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT94), .B1(new_n548), .B2(new_n538), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n540), .B1(new_n548), .B2(new_n538), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n539), .B(new_n551), .C1(new_n547), .C2(new_n546), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G134), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n543), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n543), .A2(new_n555), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n535), .A2(G107), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n556), .A2(new_n557), .B1(new_n558), .B2(new_n537), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT96), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n554), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n554), .B2(new_n559), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n545), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT9), .B(G234), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n565), .A2(new_n187), .A3(G953), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n554), .A2(new_n559), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT96), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n561), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n545), .A3(new_n566), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G478), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n573), .B(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G952), .ZN(new_n577));
  AOI211_X1 g391(.A(G953), .B(new_n577), .C1(G234), .C2(G237), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n188), .B(new_n241), .C1(G234), .C2(G237), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT21), .B(G898), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n532), .A2(new_n576), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G221), .B1(new_n565), .B2(G902), .ZN(new_n584));
  INV_X1    g398(.A(G469), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n436), .A2(new_n438), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n302), .B1(new_n330), .B2(new_n297), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n452), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n586), .A2(new_n333), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n452), .A2(new_n463), .A3(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT87), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT87), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n452), .A2(new_n463), .A3(new_n593), .A4(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n290), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n590), .A2(new_n595), .A3(new_n290), .ZN(new_n598));
  XNOR2_X1  g412(.A(G110), .B(G140), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT85), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n241), .A2(G227), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n600), .B(new_n601), .Z(new_n602));
  NAND3_X1  g416(.A1(new_n597), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n602), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n590), .A2(new_n595), .A3(new_n290), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n446), .A2(new_n342), .A3(new_n302), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n589), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n607), .A2(KEYINPUT12), .A3(new_n337), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT12), .B1(new_n607), .B2(new_n337), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n604), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n603), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n585), .B1(new_n612), .B2(new_n188), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n604), .B1(new_n605), .B2(new_n596), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n598), .B(new_n602), .C1(new_n608), .C2(new_n609), .ZN(new_n615));
  AOI211_X1 g429(.A(G469), .B(G902), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n584), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n488), .A2(new_n583), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n416), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  AOI21_X1  g434(.A(new_n257), .B1(new_n396), .B2(new_n188), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n396), .A2(new_n397), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n617), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n253), .A3(new_n255), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n417), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n472), .A2(new_n484), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n486), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n472), .A2(new_n418), .A3(new_n484), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n574), .A2(new_n188), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n573), .B2(new_n574), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n566), .B1(new_n571), .B2(new_n545), .ZN(new_n635));
  INV_X1    g449(.A(new_n545), .ZN(new_n636));
  AOI211_X1 g450(.A(new_n636), .B(new_n567), .C1(new_n570), .C2(new_n561), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT33), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n568), .A2(new_n572), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n638), .A2(G478), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT97), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n634), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n532), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n632), .A2(new_n646), .A3(KEYINPUT98), .A4(new_n582), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n582), .B(new_n417), .C1(new_n485), .C2(new_n487), .ZN(new_n649));
  INV_X1    g463(.A(new_n515), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n530), .B1(new_n526), .B2(new_n527), .ZN(new_n651));
  INV_X1    g465(.A(new_n527), .ZN(new_n652));
  AOI211_X1 g466(.A(KEYINPUT20), .B(new_n652), .C1(new_n525), .C2(new_n513), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n650), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n634), .A2(new_n641), .A3(new_n644), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n644), .B1(new_n634), .B2(new_n641), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n648), .B1(new_n649), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n647), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n627), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT34), .B(G104), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  INV_X1    g477(.A(new_n575), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n573), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n532), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n663), .B1(new_n666), .B2(new_n581), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n654), .A2(new_n576), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(KEYINPUT99), .A3(new_n582), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n632), .A3(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n670), .A2(new_n624), .A3(new_n626), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT100), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT35), .B(G107), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  NAND2_X1  g488(.A1(new_n231), .A2(new_n239), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n244), .A2(KEYINPUT36), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n675), .B(new_n676), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n254), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n253), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n625), .A3(new_n632), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n624), .A2(new_n583), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT101), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n683), .B(new_n685), .ZN(G12));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n579), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n578), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n668), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n680), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n409), .A2(new_n410), .A3(new_n414), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n410), .B1(new_n409), .B2(new_n414), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  NOR2_X1   g510(.A1(new_n485), .A2(new_n487), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT38), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT40), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n690), .B(KEYINPUT39), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n625), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n698), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n388), .B1(new_n355), .B2(new_n365), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n257), .B1(new_n704), .B2(new_n188), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n412), .B2(new_n413), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n679), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n654), .A2(new_n665), .ZN(new_n708));
  AOI211_X1 g522(.A(new_n628), .B(new_n708), .C1(new_n701), .C2(KEYINPUT40), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n703), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  NAND2_X1  g525(.A1(new_n402), .A2(new_n415), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n632), .A2(new_n646), .A3(new_n713), .A4(new_n690), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n654), .B(new_n690), .C1(new_n655), .C2(new_n656), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT102), .B1(new_n715), .B2(new_n488), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n617), .B1(new_n253), .B2(new_n678), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  INV_X1    g534(.A(new_n256), .ZN(new_n721));
  INV_X1    g535(.A(new_n616), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n614), .A2(new_n615), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n188), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n584), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n647), .B2(new_n658), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n712), .A2(new_n721), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  NOR2_X1   g547(.A1(new_n670), .A2(new_n729), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n734), .B(new_n721), .C1(new_n693), .C2(new_n694), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  NOR3_X1   g550(.A1(new_n729), .A2(new_n583), .A3(new_n488), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n679), .B(new_n737), .C1(new_n693), .C2(new_n694), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  NAND4_X1  g553(.A1(new_n632), .A2(KEYINPUT103), .A3(new_n665), .A4(new_n654), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n488), .B2(new_n708), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n729), .A2(new_n581), .ZN(new_n744));
  INV_X1    g558(.A(new_n319), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n406), .B2(new_n407), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n392), .B1(new_n746), .B2(new_n365), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n621), .B1(new_n747), .B2(new_n397), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n743), .A2(new_n744), .A3(new_n748), .A4(new_n721), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT104), .B(G122), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G24));
  INV_X1    g565(.A(new_n715), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n488), .A2(new_n726), .A3(new_n727), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n748), .A2(new_n679), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  AOI21_X1  g569(.A(new_n386), .B1(KEYINPUT106), .B2(new_n414), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n401), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n256), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n630), .A2(new_n417), .A3(new_n631), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n715), .A2(new_n760), .A3(new_n617), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(KEYINPUT42), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n712), .A2(new_n763), .A3(new_n721), .A4(new_n761), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n763), .B1(new_n416), .B2(new_n761), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G131), .ZN(G33));
  NOR3_X1   g583(.A1(new_n691), .A2(new_n760), .A3(new_n617), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n721), .B(new_n770), .C1(new_n693), .C2(new_n694), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n416), .A2(KEYINPUT107), .A3(new_n770), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  OAI21_X1  g590(.A(new_n532), .B1(new_n655), .B2(new_n656), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT43), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(KEYINPUT43), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n624), .A3(new_n679), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n612), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n603), .A2(new_n611), .A3(KEYINPUT45), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(G469), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(G469), .A2(G902), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT46), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n616), .A2(KEYINPUT46), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n787), .A3(new_n788), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n584), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n760), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n700), .A3(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n782), .A2(new_n783), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n277), .ZN(G39));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n790), .A2(KEYINPUT47), .A3(new_n584), .A4(new_n792), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n721), .A2(new_n715), .A3(new_n760), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT108), .B1(new_n804), .B2(new_n712), .ZN(new_n805));
  INV_X1    g619(.A(new_n712), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n806), .A2(new_n802), .A3(new_n807), .A4(new_n803), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  AND3_X1   g624(.A1(new_n778), .A2(new_n578), .A3(new_n779), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n729), .A2(new_n760), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n759), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT48), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n813), .A2(KEYINPUT114), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n811), .A2(new_n721), .A3(new_n748), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n815), .B1(new_n753), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n721), .A2(new_n812), .A3(new_n578), .A4(new_n706), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n646), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(G952), .A3(new_n241), .ZN(new_n822));
  XNOR2_X1  g636(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(new_n813), .B2(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n818), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n819), .B1(new_n818), .B2(new_n824), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n698), .A2(new_n628), .A3(new_n728), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT112), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OR4_X1    g645(.A1(KEYINPUT113), .A2(new_n831), .A3(KEYINPUT50), .A4(new_n816), .ZN(new_n832));
  XOR2_X1   g646(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n831), .B2(new_n816), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n820), .A2(new_n532), .A3(new_n645), .A4(new_n643), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n811), .A2(new_n812), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n747), .A2(new_n397), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n622), .A3(new_n679), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n835), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n800), .B(new_n801), .C1(new_n584), .C2(new_n726), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n840), .A2(new_n795), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n841), .B2(new_n817), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n832), .A2(new_n834), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n827), .B1(new_n828), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n828), .B2(new_n843), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n743), .A2(new_n707), .A3(new_n625), .A4(new_n690), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n719), .A2(new_n695), .A3(new_n847), .A4(new_n754), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT52), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n712), .B1(new_n718), .B2(new_n692), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n754), .A4(new_n847), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n849), .A2(KEYINPUT110), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT110), .B1(new_n849), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n731), .A2(new_n735), .A3(new_n738), .A4(new_n749), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n646), .A2(new_n668), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n649), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n681), .A2(new_n682), .B1(new_n627), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n619), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT109), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n532), .A2(new_n576), .A3(new_n690), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n862), .B1(new_n760), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n690), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n654), .A2(new_n665), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n697), .A3(KEYINPUT109), .A4(new_n417), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n864), .A2(new_n717), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n693), .B2(new_n694), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n748), .A2(new_n761), .A3(new_n679), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n773), .B2(new_n774), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n861), .A2(new_n768), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n846), .B1(new_n855), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT111), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n731), .A2(new_n735), .A3(new_n738), .A4(new_n749), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n619), .A2(KEYINPUT53), .A3(new_n859), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n768), .A2(new_n876), .A3(new_n872), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n849), .A2(new_n852), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n875), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n872), .A2(new_n876), .A3(new_n877), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n717), .A2(new_n632), .A3(new_n668), .A4(new_n690), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n882), .A2(new_n883), .B1(new_n402), .B2(new_n415), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n753), .A2(new_n752), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n838), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n851), .B1(new_n887), .B2(new_n847), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n851), .A2(new_n850), .A3(new_n754), .A4(new_n847), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n881), .A2(KEYINPUT111), .A3(new_n768), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n874), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT53), .B1(new_n855), .B2(new_n873), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n890), .A2(new_n846), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n895), .B1(new_n873), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n894), .B1(new_n897), .B2(new_n893), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n845), .A2(new_n898), .B1(G952), .B2(G953), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n726), .A2(KEYINPUT49), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n726), .A2(KEYINPUT49), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n584), .A2(new_n417), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n777), .A4(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(new_n721), .A3(new_n706), .A4(new_n698), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n899), .A2(new_n904), .ZN(G75));
  NOR2_X1   g719(.A1(new_n241), .A2(G952), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n188), .B1(new_n874), .B2(new_n892), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT56), .B1(new_n908), .B2(G210), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n456), .A2(new_n458), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(new_n467), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT55), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n907), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n908), .B2(G210), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(KEYINPUT116), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(KEYINPUT116), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(G51));
  XOR2_X1   g733(.A(new_n788), .B(KEYINPUT57), .Z(new_n920));
  INV_X1    g734(.A(new_n894), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n893), .B1(new_n874), .B2(new_n892), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n723), .B(KEYINPUT117), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n908), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n926), .A2(new_n787), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n906), .B1(new_n925), .B2(new_n927), .ZN(G54));
  NAND3_X1  g742(.A1(new_n908), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n513), .A3(new_n525), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n908), .A2(KEYINPUT58), .A3(G475), .A4(new_n526), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n930), .A2(new_n907), .A3(new_n931), .ZN(G60));
  NAND2_X1  g746(.A1(new_n638), .A2(new_n640), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n633), .B(KEYINPUT59), .Z(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n898), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  INV_X1    g750(.A(new_n922), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(new_n894), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n935), .A2(new_n938), .A3(new_n906), .ZN(G63));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n874), .B2(new_n892), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n677), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n907), .B1(new_n943), .B2(new_n250), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n940), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n943), .A2(new_n250), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n948), .A2(KEYINPUT61), .A3(new_n907), .A4(new_n944), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(G66));
  OAI21_X1  g764(.A(new_n241), .B1(new_n856), .B2(new_n860), .ZN(new_n951));
  OAI21_X1  g765(.A(G953), .B1(new_n580), .B2(new_n460), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n951), .A2(KEYINPUT118), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(KEYINPUT118), .B2(new_n951), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n910), .B1(G898), .B2(new_n241), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT119), .Z(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G69));
  AOI21_X1  g771(.A(new_n241), .B1(G227), .B2(G900), .ZN(new_n958));
  INV_X1    g772(.A(new_n305), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n374), .B1(KEYINPUT30), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT120), .Z(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n519), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n797), .B1(new_n808), .B2(new_n805), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n759), .A2(new_n700), .A3(new_n743), .A4(new_n794), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n887), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(new_n768), .A3(new_n775), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n241), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n241), .A2(G900), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT122), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n962), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(KEYINPUT124), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n887), .A2(new_n973), .A3(new_n710), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT121), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n857), .A2(new_n701), .A3(new_n760), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n416), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n887), .A2(new_n710), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n963), .B(new_n977), .C1(new_n973), .C2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n962), .B1(new_n980), .B2(G953), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT124), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n970), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n958), .B1(new_n972), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(KEYINPUT125), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n986), .B(new_n958), .C1(new_n972), .C2(new_n983), .ZN(new_n987));
  INV_X1    g801(.A(new_n958), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n971), .A2(new_n981), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT123), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n971), .A2(new_n981), .A3(KEYINPUT123), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n985), .A2(new_n987), .A3(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(new_n379), .A2(new_n380), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n388), .ZN(new_n996));
  XNOR2_X1  g810(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n257), .A2(new_n188), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n907), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n996), .A2(new_n999), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT127), .Z(new_n1002));
  NOR2_X1   g816(.A1(new_n897), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n980), .A2(new_n325), .A3(new_n379), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n375), .A2(new_n380), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n966), .B2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g820(.A(new_n1000), .B(new_n1003), .C1(new_n861), .C2(new_n1006), .ZN(G57));
endmodule


