

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595;

  INV_X1 U328 ( .A(KEYINPUT82), .ZN(n318) );
  XNOR2_X1 U329 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U330 ( .A(n447), .B(n320), .ZN(n324) );
  XNOR2_X1 U331 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n402) );
  XNOR2_X1 U332 ( .A(n403), .B(n402), .ZN(n537) );
  XNOR2_X1 U333 ( .A(n467), .B(G190GAT), .ZN(n468) );
  XNOR2_X1 U334 ( .A(n469), .B(n468), .ZN(G1351GAT) );
  XOR2_X1 U335 ( .A(G176GAT), .B(KEYINPUT89), .Z(n297) );
  XNOR2_X1 U336 ( .A(G169GAT), .B(KEYINPUT90), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U338 ( .A(KEYINPUT67), .B(KEYINPUT20), .Z(n299) );
  XNOR2_X1 U339 ( .A(G15GAT), .B(KEYINPUT91), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U341 ( .A(n301), .B(n300), .Z(n307) );
  XOR2_X1 U342 ( .A(G183GAT), .B(KEYINPUT17), .Z(n303) );
  XNOR2_X1 U343 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n302) );
  XNOR2_X1 U344 ( .A(n303), .B(n302), .ZN(n414) );
  XOR2_X1 U345 ( .A(G127GAT), .B(KEYINPUT0), .Z(n305) );
  XNOR2_X1 U346 ( .A(G113GAT), .B(KEYINPUT88), .ZN(n304) );
  XNOR2_X1 U347 ( .A(n305), .B(n304), .ZN(n420) );
  XNOR2_X1 U348 ( .A(n414), .B(n420), .ZN(n306) );
  XNOR2_X1 U349 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U350 ( .A(G190GAT), .B(G134GAT), .Z(n328) );
  XOR2_X1 U351 ( .A(G120GAT), .B(G71GAT), .Z(n356) );
  XOR2_X1 U352 ( .A(n328), .B(n356), .Z(n309) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U355 ( .A(n311), .B(n310), .Z(n313) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G99GAT), .ZN(n312) );
  XOR2_X1 U357 ( .A(n313), .B(n312), .Z(n538) );
  INV_X1 U358 ( .A(n538), .ZN(n504) );
  INV_X1 U359 ( .A(KEYINPUT83), .ZN(n332) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n314), .B(G29GAT), .ZN(n315) );
  XOR2_X1 U362 ( .A(n315), .B(KEYINPUT8), .Z(n317) );
  XNOR2_X1 U363 ( .A(G43GAT), .B(G50GAT), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n317), .B(n316), .ZN(n384) );
  XOR2_X1 U365 ( .A(G218GAT), .B(G162GAT), .Z(n447) );
  NAND2_X1 U366 ( .A1(G232GAT), .A2(G233GAT), .ZN(n319) );
  XOR2_X1 U367 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n322) );
  XNOR2_X1 U368 ( .A(KEYINPUT81), .B(KEYINPUT10), .ZN(n321) );
  XNOR2_X1 U369 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U370 ( .A(n324), .B(n323), .Z(n330) );
  XOR2_X1 U371 ( .A(KEYINPUT79), .B(G92GAT), .Z(n326) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(G85GAT), .ZN(n325) );
  XNOR2_X1 U373 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(n327), .ZN(n369) );
  XOR2_X1 U375 ( .A(n328), .B(n369), .Z(n329) );
  XNOR2_X1 U376 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U377 ( .A(n384), .B(n331), .ZN(n395) );
  XNOR2_X1 U378 ( .A(n332), .B(n395), .ZN(n466) );
  XOR2_X1 U379 ( .A(n466), .B(KEYINPUT104), .Z(n333) );
  XNOR2_X1 U380 ( .A(n333), .B(KEYINPUT36), .ZN(n593) );
  XOR2_X1 U381 ( .A(KEYINPUT15), .B(KEYINPUT87), .Z(n335) );
  XNOR2_X1 U382 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n354) );
  XOR2_X1 U384 ( .A(G78GAT), .B(G71GAT), .Z(n337) );
  XNOR2_X1 U385 ( .A(G22GAT), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U386 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U387 ( .A(KEYINPUT86), .B(G64GAT), .Z(n339) );
  XNOR2_X1 U388 ( .A(G8GAT), .B(G127GAT), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U390 ( .A(n341), .B(n340), .Z(n347) );
  XNOR2_X1 U391 ( .A(G57GAT), .B(KEYINPUT76), .ZN(n342) );
  XNOR2_X1 U392 ( .A(n342), .B(KEYINPUT13), .ZN(n357) );
  XOR2_X1 U393 ( .A(n357), .B(G211GAT), .Z(n344) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U396 ( .A(G155GAT), .B(n345), .ZN(n346) );
  XNOR2_X1 U397 ( .A(n347), .B(n346), .ZN(n349) );
  INV_X1 U398 ( .A(KEYINPUT14), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n349), .B(n348), .ZN(n352) );
  XNOR2_X1 U400 ( .A(G15GAT), .B(G1GAT), .ZN(n350) );
  XNOR2_X1 U401 ( .A(n350), .B(KEYINPUT72), .ZN(n376) );
  XNOR2_X1 U402 ( .A(n376), .B(KEYINPUT12), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U404 ( .A(n354), .B(n353), .Z(n545) );
  INV_X1 U405 ( .A(n545), .ZN(n561) );
  NOR2_X1 U406 ( .A1(n593), .A2(n561), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n355), .B(KEYINPUT45), .ZN(n389) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n359) );
  AND2_X1 U409 ( .A1(G230GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U410 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U411 ( .A(KEYINPUT77), .B(KEYINPUT33), .Z(n361) );
  XNOR2_X1 U412 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n360) );
  XOR2_X1 U413 ( .A(n361), .B(n360), .Z(n362) );
  XNOR2_X1 U414 ( .A(n363), .B(n362), .ZN(n368) );
  XOR2_X1 U415 ( .A(G78GAT), .B(G148GAT), .Z(n365) );
  XNOR2_X1 U416 ( .A(KEYINPUT78), .B(G204GAT), .ZN(n364) );
  XNOR2_X1 U417 ( .A(n365), .B(n364), .ZN(n446) );
  XNOR2_X1 U418 ( .A(G176GAT), .B(G64GAT), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n366), .B(KEYINPUT80), .ZN(n413) );
  XNOR2_X1 U420 ( .A(n446), .B(n413), .ZN(n367) );
  XOR2_X1 U421 ( .A(n368), .B(n367), .Z(n370) );
  XNOR2_X1 U422 ( .A(n370), .B(n369), .ZN(n585) );
  XOR2_X1 U423 ( .A(KEYINPUT74), .B(KEYINPUT69), .Z(n372) );
  XNOR2_X1 U424 ( .A(KEYINPUT71), .B(KEYINPUT73), .ZN(n371) );
  XNOR2_X1 U425 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U426 ( .A(n373), .B(G113GAT), .Z(n375) );
  XNOR2_X1 U427 ( .A(G169GAT), .B(G8GAT), .ZN(n404) );
  XOR2_X1 U428 ( .A(n404), .B(G197GAT), .Z(n374) );
  XNOR2_X1 U429 ( .A(n375), .B(n374), .ZN(n380) );
  XOR2_X1 U430 ( .A(G141GAT), .B(G22GAT), .Z(n453) );
  XOR2_X1 U431 ( .A(n453), .B(n376), .Z(n378) );
  NAND2_X1 U432 ( .A1(G229GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U434 ( .A(n380), .B(n379), .Z(n386) );
  XOR2_X1 U435 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n382) );
  XNOR2_X1 U436 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U439 ( .A(n386), .B(n385), .Z(n512) );
  XNOR2_X1 U440 ( .A(n512), .B(KEYINPUT75), .ZN(n568) );
  INV_X1 U441 ( .A(n568), .ZN(n387) );
  AND2_X1 U442 ( .A1(n585), .A2(n387), .ZN(n388) );
  AND2_X1 U443 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U444 ( .A(n390), .B(KEYINPUT114), .ZN(n401) );
  INV_X1 U445 ( .A(n512), .ZN(n582) );
  XNOR2_X1 U446 ( .A(n585), .B(KEYINPUT65), .ZN(n392) );
  INV_X1 U447 ( .A(KEYINPUT41), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n570) );
  NAND2_X1 U449 ( .A1(n582), .A2(n570), .ZN(n394) );
  INV_X1 U450 ( .A(KEYINPUT46), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n398) );
  INV_X1 U452 ( .A(n395), .ZN(n396) );
  NAND2_X1 U453 ( .A1(n561), .A2(n396), .ZN(n397) );
  NOR2_X1 U454 ( .A1(n398), .A2(n397), .ZN(n399) );
  XOR2_X1 U455 ( .A(KEYINPUT47), .B(n399), .Z(n400) );
  NOR2_X1 U456 ( .A1(n401), .A2(n400), .ZN(n403) );
  XNOR2_X1 U457 ( .A(G36GAT), .B(G218GAT), .ZN(n405) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n418) );
  XNOR2_X1 U459 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n406), .B(G211GAT), .ZN(n457) );
  XOR2_X1 U461 ( .A(KEYINPUT101), .B(n457), .Z(n408) );
  NAND2_X1 U462 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U464 ( .A(KEYINPUT84), .B(G92GAT), .Z(n410) );
  XNOR2_X1 U465 ( .A(G190GAT), .B(G204GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U467 ( .A(n412), .B(n411), .Z(n416) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U469 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U470 ( .A(n418), .B(n417), .Z(n528) );
  INV_X1 U471 ( .A(n528), .ZN(n502) );
  NOR2_X1 U472 ( .A1(n537), .A2(n502), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n419), .B(KEYINPUT54), .ZN(n444) );
  XOR2_X1 U474 ( .A(G85GAT), .B(n420), .Z(n422) );
  NAND2_X1 U475 ( .A1(G225GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n443) );
  XOR2_X1 U477 ( .A(G57GAT), .B(G120GAT), .Z(n424) );
  XNOR2_X1 U478 ( .A(G141GAT), .B(G1GAT), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U480 ( .A(KEYINPUT82), .B(G148GAT), .Z(n426) );
  XNOR2_X1 U481 ( .A(G134GAT), .B(G162GAT), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n440) );
  XOR2_X1 U484 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n430) );
  XNOR2_X1 U485 ( .A(KEYINPUT4), .B(KEYINPUT100), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U487 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n432) );
  XNOR2_X1 U488 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U491 ( .A(KEYINPUT92), .B(KEYINPUT2), .Z(n436) );
  XNOR2_X1 U492 ( .A(KEYINPUT93), .B(G155GAT), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U494 ( .A(KEYINPUT3), .B(n437), .ZN(n462) );
  XNOR2_X1 U495 ( .A(n438), .B(n462), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U497 ( .A(G29GAT), .B(n441), .Z(n442) );
  XOR2_X1 U498 ( .A(n443), .B(n442), .Z(n526) );
  INV_X1 U499 ( .A(n526), .ZN(n499) );
  NAND2_X1 U500 ( .A1(n444), .A2(n499), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n445), .B(KEYINPUT66), .ZN(n581) );
  XOR2_X1 U502 ( .A(n447), .B(n446), .Z(n449) );
  NAND2_X1 U503 ( .A1(G228GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(n461) );
  XOR2_X1 U505 ( .A(KEYINPUT94), .B(KEYINPUT22), .Z(n451) );
  XNOR2_X1 U506 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U508 ( .A(n452), .B(G106GAT), .Z(n455) );
  XNOR2_X1 U509 ( .A(G50GAT), .B(n453), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U511 ( .A(n456), .B(KEYINPUT23), .Z(n459) );
  XNOR2_X1 U512 ( .A(n457), .B(KEYINPUT96), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n461), .B(n460), .ZN(n463) );
  XNOR2_X1 U515 ( .A(n463), .B(n462), .ZN(n479) );
  NOR2_X1 U516 ( .A1(n581), .A2(n479), .ZN(n464) );
  XNOR2_X1 U517 ( .A(n464), .B(KEYINPUT55), .ZN(n465) );
  NOR2_X2 U518 ( .A1(n504), .A2(n465), .ZN(n575) );
  NAND2_X1 U519 ( .A1(n575), .A2(n466), .ZN(n469) );
  XOR2_X1 U520 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n467) );
  XNOR2_X1 U521 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n486) );
  NAND2_X1 U522 ( .A1(n568), .A2(n585), .ZN(n496) );
  NOR2_X1 U523 ( .A1(n561), .A2(n466), .ZN(n470) );
  XNOR2_X1 U524 ( .A(n470), .B(KEYINPUT16), .ZN(n484) );
  NOR2_X1 U525 ( .A1(n504), .A2(n502), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n479), .A2(n471), .ZN(n472) );
  XOR2_X1 U527 ( .A(KEYINPUT25), .B(n472), .Z(n475) );
  NAND2_X1 U528 ( .A1(n479), .A2(n504), .ZN(n473) );
  XOR2_X1 U529 ( .A(n473), .B(KEYINPUT26), .Z(n554) );
  INV_X1 U530 ( .A(n554), .ZN(n580) );
  XOR2_X1 U531 ( .A(n528), .B(KEYINPUT27), .Z(n477) );
  NOR2_X1 U532 ( .A1(n580), .A2(n477), .ZN(n474) );
  NOR2_X1 U533 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U534 ( .A1(n526), .A2(n476), .ZN(n482) );
  NOR2_X1 U535 ( .A1(n499), .A2(n477), .ZN(n478) );
  XOR2_X1 U536 ( .A(KEYINPUT102), .B(n478), .Z(n536) );
  XOR2_X1 U537 ( .A(KEYINPUT28), .B(n479), .Z(n508) );
  NAND2_X1 U538 ( .A1(n508), .A2(n504), .ZN(n480) );
  NOR2_X1 U539 ( .A1(n536), .A2(n480), .ZN(n481) );
  NOR2_X1 U540 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U541 ( .A(KEYINPUT103), .B(n483), .ZN(n493) );
  NAND2_X1 U542 ( .A1(n484), .A2(n493), .ZN(n513) );
  NOR2_X1 U543 ( .A1(n496), .A2(n513), .ZN(n490) );
  NAND2_X1 U544 ( .A1(n490), .A2(n526), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(G1324GAT) );
  NAND2_X1 U546 ( .A1(n528), .A2(n490), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n487), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .Z(n489) );
  NAND2_X1 U549 ( .A1(n490), .A2(n538), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  INV_X1 U551 ( .A(n508), .ZN(n541) );
  NAND2_X1 U552 ( .A1(n490), .A2(n541), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT106), .Z(n492) );
  XNOR2_X1 U555 ( .A(KEYINPUT39), .B(n492), .ZN(n501) );
  NAND2_X1 U556 ( .A1(n561), .A2(n493), .ZN(n494) );
  NOR2_X1 U557 ( .A1(n593), .A2(n494), .ZN(n495) );
  XNOR2_X1 U558 ( .A(KEYINPUT37), .B(n495), .ZN(n525) );
  NOR2_X1 U559 ( .A1(n525), .A2(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(KEYINPUT38), .B(KEYINPUT105), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n509) );
  NOR2_X1 U562 ( .A1(n499), .A2(n509), .ZN(n500) );
  XOR2_X1 U563 ( .A(n501), .B(n500), .Z(G1328GAT) );
  NOR2_X1 U564 ( .A1(n502), .A2(n509), .ZN(n503) );
  XOR2_X1 U565 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  XNOR2_X1 U566 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n506) );
  NOR2_X1 U567 ( .A1(n504), .A2(n509), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NOR2_X1 U570 ( .A1(n509), .A2(n508), .ZN(n510) );
  XOR2_X1 U571 ( .A(KEYINPUT108), .B(n510), .Z(n511) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(n511), .ZN(G1331GAT) );
  NAND2_X1 U573 ( .A1(n570), .A2(n512), .ZN(n524) );
  NOR2_X1 U574 ( .A1(n524), .A2(n513), .ZN(n514) );
  XOR2_X1 U575 ( .A(KEYINPUT109), .B(n514), .Z(n520) );
  NAND2_X1 U576 ( .A1(n520), .A2(n526), .ZN(n515) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(n515), .ZN(n516) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(n516), .ZN(G1332GAT) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(KEYINPUT110), .ZN(n518) );
  NAND2_X1 U580 ( .A1(n520), .A2(n528), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n538), .A2(n520), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n522) );
  NAND2_X1 U585 ( .A1(n520), .A2(n541), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U587 ( .A(G78GAT), .B(n523), .Z(G1335GAT) );
  NOR2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n532), .A2(n526), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n527), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n528), .A2(n532), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n529), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n538), .A2(n532), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(KEYINPUT112), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n534) );
  NAND2_X1 U597 ( .A1(n532), .A2(n541), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n553) );
  NAND2_X1 U601 ( .A1(n553), .A2(n538), .ZN(n539) );
  XOR2_X1 U602 ( .A(KEYINPUT115), .B(n539), .Z(n540) );
  NOR2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n549), .A2(n568), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U607 ( .A1(n549), .A2(n570), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n547) );
  NAND2_X1 U610 ( .A1(n549), .A2(n545), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U612 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n551) );
  NAND2_X1 U614 ( .A1(n549), .A2(n466), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U616 ( .A(G134GAT), .B(n552), .Z(G1343GAT) );
  XOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT119), .Z(n557) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U619 ( .A(KEYINPUT118), .B(n555), .Z(n565) );
  NAND2_X1 U620 ( .A1(n582), .A2(n565), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  NAND2_X1 U623 ( .A1(n570), .A2(n565), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n563) );
  INV_X1 U627 ( .A(n561), .ZN(n588) );
  NAND2_X1 U628 ( .A1(n588), .A2(n565), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(n564), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n395), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT122), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n575), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G169GAT), .B(n569), .ZN(G1348GAT) );
  NAND2_X1 U636 ( .A1(n575), .A2(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n574) );
  XOR2_X1 U639 ( .A(G176GAT), .B(KEYINPUT56), .Z(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  NAND2_X1 U641 ( .A1(n575), .A2(n588), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n576), .B(KEYINPUT124), .ZN(n577) );
  XNOR2_X1 U643 ( .A(G183GAT), .B(n577), .ZN(G1350GAT) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(KEYINPUT126), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT60), .B(n579), .Z(n584) );
  NOR2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n589) );
  NAND2_X1 U648 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .Z(n587) );
  INV_X1 U651 ( .A(n589), .ZN(n592) );
  OR2_X1 U652 ( .A1(n592), .A2(n585), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  XOR2_X1 U654 ( .A(G211GAT), .B(KEYINPUT127), .Z(n591) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1354GAT) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(n594), .Z(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

