

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777;

  XNOR2_X1 U374 ( .A(n577), .B(KEYINPUT32), .ZN(n578) );
  XNOR2_X1 U375 ( .A(n430), .B(KEYINPUT101), .ZN(n675) );
  XNOR2_X2 U376 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X2 U377 ( .A(n352), .B(n495), .ZN(n764) );
  NAND2_X1 U378 ( .A1(n413), .A2(n412), .ZN(n352) );
  NAND2_X1 U379 ( .A1(n353), .A2(n581), .ZN(n459) );
  INV_X1 U380 ( .A(n584), .ZN(n353) );
  XNOR2_X2 U381 ( .A(n579), .B(KEYINPUT82), .ZN(n584) );
  XNOR2_X2 U382 ( .A(n564), .B(KEYINPUT91), .ZN(n554) );
  NOR2_X2 U383 ( .A1(n429), .A2(n675), .ZN(n699) );
  XOR2_X1 U384 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n354) );
  XOR2_X1 U385 ( .A(n610), .B(KEYINPUT71), .Z(n355) );
  XNOR2_X2 U386 ( .A(n592), .B(KEYINPUT75), .ZN(n674) );
  INV_X1 U387 ( .A(n680), .ZN(n429) );
  NAND2_X1 U388 ( .A1(n641), .A2(n688), .ZN(n428) );
  NOR2_X1 U389 ( .A1(n409), .A2(n709), .ZN(n596) );
  INV_X1 U390 ( .A(n560), .ZN(n556) );
  XNOR2_X1 U391 ( .A(n389), .B(n390), .ZN(n386) );
  NOR2_X2 U392 ( .A1(n554), .A2(n692), .ZN(n374) );
  AND2_X1 U393 ( .A1(n365), .A2(n695), .ZN(n615) );
  INV_X1 U394 ( .A(n715), .ZN(n402) );
  NOR2_X1 U395 ( .A1(n597), .A2(n598), .ZN(n365) );
  XNOR2_X1 U396 ( .A(n555), .B(KEYINPUT100), .ZN(n680) );
  NAND2_X1 U397 ( .A1(n556), .A2(n559), .ZN(n555) );
  XNOR2_X1 U398 ( .A(n386), .B(n384), .ZN(n383) );
  XNOR2_X1 U399 ( .A(n396), .B(G125), .ZN(n504) );
  INV_X1 U400 ( .A(G953), .ZN(n388) );
  INV_X1 U401 ( .A(G146), .ZN(n396) );
  INV_X1 U402 ( .A(G953), .ZN(n405) );
  INV_X1 U403 ( .A(KEYINPUT88), .ZN(n385) );
  INV_X1 U404 ( .A(KEYINPUT66), .ZN(n404) );
  NOR2_X1 U405 ( .A1(n359), .A2(n356), .ZN(n421) );
  NAND2_X1 U406 ( .A1(n364), .A2(n363), .ZN(n362) );
  XNOR2_X1 U407 ( .A(n569), .B(KEYINPUT105), .ZN(n774) );
  NAND2_X1 U408 ( .A1(n398), .A2(n654), .ZN(n603) );
  XNOR2_X1 U409 ( .A(n401), .B(n354), .ZN(n683) );
  AND2_X1 U410 ( .A1(n377), .A2(n376), .ZN(n375) );
  NAND2_X1 U411 ( .A1(n553), .A2(n402), .ZN(n401) );
  NAND2_X1 U412 ( .A1(n400), .A2(n674), .ZN(n399) );
  OR2_X1 U413 ( .A1(n724), .A2(n444), .ZN(n613) );
  INV_X1 U414 ( .A(n699), .ZN(n400) );
  NAND2_X1 U415 ( .A1(n369), .A2(n368), .ZN(n367) );
  AND2_X1 U416 ( .A1(n372), .A2(n371), .ZN(n370) );
  INV_X1 U417 ( .A(n567), .ZN(n369) );
  XNOR2_X1 U418 ( .A(n601), .B(KEYINPUT38), .ZN(n695) );
  NOR2_X1 U419 ( .A1(n709), .A2(KEYINPUT108), .ZN(n368) );
  NAND2_X1 U420 ( .A1(n709), .A2(KEYINPUT108), .ZN(n371) );
  XNOR2_X1 U421 ( .A(n397), .B(n393), .ZN(n745) );
  XNOR2_X1 U422 ( .A(n383), .B(n382), .ZN(n423) );
  XNOR2_X1 U423 ( .A(n511), .B(n510), .ZN(n397) );
  XNOR2_X1 U424 ( .A(n763), .B(n394), .ZN(n393) );
  XNOR2_X1 U425 ( .A(n392), .B(G134), .ZN(n531) );
  XNOR2_X1 U426 ( .A(n387), .B(n385), .ZN(n384) );
  XNOR2_X1 U427 ( .A(n504), .B(n395), .ZN(n763) );
  XNOR2_X1 U428 ( .A(n403), .B(G137), .ZN(n495) );
  XNOR2_X1 U429 ( .A(n504), .B(n391), .ZN(n382) );
  NAND2_X1 U430 ( .A1(n388), .A2(G224), .ZN(n387) );
  XOR2_X1 U431 ( .A(n404), .B(KEYINPUT4), .Z(n403) );
  XNOR2_X1 U432 ( .A(n435), .B(KEYINPUT67), .ZN(n541) );
  XNOR2_X1 U433 ( .A(n507), .B(n506), .ZN(n394) );
  XNOR2_X1 U434 ( .A(G140), .B(KEYINPUT10), .ZN(n395) );
  XNOR2_X1 U435 ( .A(G122), .B(G116), .ZN(n532) );
  XNOR2_X1 U436 ( .A(G128), .B(G143), .ZN(n392) );
  XNOR2_X1 U437 ( .A(G101), .B(KEYINPUT73), .ZN(n469) );
  XNOR2_X1 U438 ( .A(G128), .B(G143), .ZN(n391) );
  NAND2_X1 U439 ( .A1(n357), .A2(n686), .ZN(n356) );
  NAND2_X1 U440 ( .A1(n358), .A2(n363), .ZN(n357) );
  INV_X1 U441 ( .A(n776), .ZN(n358) );
  NAND2_X1 U442 ( .A1(n362), .A2(n360), .ZN(n359) );
  NAND2_X1 U443 ( .A1(n361), .A2(n777), .ZN(n360) );
  AND2_X1 U444 ( .A1(n776), .A2(n617), .ZN(n361) );
  INV_X1 U445 ( .A(n617), .ZN(n363) );
  INV_X1 U446 ( .A(n777), .ZN(n364) );
  XNOR2_X2 U447 ( .A(n616), .B(KEYINPUT40), .ZN(n777) );
  AND2_X1 U448 ( .A1(n365), .A2(n599), .ZN(n602) );
  NAND2_X1 U449 ( .A1(n369), .A2(n366), .ZN(n373) );
  INV_X1 U450 ( .A(n709), .ZN(n366) );
  NAND2_X1 U451 ( .A1(n370), .A2(n367), .ZN(n528) );
  NAND2_X1 U452 ( .A1(n567), .A2(KEYINPUT108), .ZN(n372) );
  OR2_X1 U453 ( .A1(n373), .A2(n708), .ZN(n715) );
  XNOR2_X1 U454 ( .A(n374), .B(KEYINPUT34), .ZN(n551) );
  NAND2_X1 U455 ( .A1(n375), .A2(n378), .ZN(n692) );
  XNOR2_X2 U456 ( .A(n490), .B(n489), .ZN(n564) );
  NAND2_X1 U457 ( .A1(n528), .A2(n381), .ZN(n376) );
  NAND2_X1 U458 ( .A1(n618), .A2(n381), .ZN(n377) );
  NAND2_X1 U459 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U460 ( .A(n618), .ZN(n379) );
  NOR2_X1 U461 ( .A1(n528), .A2(n381), .ZN(n380) );
  INV_X1 U462 ( .A(KEYINPUT33), .ZN(n381) );
  XNOR2_X2 U463 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n389) );
  XNOR2_X2 U464 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n390) );
  INV_X1 U465 ( .A(n674), .ZN(n607) );
  NAND2_X1 U466 ( .A1(n399), .A2(KEYINPUT47), .ZN(n398) );
  NAND2_X1 U467 ( .A1(n683), .A2(n671), .ZN(n557) );
  OR2_X1 U468 ( .A1(n554), .A2(n414), .ZN(n671) );
  XOR2_X2 U469 ( .A(KEYINPUT87), .B(G110), .Z(n470) );
  XNOR2_X2 U470 ( .A(n756), .B(KEYINPUT68), .ZN(n494) );
  XNOR2_X2 U471 ( .A(n472), .B(n471), .ZN(n756) );
  XNOR2_X2 U472 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X2 U473 ( .A(n419), .B(KEYINPUT1), .ZN(n567) );
  NAND2_X1 U474 ( .A1(n437), .A2(n436), .ZN(n406) );
  NAND2_X1 U475 ( .A1(n437), .A2(n436), .ZN(n621) );
  XNOR2_X1 U476 ( .A(n478), .B(n477), .ZN(n407) );
  XNOR2_X1 U477 ( .A(n478), .B(n477), .ZN(n600) );
  XNOR2_X1 U478 ( .A(n406), .B(n481), .ZN(n408) );
  XNOR2_X1 U479 ( .A(n621), .B(n481), .ZN(n591) );
  BUF_X1 U480 ( .A(n419), .Z(n409) );
  NAND2_X1 U481 ( .A1(n531), .A2(n541), .ZN(n412) );
  NAND2_X1 U482 ( .A1(n410), .A2(n411), .ZN(n413) );
  INV_X1 U483 ( .A(n531), .ZN(n410) );
  INV_X1 U484 ( .A(n541), .ZN(n411) );
  OR2_X1 U485 ( .A1(n593), .A2(n415), .ZN(n414) );
  INV_X1 U486 ( .A(n596), .ZN(n415) );
  INV_X1 U487 ( .A(G131), .ZN(n435) );
  INV_X1 U488 ( .A(G113), .ZN(n465) );
  XNOR2_X1 U489 ( .A(KEYINPUT3), .B(G119), .ZN(n466) );
  NOR2_X1 U490 ( .A1(G237), .A2(G953), .ZN(n516) );
  XNOR2_X1 U491 ( .A(n699), .B(KEYINPUT79), .ZN(n604) );
  NAND2_X1 U492 ( .A1(n655), .A2(n578), .ZN(n579) );
  INV_X1 U493 ( .A(KEYINPUT80), .ZN(n462) );
  AND2_X1 U494 ( .A1(n455), .A2(n454), .ZN(n453) );
  XNOR2_X1 U495 ( .A(n541), .B(n433), .ZN(n432) );
  INV_X1 U496 ( .A(G122), .ZN(n434) );
  XNOR2_X1 U497 ( .A(G113), .B(G104), .ZN(n542) );
  NOR2_X1 U498 ( .A1(n480), .A2(KEYINPUT83), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n523), .B(n522), .ZN(n660) );
  XOR2_X1 U500 ( .A(G107), .B(G104), .Z(n471) );
  INV_X1 U501 ( .A(KEYINPUT28), .ZN(n425) );
  XNOR2_X1 U502 ( .A(n445), .B(n612), .ZN(n724) );
  INV_X1 U503 ( .A(n698), .ZN(n446) );
  BUF_X1 U504 ( .A(n567), .Z(n710) );
  INV_X1 U505 ( .A(KEYINPUT81), .ZN(n464) );
  NAND2_X1 U506 ( .A1(n480), .A2(KEYINPUT83), .ZN(n440) );
  XNOR2_X1 U507 ( .A(G116), .B(G101), .ZN(n519) );
  INV_X1 U508 ( .A(KEYINPUT45), .ZN(n460) );
  INV_X1 U509 ( .A(KEYINPUT19), .ZN(n481) );
  XNOR2_X1 U510 ( .A(KEYINPUT70), .B(KEYINPUT16), .ZN(n467) );
  XNOR2_X1 U511 ( .A(n509), .B(n508), .ZN(n510) );
  INV_X1 U512 ( .A(KEYINPUT93), .ZN(n508) );
  XNOR2_X1 U513 ( .A(G128), .B(G110), .ZN(n509) );
  XNOR2_X1 U514 ( .A(n544), .B(n432), .ZN(n547) );
  XNOR2_X1 U515 ( .A(n523), .B(n497), .ZN(n734) );
  XNOR2_X1 U516 ( .A(n660), .B(n659), .ZN(n661) );
  INV_X1 U517 ( .A(KEYINPUT126), .ZN(n427) );
  XNOR2_X1 U518 ( .A(n645), .B(KEYINPUT59), .ZN(n646) );
  INV_X1 U519 ( .A(n611), .ZN(n444) );
  NAND2_X1 U520 ( .A1(n560), .A2(n431), .ZN(n430) );
  NAND2_X1 U521 ( .A1(n568), .A2(n442), .ZN(n569) );
  AND2_X1 U522 ( .A1(n417), .A2(n710), .ZN(n442) );
  XNOR2_X1 U523 ( .A(n743), .B(n742), .ZN(n422) );
  INV_X1 U524 ( .A(KEYINPUT56), .ZN(n463) );
  XNOR2_X1 U525 ( .A(n578), .B(n418), .ZN(G21) );
  XOR2_X1 U526 ( .A(n657), .B(n658), .Z(n416) );
  AND2_X1 U527 ( .A1(n618), .A2(n704), .ZN(n417) );
  XOR2_X1 U528 ( .A(G119), .B(KEYINPUT127), .Z(n418) );
  NOR2_X1 U529 ( .A1(n590), .A2(n409), .ZN(n611) );
  XNOR2_X2 U530 ( .A(n498), .B(G469), .ZN(n419) );
  NAND2_X1 U531 ( .A1(n739), .A2(G210), .ZN(n452) );
  XNOR2_X1 U532 ( .A(G143), .B(n434), .ZN(n433) );
  NOR2_X1 U533 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U534 ( .A1(n451), .A2(n663), .ZN(n450) );
  XNOR2_X1 U535 ( .A(n452), .B(n416), .ZN(n451) );
  NAND2_X1 U536 ( .A1(n751), .A2(n638), .ZN(n420) );
  NAND2_X1 U537 ( .A1(n750), .A2(n638), .ZN(n690) );
  NAND2_X1 U538 ( .A1(n421), .A2(n355), .ZN(n625) );
  NOR2_X1 U539 ( .A1(n422), .A2(n748), .ZN(G63) );
  OR2_X1 U540 ( .A1(n708), .A2(n480), .ZN(n594) );
  XNOR2_X1 U541 ( .A(n552), .B(KEYINPUT35), .ZN(n580) );
  XNOR2_X1 U542 ( .A(n423), .B(n757), .ZN(n473) );
  NAND2_X1 U543 ( .A1(n424), .A2(n596), .ZN(n597) );
  XNOR2_X1 U544 ( .A(n594), .B(n595), .ZN(n424) );
  XNOR2_X1 U545 ( .A(n625), .B(KEYINPUT48), .ZN(n633) );
  XNOR2_X1 U546 ( .A(n589), .B(n425), .ZN(n590) );
  XNOR2_X2 U547 ( .A(n426), .B(n460), .ZN(n642) );
  NAND2_X1 U548 ( .A1(n448), .A2(n458), .ZN(n426) );
  NOR2_X2 U549 ( .A1(G902), .A2(n734), .ZN(n498) );
  NOR2_X2 U550 ( .A1(n642), .A2(n428), .ZN(n643) );
  XNOR2_X1 U551 ( .A(n428), .B(n427), .ZN(n766) );
  INV_X1 U552 ( .A(n559), .ZN(n431) );
  NAND2_X1 U553 ( .A1(n439), .A2(n438), .ZN(n436) );
  AND2_X2 U554 ( .A1(n441), .A2(n440), .ZN(n437) );
  INV_X1 U555 ( .A(n407), .ZN(n439) );
  NAND2_X1 U556 ( .A1(n600), .A2(KEYINPUT83), .ZN(n441) );
  NAND2_X1 U557 ( .A1(n568), .A2(n710), .ZN(n443) );
  XNOR2_X1 U558 ( .A(n443), .B(KEYINPUT107), .ZN(n572) );
  INV_X1 U559 ( .A(n601), .ZN(n631) );
  NAND2_X1 U560 ( .A1(n447), .A2(n446), .ZN(n445) );
  INV_X1 U561 ( .A(n697), .ZN(n447) );
  XNOR2_X1 U562 ( .A(n449), .B(n462), .ZN(n448) );
  NAND2_X1 U563 ( .A1(n456), .A2(n453), .ZN(n449) );
  XNOR2_X1 U564 ( .A(n450), .B(n463), .ZN(G51) );
  XNOR2_X1 U565 ( .A(n558), .B(KEYINPUT102), .ZN(n454) );
  INV_X1 U566 ( .A(n774), .ZN(n455) );
  XNOR2_X1 U567 ( .A(n457), .B(n464), .ZN(n456) );
  NAND2_X1 U568 ( .A1(n580), .A2(KEYINPUT44), .ZN(n457) );
  NAND2_X1 U569 ( .A1(n459), .A2(n461), .ZN(n458) );
  NAND2_X1 U570 ( .A1(n584), .A2(n583), .ZN(n461) );
  BUF_X1 U571 ( .A(n739), .Z(n744) );
  XNOR2_X1 U572 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U573 ( .A(n741), .B(n740), .ZN(n742) );
  INV_X1 U574 ( .A(n655), .ZN(n656) );
  XNOR2_X1 U575 ( .A(n466), .B(n465), .ZN(n517) );
  XNOR2_X1 U576 ( .A(n532), .B(n467), .ZN(n468) );
  XNOR2_X1 U577 ( .A(n517), .B(n468), .ZN(n757) );
  XNOR2_X1 U578 ( .A(n494), .B(n473), .ZN(n657) );
  XNOR2_X1 U579 ( .A(G902), .B(KEYINPUT15), .ZN(n639) );
  NAND2_X1 U580 ( .A1(n657), .A2(n639), .ZN(n478) );
  INV_X1 U581 ( .A(G902), .ZN(n524) );
  INV_X1 U582 ( .A(G237), .ZN(n474) );
  NAND2_X1 U583 ( .A1(n524), .A2(n474), .ZN(n479) );
  NAND2_X1 U584 ( .A1(n479), .A2(G210), .ZN(n476) );
  INV_X1 U585 ( .A(KEYINPUT89), .ZN(n475) );
  NAND2_X1 U586 ( .A1(n479), .A2(G214), .ZN(n694) );
  INV_X1 U587 ( .A(n694), .ZN(n480) );
  NAND2_X1 U588 ( .A1(G234), .A2(G237), .ZN(n482) );
  XNOR2_X1 U589 ( .A(n482), .B(KEYINPUT14), .ZN(n483) );
  XNOR2_X1 U590 ( .A(KEYINPUT72), .B(n483), .ZN(n486) );
  AND2_X1 U591 ( .A1(n486), .A2(G953), .ZN(n484) );
  NAND2_X1 U592 ( .A1(G902), .A2(n484), .ZN(n585) );
  NOR2_X1 U593 ( .A1(G898), .A2(n585), .ZN(n485) );
  XNOR2_X1 U594 ( .A(n485), .B(KEYINPUT90), .ZN(n487) );
  NAND2_X1 U595 ( .A1(G952), .A2(n486), .ZN(n723) );
  NOR2_X1 U596 ( .A1(n723), .A2(G953), .ZN(n587) );
  OR2_X1 U597 ( .A1(n487), .A2(n587), .ZN(n488) );
  NAND2_X1 U598 ( .A1(n591), .A2(n488), .ZN(n490) );
  INV_X1 U599 ( .A(KEYINPUT0), .ZN(n489) );
  XOR2_X1 U600 ( .A(G140), .B(KEYINPUT92), .Z(n492) );
  NAND2_X1 U601 ( .A1(G227), .A2(n405), .ZN(n491) );
  XNOR2_X1 U602 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U603 ( .A(n494), .B(n493), .ZN(n497) );
  XNOR2_X2 U604 ( .A(n764), .B(G146), .ZN(n523) );
  NAND2_X1 U605 ( .A1(n639), .A2(G234), .ZN(n500) );
  XNOR2_X1 U606 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n499) );
  XNOR2_X1 U607 ( .A(n500), .B(n499), .ZN(n512) );
  NAND2_X1 U608 ( .A1(n512), .A2(G221), .ZN(n503) );
  INV_X1 U609 ( .A(KEYINPUT95), .ZN(n501) );
  XNOR2_X1 U610 ( .A(n501), .B(KEYINPUT21), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n503), .B(n502), .ZN(n563) );
  INV_X1 U612 ( .A(n563), .ZN(n705) );
  NAND2_X1 U613 ( .A1(G234), .A2(n405), .ZN(n505) );
  XOR2_X1 U614 ( .A(KEYINPUT8), .B(n505), .Z(n537) );
  NAND2_X1 U615 ( .A1(n537), .A2(G221), .ZN(n511) );
  XOR2_X1 U616 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n507) );
  XNOR2_X1 U617 ( .A(G119), .B(G137), .ZN(n506) );
  NOR2_X1 U618 ( .A1(G902), .A2(n745), .ZN(n515) );
  NAND2_X1 U619 ( .A1(G217), .A2(n512), .ZN(n513) );
  XNOR2_X1 U620 ( .A(n513), .B(KEYINPUT25), .ZN(n514) );
  XNOR2_X2 U621 ( .A(n515), .B(n514), .ZN(n704) );
  NAND2_X1 U622 ( .A1(n705), .A2(n704), .ZN(n709) );
  XNOR2_X1 U623 ( .A(n516), .B(KEYINPUT74), .ZN(n545) );
  NAND2_X1 U624 ( .A1(n545), .A2(G210), .ZN(n518) );
  XNOR2_X1 U625 ( .A(n518), .B(n517), .ZN(n521) );
  XNOR2_X1 U626 ( .A(n519), .B(KEYINPUT5), .ZN(n520) );
  NAND2_X1 U627 ( .A1(n660), .A2(n524), .ZN(n526) );
  INV_X1 U628 ( .A(G472), .ZN(n525) );
  XNOR2_X2 U629 ( .A(n526), .B(n525), .ZN(n708) );
  INV_X1 U630 ( .A(n708), .ZN(n593) );
  XOR2_X1 U631 ( .A(KEYINPUT6), .B(KEYINPUT103), .Z(n527) );
  XNOR2_X1 U632 ( .A(n593), .B(n527), .ZN(n618) );
  XOR2_X1 U633 ( .A(KEYINPUT98), .B(KEYINPUT9), .Z(n530) );
  XNOR2_X1 U634 ( .A(KEYINPUT97), .B(KEYINPUT99), .ZN(n529) );
  XNOR2_X1 U635 ( .A(n530), .B(n529), .ZN(n536) );
  XNOR2_X1 U636 ( .A(n531), .B(G107), .ZN(n534) );
  XNOR2_X1 U637 ( .A(n532), .B(KEYINPUT7), .ZN(n533) );
  XNOR2_X1 U638 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U639 ( .A(n536), .B(n535), .Z(n539) );
  NAND2_X1 U640 ( .A1(G217), .A2(n537), .ZN(n538) );
  XNOR2_X1 U641 ( .A(n539), .B(n538), .ZN(n741) );
  NOR2_X1 U642 ( .A1(n741), .A2(G902), .ZN(n540) );
  XOR2_X1 U643 ( .A(n540), .B(G478), .Z(n560) );
  XOR2_X1 U644 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n543) );
  XNOR2_X1 U645 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U646 ( .A1(G214), .A2(n545), .ZN(n546) );
  XNOR2_X1 U647 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U648 ( .A(n763), .B(n548), .ZN(n645) );
  NOR2_X1 U649 ( .A1(G902), .A2(n645), .ZN(n550) );
  XNOR2_X1 U650 ( .A(KEYINPUT13), .B(G475), .ZN(n549) );
  XNOR2_X1 U651 ( .A(n550), .B(n549), .ZN(n559) );
  AND2_X1 U652 ( .A1(n560), .A2(n559), .ZN(n599) );
  NAND2_X1 U653 ( .A1(n551), .A2(n599), .ZN(n552) );
  BUF_X1 U654 ( .A(n564), .Z(n553) );
  NAND2_X1 U655 ( .A1(n557), .A2(n604), .ZN(n558) );
  NOR2_X1 U656 ( .A1(n560), .A2(n559), .ZN(n562) );
  INV_X1 U657 ( .A(KEYINPUT104), .ZN(n561) );
  XNOR2_X1 U658 ( .A(n562), .B(n561), .ZN(n697) );
  NOR2_X1 U659 ( .A1(n697), .A2(n563), .ZN(n565) );
  NAND2_X1 U660 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U661 ( .A(n566), .B(KEYINPUT22), .ZN(n576) );
  INV_X1 U662 ( .A(n576), .ZN(n568) );
  INV_X1 U663 ( .A(n704), .ZN(n570) );
  AND2_X1 U664 ( .A1(n708), .A2(n570), .ZN(n571) );
  NAND2_X1 U665 ( .A1(n572), .A2(n571), .ZN(n655) );
  NOR2_X1 U666 ( .A1(n710), .A2(n704), .ZN(n573) );
  XNOR2_X1 U667 ( .A(n573), .B(KEYINPUT106), .ZN(n574) );
  NAND2_X1 U668 ( .A1(n574), .A2(n618), .ZN(n575) );
  OR2_X1 U669 ( .A1(n576), .A2(n575), .ZN(n577) );
  BUF_X1 U670 ( .A(n580), .Z(n773) );
  OR2_X1 U671 ( .A1(n773), .A2(KEYINPUT44), .ZN(n581) );
  INV_X1 U672 ( .A(KEYINPUT44), .ZN(n583) );
  INV_X1 U673 ( .A(n642), .ZN(n750) );
  NOR2_X1 U674 ( .A1(G900), .A2(n585), .ZN(n586) );
  NOR2_X1 U675 ( .A1(n587), .A2(n586), .ZN(n598) );
  NOR2_X1 U676 ( .A1(n598), .A2(n704), .ZN(n588) );
  NAND2_X1 U677 ( .A1(n588), .A2(n705), .ZN(n619) );
  NOR2_X1 U678 ( .A1(n708), .A2(n619), .ZN(n589) );
  NAND2_X1 U679 ( .A1(n611), .A2(n408), .ZN(n592) );
  XOR2_X1 U680 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n595) );
  BUF_X1 U681 ( .A(n407), .Z(n601) );
  NAND2_X1 U682 ( .A1(n602), .A2(n631), .ZN(n654) );
  XNOR2_X1 U683 ( .A(n603), .B(KEYINPUT78), .ZN(n609) );
  XNOR2_X1 U684 ( .A(KEYINPUT65), .B(KEYINPUT47), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n695), .A2(n694), .ZN(n698) );
  XNOR2_X1 U688 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n613), .B(KEYINPUT42), .ZN(n776) );
  XNOR2_X1 U690 ( .A(KEYINPUT69), .B(KEYINPUT39), .ZN(n614) );
  XNOR2_X1 U691 ( .A(n615), .B(n614), .ZN(n634) );
  NAND2_X1 U692 ( .A1(n634), .A2(n429), .ZN(n616) );
  XOR2_X1 U693 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n617) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n620), .A2(n429), .ZN(n626) );
  INV_X1 U696 ( .A(n406), .ZN(n622) );
  NOR2_X1 U697 ( .A1(n626), .A2(n622), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(KEYINPUT36), .ZN(n624) );
  INV_X1 U699 ( .A(n710), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n624), .A2(n627), .ZN(n686) );
  XOR2_X1 U701 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n630) );
  NOR2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n628), .A2(n694), .ZN(n629) );
  XOR2_X1 U704 ( .A(n630), .B(n629), .Z(n632) );
  NOR2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n653) );
  NOR2_X2 U706 ( .A1(n633), .A2(n653), .ZN(n641) );
  NAND2_X1 U707 ( .A1(n634), .A2(n675), .ZN(n688) );
  NAND2_X1 U708 ( .A1(n688), .A2(KEYINPUT2), .ZN(n636) );
  INV_X1 U709 ( .A(KEYINPUT76), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(n637) );
  AND2_X1 U711 ( .A1(n641), .A2(n637), .ZN(n638) );
  INV_X1 U712 ( .A(n639), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n690), .A2(n640), .ZN(n644) );
  NOR2_X2 U714 ( .A1(n643), .A2(KEYINPUT2), .ZN(n689) );
  NOR2_X4 U715 ( .A1(n644), .A2(n689), .ZN(n739) );
  NAND2_X1 U716 ( .A1(n739), .A2(G475), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(n650) );
  INV_X1 U718 ( .A(G952), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n648), .A2(G953), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n649), .B(KEYINPUT86), .ZN(n663) );
  NAND2_X1 U721 ( .A1(n650), .A2(n663), .ZN(n652) );
  INV_X1 U722 ( .A(KEYINPUT60), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(G60) );
  XOR2_X1 U724 ( .A(n653), .B(G140), .Z(G42) );
  XNOR2_X1 U725 ( .A(n654), .B(G143), .ZN(G45) );
  XOR2_X1 U726 ( .A(n656), .B(G110), .Z(G12) );
  XNOR2_X1 U727 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n658) );
  INV_X1 U728 ( .A(n663), .ZN(n748) );
  NAND2_X1 U729 ( .A1(n739), .A2(G472), .ZN(n662) );
  XNOR2_X1 U730 ( .A(KEYINPUT84), .B(KEYINPUT62), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n662), .B(n661), .ZN(n664) );
  NAND2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n667) );
  XNOR2_X1 U733 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n665) );
  XOR2_X1 U734 ( .A(n665), .B(KEYINPUT85), .Z(n666) );
  XNOR2_X1 U735 ( .A(n667), .B(n666), .ZN(G57) );
  NOR2_X1 U736 ( .A1(n680), .A2(n671), .ZN(n668) );
  XOR2_X1 U737 ( .A(G104), .B(n668), .Z(G6) );
  XOR2_X1 U738 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n670) );
  XNOR2_X1 U739 ( .A(G107), .B(KEYINPUT114), .ZN(n669) );
  XNOR2_X1 U740 ( .A(n670), .B(n669), .ZN(n673) );
  INV_X1 U741 ( .A(n675), .ZN(n682) );
  NOR2_X1 U742 ( .A1(n682), .A2(n671), .ZN(n672) );
  XOR2_X1 U743 ( .A(n673), .B(n672), .Z(G9) );
  XOR2_X1 U744 ( .A(G128), .B(KEYINPUT29), .Z(n677) );
  NAND2_X1 U745 ( .A1(n674), .A2(n675), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n677), .B(n676), .ZN(G30) );
  XOR2_X1 U747 ( .A(G146), .B(KEYINPUT115), .Z(n679) );
  NAND2_X1 U748 ( .A1(n674), .A2(n429), .ZN(n678) );
  XNOR2_X1 U749 ( .A(n679), .B(n678), .ZN(G48) );
  NOR2_X1 U750 ( .A1(n680), .A2(n683), .ZN(n681) );
  XOR2_X1 U751 ( .A(G113), .B(n681), .Z(G15) );
  NOR2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U753 ( .A(G116), .B(n684), .Z(G18) );
  XOR2_X1 U754 ( .A(KEYINPUT116), .B(KEYINPUT37), .Z(n685) );
  XNOR2_X1 U755 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U756 ( .A(G125), .B(n687), .ZN(G27) );
  XNOR2_X1 U757 ( .A(G134), .B(n688), .ZN(G36) );
  XNOR2_X1 U758 ( .A(n689), .B(KEYINPUT77), .ZN(n691) );
  NAND2_X1 U759 ( .A1(n691), .A2(n420), .ZN(n729) );
  BUF_X1 U760 ( .A(n692), .Z(n693) );
  NOR2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n701) );
  NOR2_X1 U763 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U765 ( .A(n702), .B(KEYINPUT118), .ZN(n703) );
  NOR2_X1 U766 ( .A1(n693), .A2(n703), .ZN(n720) );
  NOR2_X1 U767 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U768 ( .A(n706), .B(KEYINPUT49), .ZN(n707) );
  NAND2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n713) );
  NAND2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U771 ( .A(KEYINPUT50), .B(n711), .Z(n712) );
  NOR2_X1 U772 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U773 ( .A(n714), .B(KEYINPUT117), .ZN(n716) );
  NAND2_X1 U774 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U775 ( .A(KEYINPUT51), .B(n717), .ZN(n718) );
  NOR2_X1 U776 ( .A1(n724), .A2(n718), .ZN(n719) );
  NOR2_X1 U777 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U778 ( .A(n721), .B(KEYINPUT52), .ZN(n722) );
  NOR2_X1 U779 ( .A1(n723), .A2(n722), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n724), .A2(n693), .ZN(n725) );
  XOR2_X1 U781 ( .A(KEYINPUT119), .B(n725), .Z(n726) );
  NOR2_X1 U782 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U783 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U784 ( .A1(n730), .A2(G953), .ZN(n731) );
  XNOR2_X1 U785 ( .A(n731), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U786 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n733) );
  XNOR2_X1 U787 ( .A(KEYINPUT121), .B(KEYINPUT120), .ZN(n732) );
  XNOR2_X1 U788 ( .A(n733), .B(n732), .ZN(n735) );
  XNOR2_X1 U789 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U790 ( .A1(n739), .A2(G469), .ZN(n736) );
  XOR2_X1 U791 ( .A(n737), .B(n736), .Z(n738) );
  NOR2_X1 U792 ( .A1(n748), .A2(n738), .ZN(G54) );
  NAND2_X1 U793 ( .A1(n744), .A2(G478), .ZN(n743) );
  XOR2_X1 U794 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n740) );
  NAND2_X1 U795 ( .A1(n744), .A2(G217), .ZN(n747) );
  XNOR2_X1 U796 ( .A(n745), .B(KEYINPUT124), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n747), .B(n746), .ZN(n749) );
  NOR2_X1 U798 ( .A1(n749), .A2(n748), .ZN(G66) );
  BUF_X1 U799 ( .A(n750), .Z(n751) );
  NAND2_X1 U800 ( .A1(n751), .A2(n405), .ZN(n755) );
  NAND2_X1 U801 ( .A1(G953), .A2(G224), .ZN(n752) );
  XNOR2_X1 U802 ( .A(KEYINPUT61), .B(n752), .ZN(n753) );
  NAND2_X1 U803 ( .A1(n753), .A2(G898), .ZN(n754) );
  NAND2_X1 U804 ( .A1(n755), .A2(n754), .ZN(n761) );
  XOR2_X1 U805 ( .A(n757), .B(n756), .Z(n759) );
  NOR2_X1 U806 ( .A1(G898), .A2(n405), .ZN(n758) );
  NOR2_X1 U807 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U808 ( .A(n761), .B(n760), .ZN(n762) );
  XOR2_X1 U809 ( .A(KEYINPUT125), .B(n762), .Z(G69) );
  XOR2_X1 U810 ( .A(n764), .B(n763), .Z(n768) );
  INV_X1 U811 ( .A(n768), .ZN(n765) );
  XOR2_X1 U812 ( .A(n766), .B(n765), .Z(n767) );
  NAND2_X1 U813 ( .A1(n767), .A2(n405), .ZN(n772) );
  XOR2_X1 U814 ( .A(G227), .B(n768), .Z(n769) );
  NAND2_X1 U815 ( .A1(n769), .A2(G900), .ZN(n770) );
  NAND2_X1 U816 ( .A1(n770), .A2(G953), .ZN(n771) );
  NAND2_X1 U817 ( .A1(n772), .A2(n771), .ZN(G72) );
  XOR2_X1 U818 ( .A(n773), .B(G122), .Z(G24) );
  XNOR2_X1 U819 ( .A(G101), .B(n774), .ZN(n775) );
  XNOR2_X1 U820 ( .A(n775), .B(KEYINPUT113), .ZN(G3) );
  XNOR2_X1 U821 ( .A(G137), .B(n776), .ZN(G39) );
  XNOR2_X1 U822 ( .A(G131), .B(n777), .ZN(G33) );
endmodule

