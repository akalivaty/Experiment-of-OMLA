//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(new_n190), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(G237), .A2(G953), .ZN(new_n197));
  AOI21_X1  g011(.A(G143), .B1(new_n197), .B2(G214), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(G143), .A3(G214), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT18), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n199), .B(new_n200), .C1(new_n201), .C2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n200), .ZN(new_n204));
  OAI21_X1  g018(.A(G131), .B1(new_n204), .B2(new_n198), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n196), .B(new_n203), .C1(new_n201), .C2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n199), .A2(new_n202), .A3(new_n200), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n209));
  OR3_X1    g023(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n191), .A2(KEYINPUT91), .A3(KEYINPUT19), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT19), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT91), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n194), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(G146), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n206), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G113), .B(G122), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n219), .B(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n205), .A2(new_n207), .A3(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n209), .A2(G146), .A3(new_n210), .ZN(new_n226));
  AOI21_X1  g040(.A(G146), .B1(new_n209), .B2(new_n210), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n225), .B(new_n228), .C1(new_n224), .C2(new_n205), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n221), .A3(new_n206), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G475), .ZN(new_n232));
  INV_X1    g046(.A(G902), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  XOR2_X1   g048(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT92), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(KEYINPUT92), .A3(new_n235), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n234), .A2(KEYINPUT20), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n229), .A2(new_n206), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n222), .ZN(new_n243));
  AOI21_X1  g057(.A(G902), .B1(new_n243), .B2(new_n230), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT93), .B(G475), .ZN(new_n245));
  OR2_X1    g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT94), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT94), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n241), .A2(new_n249), .A3(new_n246), .ZN(new_n250));
  INV_X1    g064(.A(G953), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n251), .A2(G952), .ZN(new_n252));
  INV_X1    g066(.A(G234), .ZN(new_n253));
  INV_X1    g067(.A(G237), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(G902), .B(G953), .C1(new_n253), .C2(new_n254), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT96), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT21), .B(G898), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(G143), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G116), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT14), .A3(G122), .ZN(new_n270));
  XNOR2_X1  g084(.A(G116), .B(G122), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(G107), .B(new_n270), .C1(new_n272), .C2(KEYINPUT14), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n268), .B(new_n273), .C1(G107), .C2(new_n272), .ZN(new_n274));
  INV_X1    g088(.A(G143), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT13), .A3(G128), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n276), .B(KEYINPUT95), .Z(new_n277));
  OAI21_X1  g091(.A(new_n265), .B1(new_n263), .B2(KEYINPUT13), .ZN(new_n278));
  OAI21_X1  g092(.A(G134), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n266), .A2(new_n267), .ZN(new_n280));
  INV_X1    g094(.A(G107), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n271), .B(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(KEYINPUT9), .B(G234), .Z(new_n285));
  AND3_X1   g099(.A1(new_n285), .A2(G217), .A3(new_n251), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n284), .B(new_n286), .Z(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n233), .ZN(new_n288));
  INV_X1    g102(.A(G478), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(KEYINPUT15), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n284), .B(new_n286), .ZN(new_n292));
  OR3_X1    g106(.A1(new_n292), .A2(G902), .A3(new_n290), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n248), .A2(new_n250), .A3(new_n261), .A4(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G469), .ZN(new_n297));
  XNOR2_X1  g111(.A(G110), .B(G140), .ZN(new_n298));
  INV_X1    g112(.A(G227), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(G953), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n298), .B(new_n300), .Z(new_n301));
  INV_X1    g115(.A(KEYINPUT10), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT1), .B1(new_n275), .B2(G146), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n262), .B1(new_n303), .B2(KEYINPUT66), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n192), .A2(G143), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT1), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n275), .A2(G146), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G143), .B(G146), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(G128), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n302), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT82), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n281), .A2(G104), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n281), .A2(G104), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(KEYINPUT3), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G101), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n281), .A3(G104), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n319), .A2(KEYINPUT81), .A3(new_n320), .A4(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT3), .B1(new_n220), .B2(G107), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n220), .A2(G107), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n324), .A2(new_n322), .A3(new_n320), .A4(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n320), .B1(new_n318), .B2(new_n325), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n316), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  AOI211_X1 g146(.A(KEYINPUT82), .B(new_n330), .C1(new_n323), .C2(new_n328), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n315), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT0), .A2(G128), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT64), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(KEYINPUT0), .B2(G128), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT0), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n262), .A3(KEYINPUT64), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n310), .A2(new_n335), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n312), .A2(KEYINPUT0), .A3(G128), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n324), .A2(new_n322), .A3(new_n325), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G101), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n343), .B1(new_n329), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n343), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n342), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n262), .B1(new_n305), .B2(KEYINPUT1), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n314), .B1(new_n350), .B2(new_n312), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n326), .A2(new_n327), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n326), .A2(new_n327), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n331), .B(new_n351), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n302), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n334), .A2(new_n349), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT65), .ZN(new_n357));
  INV_X1    g171(.A(G137), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(G134), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n267), .A2(KEYINPUT65), .A3(G137), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT11), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n267), .B2(G137), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n358), .A2(KEYINPUT11), .A3(G134), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G131), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n360), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n367), .A2(new_n202), .A3(new_n363), .A4(new_n364), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n356), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n365), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n202), .B1(new_n371), .B2(new_n367), .ZN(new_n372));
  INV_X1    g186(.A(new_n368), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n334), .A2(new_n349), .A3(new_n374), .A4(new_n355), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n301), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n301), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n311), .A2(new_n314), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n330), .B1(new_n323), .B2(new_n328), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n354), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT12), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT83), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(new_n374), .B2(new_n382), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n380), .A2(new_n383), .A3(new_n369), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n383), .B1(new_n380), .B2(new_n369), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n297), .B(new_n233), .C1(new_n376), .C2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n301), .ZN(new_n390));
  INV_X1    g204(.A(new_n375), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n390), .B1(new_n391), .B2(new_n386), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n370), .A2(new_n375), .A3(new_n301), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(G469), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(G469), .A2(G902), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n285), .ZN(new_n398));
  OAI21_X1  g212(.A(G221), .B1(new_n398), .B2(G902), .ZN(new_n399));
  XOR2_X1   g213(.A(new_n399), .B(KEYINPUT79), .Z(new_n400));
  XOR2_X1   g214(.A(new_n400), .B(KEYINPUT80), .Z(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT84), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n404), .B(new_n401), .C1(new_n389), .C2(new_n396), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n296), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT32), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n342), .B1(new_n373), .B2(new_n372), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT68), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT68), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n369), .A2(new_n410), .A3(new_n342), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n267), .A2(G137), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n358), .A2(G134), .ZN(new_n414));
  OAI21_X1  g228(.A(G131), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n368), .A2(KEYINPUT69), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT69), .B1(new_n368), .B2(new_n415), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n378), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT70), .ZN(new_n419));
  XNOR2_X1  g233(.A(G116), .B(G119), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT2), .B(G113), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n422), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT70), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n378), .B(new_n427), .C1(new_n416), .C2(new_n417), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n412), .A2(new_n419), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n197), .A2(G210), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(new_n320), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n431), .B(new_n432), .Z(new_n433));
  NAND4_X1  g247(.A1(new_n412), .A2(new_n419), .A3(KEYINPUT30), .A4(new_n428), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n312), .B1(new_n304), .B2(new_n307), .ZN(new_n436));
  INV_X1    g250(.A(new_n314), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n368), .B(new_n415), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n408), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT30), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT67), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT67), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n442), .B(KEYINPUT30), .C1(new_n408), .C2(new_n438), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n425), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n429), .B(new_n433), .C1(new_n435), .C2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT31), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n368), .A2(new_n415), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n378), .A2(new_n448), .B1(new_n369), .B2(new_n342), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n442), .B1(new_n449), .B2(KEYINPUT30), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n439), .A2(KEYINPUT67), .A3(new_n440), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n434), .A3(new_n425), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n453), .A2(KEYINPUT31), .A3(new_n429), .A4(new_n433), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n439), .A2(new_n425), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n429), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT28), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n418), .A2(new_n408), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT28), .B1(new_n458), .B2(new_n426), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n433), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n447), .A2(new_n454), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(G472), .A2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n407), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n462), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n426), .B1(new_n450), .B2(new_n451), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n412), .A2(new_n419), .A3(new_n428), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n468), .A2(new_n434), .B1(new_n469), .B2(new_n426), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT31), .B1(new_n470), .B2(new_n433), .ZN(new_n471));
  AND4_X1   g285(.A1(KEYINPUT31), .A2(new_n453), .A3(new_n429), .A4(new_n433), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(KEYINPUT32), .A3(new_n464), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n466), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G472), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT29), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT71), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n457), .A2(new_n478), .A3(new_n460), .A4(new_n433), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n453), .A2(new_n429), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT71), .B1(new_n480), .B2(new_n462), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n462), .B(new_n459), .C1(new_n456), .C2(KEYINPUT28), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n477), .B(new_n479), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT28), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n412), .A2(new_n419), .A3(new_n428), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n425), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n484), .B1(new_n486), .B2(new_n429), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n459), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n462), .A2(new_n477), .ZN(new_n489));
  AOI21_X1  g303(.A(G902), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n476), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n475), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G217), .B1(new_n253), .B2(G902), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n494), .B(KEYINPUT72), .Z(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT22), .B(G137), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n251), .A2(G221), .A3(G234), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT74), .ZN(new_n500));
  NAND2_X1  g314(.A1(KEYINPUT24), .A2(G110), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(KEYINPUT24), .A2(G110), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT73), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n262), .B2(G119), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n262), .A2(G119), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OR2_X1    g322(.A1(KEYINPUT24), .A2(G110), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT74), .A3(new_n501), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n262), .A3(G119), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n504), .A2(new_n508), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n262), .A2(KEYINPUT23), .A3(G119), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT23), .ZN(new_n514));
  INV_X1    g328(.A(G119), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n514), .B1(new_n515), .B2(G128), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(G128), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G110), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n512), .B(new_n519), .C1(new_n226), .C2(new_n227), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT75), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n209), .A2(new_n210), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n192), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n211), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT75), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n512), .A4(new_n519), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n504), .A2(new_n510), .B1(new_n508), .B2(new_n511), .ZN(new_n528));
  INV_X1    g342(.A(G110), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n529), .B(new_n513), .C1(new_n516), .C2(new_n517), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n211), .B(new_n193), .C1(new_n528), .C2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT76), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n504), .A2(new_n510), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT73), .B1(new_n515), .B2(G128), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n511), .B1(new_n536), .B2(new_n517), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n530), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n539), .A2(KEYINPUT76), .A3(new_n211), .A4(new_n193), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT77), .B1(new_n527), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n521), .A2(new_n526), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT77), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n534), .A4(new_n540), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n499), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n545), .A2(new_n499), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n546), .A2(new_n547), .A3(G902), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT25), .B1(new_n548), .B2(KEYINPUT78), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n542), .A2(new_n545), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n498), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n499), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n233), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT25), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n495), .B1(new_n549), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n551), .A2(new_n552), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n494), .A2(new_n233), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G214), .B1(G237), .B2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G210), .B1(G237), .B2(G902), .ZN(new_n564));
  OR3_X1    g378(.A1(new_n378), .A2(KEYINPUT89), .A3(G125), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n340), .A2(new_n341), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G125), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT88), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT89), .B1(new_n378), .B2(G125), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n565), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G224), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G953), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n570), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT5), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n515), .A3(G116), .ZN(new_n575));
  OAI211_X1 g389(.A(G113), .B(new_n575), .C1(new_n421), .C2(new_n574), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n423), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n331), .B1(new_n352), .B2(new_n353), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT82), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n379), .A2(new_n316), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n345), .B1(new_n352), .B2(new_n353), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT4), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n426), .B1(new_n583), .B2(new_n347), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT85), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n323), .A2(new_n328), .B1(G101), .B2(new_n344), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n347), .B1(new_n586), .B2(new_n343), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n425), .ZN(new_n588));
  INV_X1    g402(.A(new_n577), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n332), .B2(new_n333), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT85), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(G110), .B(G122), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT86), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n585), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  OR3_X1    g409(.A1(new_n581), .A2(new_n584), .A3(new_n593), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(KEYINPUT6), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT6), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n585), .A2(new_n598), .A3(new_n592), .A4(new_n594), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT87), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n573), .B(new_n597), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT7), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n570), .B1(new_n604), .B2(new_n572), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n593), .B(KEYINPUT8), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n379), .B(new_n577), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n570), .A2(new_n604), .A3(new_n572), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n610), .B2(new_n596), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n564), .B1(new_n603), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n603), .A2(new_n611), .A3(new_n564), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n563), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n406), .A2(new_n493), .A3(new_n561), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G101), .ZN(G3));
  AND3_X1   g431(.A1(new_n603), .A2(new_n564), .A3(new_n611), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n562), .B(new_n261), .C1(new_n618), .C2(new_n612), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n292), .A2(KEYINPUT33), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n292), .A2(KEYINPUT33), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n289), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n288), .A2(G478), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n289), .A2(new_n233), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n241), .A2(new_n249), .A3(new_n246), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n249), .B1(new_n241), .B2(new_n246), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n619), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n447), .A2(new_n454), .ZN(new_n630));
  AOI21_X1  g444(.A(G902), .B1(new_n630), .B2(new_n467), .ZN(new_n631));
  OAI22_X1  g445(.A1(new_n631), .A2(new_n476), .B1(new_n463), .B2(new_n465), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n403), .B2(new_n405), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n629), .A2(new_n561), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT97), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  OAI211_X1 g451(.A(new_n238), .B(new_n239), .C1(new_n235), .C2(new_n234), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n294), .A2(new_n246), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n619), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(new_n561), .A3(new_n633), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  INV_X1    g457(.A(new_n495), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n548), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n555), .B1(new_n553), .B2(new_n554), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n541), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n543), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n499), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n233), .A3(new_n494), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n647), .A2(KEYINPUT98), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT98), .ZN(new_n654));
  INV_X1    g468(.A(new_n652), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n654), .B1(new_n557), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n632), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n406), .A2(new_n657), .A3(new_n615), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT37), .B(G110), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT99), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n659), .B(new_n661), .ZN(G12));
  NAND2_X1  g476(.A1(new_n403), .A2(new_n405), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n493), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n562), .B1(new_n618), .B2(new_n612), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n653), .A2(new_n656), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT100), .B(G900), .Z(new_n668));
  NAND2_X1  g482(.A1(new_n258), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n255), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n639), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XOR2_X1   g488(.A(new_n670), .B(KEYINPUT39), .Z(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n663), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT40), .Z(new_n678));
  OAI21_X1  g492(.A(new_n294), .B1(new_n626), .B2(new_n627), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n657), .A2(new_n563), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n470), .A2(new_n462), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n486), .A2(new_n429), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n233), .B1(new_n684), .B2(new_n433), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n475), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n618), .A2(new_n612), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT38), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n680), .B2(new_n681), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n678), .A2(new_n682), .A3(new_n687), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  NOR2_X1   g506(.A1(new_n628), .A2(new_n671), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n667), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  OAI21_X1  g509(.A(new_n233), .B1(new_n376), .B2(new_n387), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(KEYINPUT102), .A3(new_n388), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n696), .A2(new_n699), .A3(G469), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n400), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n466), .A2(new_n474), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n701), .B(new_n561), .C1(new_n702), .C2(new_n491), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n629), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n640), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NOR2_X1   g523(.A1(new_n666), .A2(new_n665), .ZN(new_n710));
  INV_X1    g524(.A(new_n400), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n388), .A2(KEYINPUT102), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n579), .A2(new_n580), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n713), .A2(new_n315), .B1(new_n587), .B2(new_n342), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n374), .B1(new_n714), .B2(new_n355), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n390), .B1(new_n715), .B2(new_n391), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n375), .B(new_n301), .C1(new_n384), .C2(new_n385), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n297), .B1(new_n718), .B2(new_n233), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n700), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n711), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n475), .B2(new_n492), .ZN(new_n723));
  INV_X1    g537(.A(new_n296), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n710), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(new_n631), .B2(new_n476), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n684), .A2(KEYINPUT28), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n460), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT103), .B1(new_n487), .B2(new_n459), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n462), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n630), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n464), .ZN(new_n735));
  OAI211_X1 g549(.A(KEYINPUT104), .B(G472), .C1(new_n463), .C2(G902), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n728), .A2(new_n561), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n260), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n665), .A2(new_n722), .A3(new_n679), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  NOR2_X1   g555(.A1(new_n665), .A2(new_n722), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n728), .A2(new_n735), .A3(new_n736), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT105), .B1(new_n743), .B2(new_n657), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n728), .A2(new_n735), .A3(new_n736), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n745), .A2(new_n666), .A3(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n693), .B(new_n742), .C1(new_n744), .C2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  NOR3_X1   g563(.A1(new_n618), .A2(new_n612), .A3(new_n563), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n693), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n397), .A2(new_n400), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n561), .B(new_n753), .C1(new_n702), .C2(new_n491), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n752), .A2(new_n755), .A3(KEYINPUT42), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n751), .B2(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  NAND3_X1  g574(.A1(new_n755), .A2(new_n672), .A3(new_n750), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT106), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n755), .A2(new_n750), .A3(new_n763), .A4(new_n672), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  NAND3_X1  g580(.A1(new_n653), .A2(new_n632), .A3(new_n656), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT109), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n248), .A2(new_n625), .A3(new_n250), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(KEYINPUT43), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n626), .A2(new_n627), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n771), .B1(new_n772), .B2(new_n625), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT108), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n769), .A2(KEYINPUT43), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n771), .A3(new_n625), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n768), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT110), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n750), .B(KEYINPUT111), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n780), .B2(new_n781), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n768), .A2(new_n785), .A3(KEYINPUT44), .A4(new_n779), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n782), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT107), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n392), .A2(new_n393), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n788), .B(G469), .C1(new_n789), .C2(KEYINPUT45), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(KEYINPUT45), .ZN(new_n791));
  NAND2_X1  g605(.A1(KEYINPUT45), .A2(G469), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n394), .A2(KEYINPUT107), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n395), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n388), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT46), .B1(new_n794), .B2(new_n395), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n711), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n798), .A2(new_n675), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n787), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G137), .ZN(G39));
  NAND2_X1  g615(.A1(new_n798), .A2(KEYINPUT47), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n493), .A2(new_n561), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT47), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n804), .B(new_n711), .C1(new_n796), .C2(new_n797), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n802), .A2(new_n752), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(KEYINPUT112), .B(G140), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(G42));
  NOR2_X1   g622(.A1(G952), .A2(G953), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT119), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n775), .A2(new_n776), .A3(new_n256), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n737), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n701), .A2(KEYINPUT116), .A3(new_n563), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n722), .B2(new_n562), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n813), .A2(new_n689), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n817), .A2(KEYINPUT118), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT117), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT118), .B1(new_n817), .B2(new_n818), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(new_n823), .A3(new_n818), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n819), .A2(new_n821), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n802), .A2(new_n805), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n698), .A2(new_n700), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n828), .A2(KEYINPUT115), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(KEYINPUT115), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n402), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n783), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n813), .ZN(new_n834));
  INV_X1    g648(.A(new_n750), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n687), .A2(new_n835), .A3(new_n722), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n561), .A3(new_n256), .ZN(new_n837));
  INV_X1    g651(.A(new_n772), .ZN(new_n838));
  OR3_X1    g652(.A1(new_n837), .A2(new_n838), .A3(new_n625), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n812), .A2(new_n722), .A3(new_n835), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n744), .B2(new_n747), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n834), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n811), .B1(new_n826), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n834), .A2(new_n841), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(KEYINPUT51), .A3(new_n825), .A4(new_n839), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n813), .A2(new_n742), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n845), .A3(new_n252), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n702), .A2(new_n491), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n557), .A3(new_n560), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n840), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT48), .Z(new_n851));
  NOR2_X1   g665(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n619), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n772), .A2(new_n294), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n628), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n633), .A3(new_n855), .A4(new_n561), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n708), .A2(new_n856), .A3(new_n659), .A4(new_n616), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n725), .A2(new_n740), .A3(new_n705), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n762), .A2(new_n764), .B1(new_n756), .B2(new_n758), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n295), .A2(new_n246), .A3(new_n638), .A4(new_n670), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n664), .A2(new_n666), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n838), .A2(new_n625), .A3(new_n670), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n743), .A2(new_n657), .A3(KEYINPUT105), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n746), .B1(new_n745), .B2(new_n666), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n862), .B1(new_n866), .B2(new_n753), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n859), .B(new_n860), .C1(new_n835), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n664), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n869), .B(new_n710), .C1(new_n672), .C2(new_n693), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n615), .A2(new_n838), .A3(new_n294), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n557), .A2(new_n655), .A3(new_n671), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n687), .A3(new_n753), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n748), .A2(new_n870), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT52), .B1(new_n875), .B2(KEYINPUT113), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n868), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT53), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n875), .A2(KEYINPUT52), .ZN(new_n880));
  INV_X1    g694(.A(new_n753), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n863), .B(new_n881), .C1(new_n864), .C2(new_n865), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n750), .B1(new_n882), .B2(new_n862), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n880), .A2(new_n860), .A3(new_n883), .A4(new_n859), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n875), .A2(KEYINPUT52), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT54), .B1(new_n879), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT114), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n885), .B1(new_n884), .B2(new_n886), .ZN(new_n890));
  INV_X1    g704(.A(new_n868), .ZN(new_n891));
  INV_X1    g705(.A(new_n876), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT53), .A4(new_n878), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n890), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n897), .B(KEYINPUT54), .C1(new_n879), .C2(new_n887), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n852), .A2(new_n889), .A3(new_n896), .A4(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n837), .A2(new_n628), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n810), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n828), .B(KEYINPUT49), .Z(new_n902));
  NOR4_X1   g716(.A1(new_n902), .A2(new_n563), .A3(new_n402), .A4(new_n769), .ZN(new_n903));
  INV_X1    g717(.A(new_n687), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n561), .A3(new_n904), .A4(new_n689), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n905), .ZN(G75));
  AOI21_X1  g720(.A(new_n233), .B1(new_n890), .B2(new_n893), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT56), .B1(new_n907), .B2(G210), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n597), .B1(new_n601), .B2(new_n602), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n573), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT55), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n908), .A2(new_n911), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n251), .A2(G952), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(G51));
  XOR2_X1   g729(.A(new_n395), .B(KEYINPUT57), .Z(new_n916));
  AOI21_X1  g730(.A(new_n894), .B1(new_n890), .B2(new_n893), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n916), .B1(new_n895), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(KEYINPUT120), .B(new_n916), .C1(new_n895), .C2(new_n917), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n718), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n794), .B(KEYINPUT121), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n907), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n914), .B1(new_n922), .B2(new_n924), .ZN(G54));
  NAND3_X1  g739(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  INV_X1    g740(.A(new_n231), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n914), .ZN(G60));
  AND2_X1   g744(.A1(new_n620), .A2(new_n621), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n889), .A2(new_n896), .A3(new_n898), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n624), .B(KEYINPUT59), .Z(new_n933));
  AOI21_X1  g747(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n931), .B(new_n933), .C1(new_n895), .C2(new_n917), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n914), .A3(new_n936), .ZN(G63));
  NAND2_X1  g751(.A1(new_n890), .A2(new_n893), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n651), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  INV_X1    g756(.A(new_n914), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n938), .A2(new_n940), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n558), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n947), .A2(new_n943), .A3(new_n941), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n945), .B(new_n948), .ZN(G66));
  OAI21_X1  g763(.A(G953), .B1(new_n259), .B2(new_n571), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n859), .B2(G953), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n909), .B1(G898), .B2(new_n251), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G69));
  NAND2_X1  g767(.A1(new_n452), .A2(new_n434), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n213), .A2(new_n216), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(new_n957), .Z(new_n958));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n748), .A2(new_n870), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n860), .A2(new_n806), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n872), .A2(new_n849), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n787), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n961), .B(new_n963), .C1(new_n965), .C2(new_n799), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n251), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n251), .A2(G900), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n959), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n799), .B1(new_n787), .B2(new_n964), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n971), .A2(new_n960), .A3(new_n962), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n959), .B(new_n969), .C1(new_n972), .C2(G953), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n958), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n968), .B1(new_n299), .B2(G953), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT126), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n961), .A2(new_n691), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT62), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n961), .A2(new_n691), .A3(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n849), .A2(new_n855), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n984), .A2(new_n677), .A3(new_n835), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n983), .A2(new_n800), .A3(new_n806), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n958), .B1(new_n986), .B2(new_n251), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n975), .A2(new_n978), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n958), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n969), .B1(new_n972), .B2(G953), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT125), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(new_n992), .B2(new_n973), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n977), .B1(new_n993), .B2(new_n987), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n989), .A2(new_n994), .ZN(G72));
  NAND2_X1  g809(.A1(G472), .A2(G902), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT63), .Z(new_n997));
  INV_X1    g811(.A(new_n859), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n997), .B1(new_n986), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n914), .B1(new_n999), .B2(new_n683), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n997), .B1(new_n966), .B2(new_n998), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n1001), .A2(new_n462), .A3(new_n470), .ZN(new_n1002));
  AOI21_X1  g816(.A(KEYINPUT127), .B1(new_n470), .B2(new_n433), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n470), .A2(new_n433), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n997), .B(new_n1005), .C1(new_n879), .C2(new_n887), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n1000), .A2(new_n1002), .A3(new_n1006), .ZN(G57));
endmodule


