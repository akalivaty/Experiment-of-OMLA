//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n575, new_n576, new_n577, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n590, new_n591, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n634, new_n635, new_n637, new_n638, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n463), .A2(G2105), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n467), .A2(G2105), .B1(G101), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(new_n461), .A3(G2104), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(new_n464), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT64), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n472), .A2(G137), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  INV_X1    g052(.A(G100), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n478), .A2(new_n473), .A3(KEYINPUT65), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT65), .B1(new_n478), .B2(new_n473), .ZN(new_n480));
  OAI221_X1 g055(.A(G2104), .B1(G112), .B2(new_n473), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n474), .A2(new_n471), .A3(G2105), .A4(new_n464), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n474), .A2(new_n471), .A3(new_n473), .A4(new_n464), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n484), .B1(G136), .B2(new_n486), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n474), .A2(new_n471), .A3(new_n464), .A4(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n462), .A2(new_n464), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n488), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n490), .A2(KEYINPUT4), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(G114), .B2(new_n473), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n483), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n493), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G62), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(KEYINPUT67), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n501), .A2(new_n504), .A3(G62), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n500), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(new_n500), .B2(KEYINPUT66), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .A3(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(new_n511), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n501), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n513), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n506), .A2(new_n517), .ZN(G166));
  AND2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT68), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(new_n507), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n521), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n510), .A2(KEYINPUT6), .A3(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT6), .B1(new_n510), .B2(G651), .ZN(new_n530));
  OAI211_X1 g105(.A(G51), .B(G543), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n509), .A2(new_n511), .B1(new_n523), .B2(new_n525), .ZN(new_n533));
  AND3_X1   g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(new_n540), .A3(new_n535), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n533), .A2(G89), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(KEYINPUT70), .B1(new_n532), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n515), .A2(G89), .A3(new_n501), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n538), .A2(new_n541), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n528), .A2(new_n544), .A3(new_n545), .A4(new_n531), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n543), .A2(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  XOR2_X1   g125(.A(KEYINPUT71), .B(G90), .Z(new_n551));
  NAND2_X1  g126(.A1(new_n533), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n512), .A2(G52), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n521), .A2(new_n526), .ZN(new_n556));
  INV_X1    g131(.A(G64), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n554), .B1(G651), .B2(new_n558), .ZN(G171));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n521), .A2(new_n526), .A3(G56), .ZN(new_n561));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n561), .A2(KEYINPUT72), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT72), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  NOR3_X1   g139(.A1(new_n563), .A2(new_n564), .A3(new_n500), .ZN(new_n565));
  AOI22_X1  g140(.A1(G81), .A2(new_n533), .B1(new_n512), .B2(G43), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n560), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n561), .A2(new_n562), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n569), .B2(KEYINPUT72), .ZN(new_n570));
  OAI211_X1 g145(.A(KEYINPUT73), .B(new_n566), .C1(new_n570), .C2(new_n563), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(G153));
  NAND4_X1  g148(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT8), .ZN(new_n576));
  NAND4_X1  g151(.A1(G319), .A2(G483), .A3(G661), .A4(new_n576), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT74), .Z(G188));
  NAND2_X1  g153(.A1(new_n515), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT9), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n512), .A2(new_n582), .A3(G53), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n581), .A2(new_n583), .B1(G91), .B2(new_n533), .ZN(new_n584));
  OAI21_X1  g159(.A(G65), .B1(new_n519), .B2(new_n520), .ZN(new_n585));
  NAND2_X1  g160(.A1(G78), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n500), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT75), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G299));
  NAND2_X1  g164(.A1(new_n558), .A2(G651), .ZN(new_n590));
  INV_X1    g165(.A(new_n554), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G301));
  INV_X1    g167(.A(G166), .ZN(G303));
  AND2_X1   g168(.A1(new_n521), .A2(new_n526), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n594), .B2(G74), .ZN(new_n595));
  AOI22_X1  g170(.A1(G87), .A2(new_n533), .B1(new_n512), .B2(G49), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G288));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n519), .A2(new_n520), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n533), .A2(G86), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n512), .A2(G48), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT76), .ZN(G305));
  NAND2_X1  g181(.A1(new_n594), .A2(G60), .ZN(new_n607));
  NAND2_X1  g182(.A1(G72), .A2(G543), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n500), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n512), .A2(G47), .ZN(new_n610));
  INV_X1    g185(.A(G85), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(new_n516), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G290));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n516), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n533), .A2(KEYINPUT10), .A3(G92), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT77), .ZN(new_n620));
  INV_X1    g195(.A(G79), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n507), .ZN(new_n622));
  NAND3_X1  g197(.A1(KEYINPUT77), .A2(G79), .A3(G543), .ZN(new_n623));
  INV_X1    g198(.A(G66), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n622), .B(new_n623), .C1(new_n599), .C2(new_n624), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n625), .A2(G651), .B1(G54), .B2(new_n512), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n628), .B2(G171), .ZN(G284));
  OAI21_X1  g205(.A(new_n629), .B1(new_n628), .B2(G171), .ZN(G321));
  MUX2_X1   g206(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g207(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g208(.A(new_n627), .ZN(new_n634));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G860), .ZN(G148));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n572), .B2(G868), .ZN(G323));
  XOR2_X1   g214(.A(KEYINPUT78), .B(KEYINPUT11), .Z(new_n640));
  XNOR2_X1  g215(.A(G323), .B(new_n640), .ZN(G282));
  NAND2_X1  g216(.A1(new_n491), .A2(new_n468), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2100), .Z(new_n646));
  OR2_X1    g221(.A1(G99), .A2(G2105), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n647), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n648));
  INV_X1    g223(.A(G123), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n483), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n486), .B2(G135), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n652), .A2(G2096), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(G2096), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n646), .A2(new_n653), .A3(new_n654), .ZN(G156));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT80), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT14), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n660), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n669), .ZN(new_n671));
  AND3_X1   g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(G401));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT81), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2084), .B(G2090), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n674), .B2(new_n677), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n676), .B2(new_n677), .ZN(new_n681));
  INV_X1    g256(.A(new_n677), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n682), .A2(new_n678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT18), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n679), .A2(new_n681), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G2096), .B(G2100), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT19), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  AND2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n695), .A2(new_n696), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(new_n702), .B(new_n701), .S(new_n694), .Z(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1991), .B(G1996), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1981), .B(G1986), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n706), .A2(new_n707), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n706), .A2(new_n707), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n712), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(G229));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G22), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G166), .B2(new_n717), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1971), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n717), .A2(G23), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G288), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT33), .B(G1976), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G6), .A2(G16), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT76), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n605), .B(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n726), .B1(new_n728), .B2(G16), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT32), .B(G1981), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n725), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(KEYINPUT34), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT34), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n725), .A2(new_n735), .A3(new_n731), .A4(new_n732), .ZN(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G25), .ZN(new_n738));
  INV_X1    g313(.A(G119), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n473), .A2(G107), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n483), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G131), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n485), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n738), .B1(new_n745), .B2(new_n737), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT35), .B(G1991), .Z(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n746), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(G290), .A2(G16), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n717), .A2(G24), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G1986), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n750), .A2(G1986), .A3(new_n751), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n749), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n734), .A2(new_n736), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(KEYINPUT36), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT83), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(KEYINPUT83), .A3(KEYINPUT36), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT36), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n734), .A2(new_n736), .A3(new_n763), .A4(new_n756), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(KEYINPUT84), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(KEYINPUT84), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n737), .A2(G35), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G162), .B2(new_n737), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT29), .Z(new_n770));
  INV_X1    g345(.A(G2090), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT88), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n717), .A2(G19), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n572), .B2(new_n717), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(G1341), .Z(new_n776));
  NOR2_X1   g351(.A1(new_n770), .A2(new_n771), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G21), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G168), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1966), .ZN(new_n780));
  NOR2_X1   g355(.A1(G4), .A2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n634), .B2(G16), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(G1348), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(G1348), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n737), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  INV_X1    g361(.A(G128), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n473), .A2(G116), .ZN(new_n788));
  OAI21_X1  g363(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n483), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G140), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n485), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n786), .B1(new_n793), .B2(new_n737), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n783), .B(new_n784), .C1(G2067), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n717), .A2(G20), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT23), .Z(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G299), .B2(G16), .ZN(new_n798));
  INV_X1    g373(.A(G1956), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n777), .A2(new_n780), .A3(new_n795), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n737), .A2(G33), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT25), .Z(new_n804));
  AOI22_X1  g379(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n473), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G139), .B2(new_n486), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n802), .B1(new_n807), .B2(new_n737), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT85), .ZN(new_n809));
  INV_X1    g384(.A(G2072), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G28), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(KEYINPUT30), .ZN(new_n813));
  AOI21_X1  g388(.A(G29), .B1(new_n812), .B2(KEYINPUT30), .ZN(new_n814));
  OR2_X1    g389(.A1(KEYINPUT31), .A2(G11), .ZN(new_n815));
  NAND2_X1  g390(.A1(KEYINPUT31), .A2(G11), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n813), .A2(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT24), .B(G34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(new_n737), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT86), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n476), .B2(new_n737), .ZN(new_n821));
  INV_X1    g396(.A(G2084), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n817), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n822), .B2(new_n821), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n811), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n651), .A2(G29), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT87), .ZN(new_n827));
  NOR2_X1   g402(.A1(G27), .A2(G29), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G164), .B2(G29), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n827), .B1(G2078), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n737), .A2(G32), .ZN(new_n831));
  NAND3_X1  g406(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT26), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n834), .A2(new_n835), .B1(G105), .B2(new_n468), .ZN(new_n836));
  INV_X1    g411(.A(G129), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n483), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n486), .B2(G141), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n831), .B1(new_n839), .B2(new_n737), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT27), .B(G1996), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n841), .A2(new_n842), .B1(G2067), .B2(new_n794), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n717), .A2(G5), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(G171), .B2(new_n717), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G1961), .ZN(new_n847));
  INV_X1    g422(.A(new_n842), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n846), .A2(new_n847), .B1(new_n840), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n829), .ZN(new_n850));
  INV_X1    g425(.A(G2078), .ZN(new_n851));
  AOI22_X1  g426(.A1(G1961), .A2(new_n845), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n830), .A2(new_n843), .A3(new_n849), .A4(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n809), .A2(new_n810), .ZN(new_n854));
  NOR3_X1   g429(.A1(new_n825), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n773), .A2(new_n776), .A3(new_n801), .A4(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT89), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n762), .A2(new_n767), .B1(new_n858), .B2(new_n859), .ZN(G311));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n760), .A2(new_n765), .A3(new_n766), .A4(new_n761), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(G150));
  XOR2_X1   g438(.A(KEYINPUT93), .B(G860), .Z(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT91), .B(G55), .Z(new_n866));
  AOI22_X1  g441(.A1(G93), .A2(new_n533), .B1(new_n512), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g442(.A1(new_n594), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(new_n500), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n568), .A2(new_n571), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT92), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g447(.A(KEYINPUT92), .B(new_n867), .C1(new_n868), .C2(new_n500), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n872), .B(new_n873), .C1(new_n565), .C2(new_n567), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n634), .A2(G559), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(KEYINPUT90), .B(KEYINPUT38), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n865), .B1(new_n879), .B2(KEYINPUT39), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(KEYINPUT39), .B2(new_n879), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n872), .A2(new_n873), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n865), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT37), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(G145));
  XOR2_X1   g460(.A(KEYINPUT98), .B(G37), .Z(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n644), .ZN(new_n888));
  OR2_X1    g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n889), .B(G2104), .C1(G118), .C2(new_n473), .ZN(new_n890));
  INV_X1    g465(.A(G142), .ZN(new_n891));
  INV_X1    g466(.A(G130), .ZN(new_n892));
  OAI221_X1 g467(.A(new_n890), .B1(new_n485), .B2(new_n891), .C1(new_n892), .C2(new_n483), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n893), .A2(new_n745), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT96), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n745), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n888), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(new_n644), .A3(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT97), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(new_n902), .A3(KEYINPUT97), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G114), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n494), .B1(new_n908), .B2(G2105), .ZN(new_n909));
  AND4_X1   g484(.A1(G2105), .A2(new_n474), .A3(new_n471), .A4(new_n464), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(G126), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n491), .A2(new_n492), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT94), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT94), .B1(new_n493), .B2(new_n498), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n793), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n793), .B1(new_n916), .B2(new_n917), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n839), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n920), .ZN(new_n922));
  INV_X1    g497(.A(new_n839), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n918), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT95), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n807), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n921), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n921), .A2(new_n924), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n807), .B(KEYINPUT95), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n907), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n927), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n905), .A2(new_n932), .A3(new_n906), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n651), .B(new_n476), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(G162), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n887), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n932), .A2(new_n903), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n936), .B(KEYINPUT99), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n933), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT100), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT100), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n938), .A2(new_n933), .A3(new_n942), .A4(new_n939), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n937), .A2(new_n944), .A3(KEYINPUT40), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT40), .B1(new_n937), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(G395));
  NOR2_X1   g522(.A1(new_n882), .A2(G868), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n875), .B(new_n637), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n533), .A2(G91), .ZN(new_n950));
  INV_X1    g525(.A(new_n583), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n582), .B1(new_n512), .B2(G53), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT75), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n587), .B(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n627), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n584), .A2(new_n588), .A3(new_n619), .A4(new_n626), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n949), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(G290), .A2(G305), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n728), .A2(new_n613), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G288), .ZN(new_n964));
  NAND2_X1  g539(.A1(G303), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(G166), .A2(G288), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT101), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n961), .A2(new_n962), .B1(new_n965), .B2(new_n966), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n971), .ZN(new_n975));
  NAND2_X1  g550(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n975), .B(new_n976), .C1(new_n968), .C2(new_n972), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n958), .A2(KEYINPUT41), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT41), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n956), .A2(new_n957), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n949), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n960), .A2(new_n974), .A3(new_n977), .A4(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT102), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n974), .A2(new_n977), .ZN(new_n986));
  INV_X1    g561(.A(new_n982), .ZN(new_n987));
  OAI211_X1 g562(.A(KEYINPUT103), .B(new_n986), .C1(new_n987), .C2(new_n959), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n959), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n985), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n983), .A2(new_n984), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(new_n628), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n948), .B1(new_n992), .B2(new_n994), .ZN(G295));
  AOI21_X1  g570(.A(new_n948), .B1(new_n992), .B2(new_n994), .ZN(G331));
  INV_X1    g571(.A(new_n958), .ZN(new_n997));
  OAI21_X1  g572(.A(G171), .B1(new_n543), .B2(new_n548), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n532), .A2(KEYINPUT70), .A3(new_n542), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n546), .A2(new_n547), .ZN(new_n1000));
  NAND3_X1  g575(.A1(G301), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n870), .A2(new_n1002), .A3(new_n874), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n870), .B2(new_n874), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n997), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1002), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n875), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n870), .A2(new_n1002), .A3(new_n874), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n981), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n968), .A2(new_n972), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1005), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G37), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1010), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT43), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1010), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT104), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n980), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT104), .A4(new_n979), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n978), .A3(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1007), .A2(new_n1008), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n958), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1016), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n886), .A4(new_n1011), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1015), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT105), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT105), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1029), .B(KEYINPUT44), .C1(new_n1015), .C2(new_n1025), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1023), .A2(new_n886), .A3(new_n1011), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1027), .B1(new_n1031), .B2(KEYINPUT43), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1016), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(new_n1024), .A3(new_n1012), .A4(new_n1011), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT106), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1011), .A2(new_n886), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1007), .A2(new_n1008), .A3(new_n1020), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1010), .B1(new_n1005), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT43), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AND4_X1   g615(.A1(KEYINPUT106), .A2(new_n1040), .A3(KEYINPUT44), .A4(new_n1035), .ZN(new_n1041));
  OAI22_X1  g616(.A1(new_n1028), .A2(new_n1030), .B1(new_n1036), .B2(new_n1041), .ZN(G397));
  INV_X1    g617(.A(G1384), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n916), .A2(new_n917), .A3(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n467), .A2(G2105), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n468), .A2(G101), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n475), .A2(new_n1047), .A3(G40), .A4(new_n1048), .ZN(new_n1049));
  OR3_X1    g624(.A1(new_n1046), .A2(KEYINPUT108), .A3(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT108), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1051));
  INV_X1    g626(.A(G2067), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n793), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(G2067), .B1(new_n790), .B2(new_n792), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1053), .A2(KEYINPUT109), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT109), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n839), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1996), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1050), .A2(new_n1051), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1050), .A2(new_n1058), .A3(new_n839), .A4(new_n1051), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT110), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1061), .A3(KEYINPUT110), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n745), .B(new_n747), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1063), .A2(new_n1064), .A3(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n613), .B(new_n753), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1043), .B1(new_n493), .B2(new_n498), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT45), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1049), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1384), .B1(new_n911), .B2(new_n914), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1045), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1077), .A3(new_n851), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT122), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1074), .A2(new_n1077), .A3(new_n1080), .A4(new_n851), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(KEYINPUT53), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n1075), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1049), .B1(new_n1075), .B2(new_n1084), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1072), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT45), .A4(new_n1043), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1049), .B1(new_n1072), .B2(new_n1045), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n851), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1088), .A2(new_n847), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1082), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1088), .A2(new_n847), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1049), .A2(new_n1092), .A3(G2078), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1046), .A2(new_n1089), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1096), .A2(new_n1097), .A3(G301), .A4(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT123), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1093), .A2(new_n1102), .A3(G301), .A4(new_n1099), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1095), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1107));
  INV_X1    g682(.A(G1971), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1088), .B2(G2090), .ZN(new_n1110));
  INV_X1    g685(.A(G8), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G166), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1110), .A2(new_n1114), .A3(G8), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1072), .A2(new_n1049), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n595), .A2(G1976), .A3(new_n596), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(G8), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT113), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1072), .A2(new_n1049), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(new_n1111), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT113), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(new_n1117), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1119), .A2(KEYINPUT52), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1976), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT52), .B1(G288), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1121), .A2(new_n1117), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n605), .A2(G1981), .ZN(new_n1128));
  INV_X1    g703(.A(G1981), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n602), .A2(new_n1129), .A3(new_n603), .A4(new_n604), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(KEYINPUT49), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT49), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g709(.A(KEYINPUT114), .B(KEYINPUT49), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1121), .B(new_n1131), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1115), .A2(new_n1124), .A3(new_n1127), .A4(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1049), .B1(new_n1072), .B2(KEYINPUT50), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1138), .A2(KEYINPUT116), .B1(new_n1084), .B2(new_n1075), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(KEYINPUT116), .B2(new_n1138), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1109), .B1(new_n1140), .B2(G2090), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1114), .B1(new_n1141), .B2(G8), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT117), .B(G2084), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1146));
  INV_X1    g721(.A(G1966), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(G8), .B1(new_n1149), .B2(G286), .ZN(new_n1150));
  AOI21_X1  g725(.A(G168), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT51), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT51), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1153), .B(G8), .C1(new_n1149), .C2(G286), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1093), .A2(new_n1099), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(G171), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1157), .B(KEYINPUT54), .C1(G171), .C2(new_n1094), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1106), .A2(new_n1143), .A3(new_n1155), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1138), .A2(KEYINPUT116), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(KEYINPUT50), .B2(new_n1072), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1138), .A2(KEYINPUT116), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n799), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(KEYINPUT56), .B(G2072), .Z(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT119), .B1(new_n1107), .B2(new_n1164), .ZN(new_n1165));
  OR3_X1    g740(.A1(new_n1107), .A2(KEYINPUT119), .A3(new_n1164), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1163), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1163), .A2(KEYINPUT120), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1170));
  XOR2_X1   g745(.A(G299), .B(KEYINPUT57), .Z(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1163), .A2(new_n1165), .A3(new_n1166), .A4(new_n1171), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1174), .A2(KEYINPUT61), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1174), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(G1348), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1088), .A2(new_n1181), .B1(new_n1052), .B2(new_n1120), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1182), .A2(new_n1183), .A3(new_n634), .ZN(new_n1184));
  XOR2_X1   g759(.A(KEYINPUT58), .B(G1341), .Z(new_n1185));
  NAND2_X1  g760(.A1(new_n1116), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1089), .A2(new_n1090), .A3(new_n1058), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1116), .A2(KEYINPUT121), .A3(new_n1185), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT59), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1191), .A2(new_n1192), .A3(new_n572), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1192), .B1(new_n1191), .B2(new_n572), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1184), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1182), .A2(new_n627), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1182), .A2(new_n627), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1183), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1176), .A2(new_n1180), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1173), .A2(new_n1196), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1174), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1159), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1115), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1124), .A2(new_n1127), .A3(new_n1136), .ZN(new_n1205));
  NOR2_X1   g780(.A1(G286), .A2(new_n1111), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1149), .A2(KEYINPUT63), .A3(new_n1206), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1110), .A2(G8), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT118), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1114), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1110), .A2(KEYINPUT118), .A3(G8), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1208), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1149), .A2(new_n1206), .ZN(new_n1215));
  NOR3_X1   g790(.A1(new_n1137), .A2(new_n1142), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1214), .B1(new_n1216), .B2(KEYINPUT63), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1136), .A2(new_n1125), .A3(new_n964), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(new_n1130), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1219), .A2(new_n1121), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT115), .ZN(new_n1221));
  OAI211_X1 g796(.A(new_n1220), .B(new_n1221), .C1(new_n1115), .C2(new_n1205), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1121), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1223), .B1(new_n1218), .B2(new_n1130), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1205), .A2(new_n1115), .ZN(new_n1225));
  OAI21_X1  g800(.A(KEYINPUT115), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1222), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1155), .A2(KEYINPUT62), .ZN(new_n1228));
  NOR3_X1   g803(.A1(new_n1137), .A2(new_n1142), .A3(new_n1095), .ZN(new_n1229));
  INV_X1    g804(.A(KEYINPUT62), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1152), .A2(new_n1230), .A3(new_n1154), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1228), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1217), .A2(new_n1227), .A3(new_n1232), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1071), .B1(new_n1203), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g809(.A(new_n1064), .ZN(new_n1235));
  NOR2_X1   g810(.A1(new_n1235), .A2(new_n1062), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n745), .A2(new_n747), .ZN(new_n1237));
  XOR2_X1   g812(.A(new_n1237), .B(KEYINPUT124), .Z(new_n1238));
  AOI22_X1  g813(.A1(new_n1236), .A2(new_n1238), .B1(new_n1052), .B2(new_n793), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1066), .A2(new_n1057), .ZN(new_n1240));
  INV_X1    g815(.A(KEYINPUT46), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1241), .B1(new_n1066), .B2(new_n1058), .ZN(new_n1242));
  NOR3_X1   g817(.A1(new_n1065), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1243));
  OAI21_X1  g818(.A(new_n1240), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  AND2_X1   g819(.A1(new_n1244), .A2(KEYINPUT47), .ZN(new_n1245));
  NOR2_X1   g820(.A1(new_n1244), .A2(KEYINPUT47), .ZN(new_n1246));
  OAI22_X1  g821(.A1(new_n1239), .A2(new_n1065), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NOR3_X1   g822(.A1(new_n1065), .A2(G1986), .A3(G290), .ZN(new_n1248));
  XNOR2_X1  g823(.A(new_n1248), .B(KEYINPUT48), .ZN(new_n1249));
  INV_X1    g824(.A(KEYINPUT125), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1069), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g826(.A1(new_n1236), .A2(KEYINPUT125), .A3(new_n1068), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1249), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g828(.A1(new_n1247), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1234), .A2(new_n1254), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g830(.A1(new_n689), .A2(G319), .A3(new_n690), .ZN(new_n1257));
  OR3_X1    g831(.A1(new_n1257), .A2(G401), .A3(KEYINPUT126), .ZN(new_n1258));
  OAI21_X1  g832(.A(KEYINPUT126), .B1(new_n1257), .B2(G401), .ZN(new_n1259));
  NAND3_X1  g833(.A1(new_n715), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  AOI21_X1  g834(.A(new_n1260), .B1(new_n937), .B2(new_n944), .ZN(new_n1261));
  NAND2_X1  g835(.A1(new_n1261), .A2(new_n1026), .ZN(G225));
  INV_X1    g836(.A(G225), .ZN(G308));
endmodule


