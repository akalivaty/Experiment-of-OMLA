//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n193), .A3(new_n196), .A4(new_n191), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(KEYINPUT66), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT64), .B1(new_n204), .B2(G146), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(G146), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n201), .B(new_n203), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n200), .A2(G143), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n202), .B(new_n208), .C1(new_n206), .C2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n194), .A2(new_n212), .A3(G131), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n198), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT2), .A2(G113), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT2), .A2(G113), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G119), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G116), .ZN(new_n219));
  INV_X1    g033(.A(G116), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G119), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n215), .A2(new_n219), .A3(new_n221), .A4(new_n216), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(KEYINPUT69), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n217), .A2(new_n222), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n201), .B1(new_n205), .B2(new_n206), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT67), .ZN(new_n233));
  OAI21_X1  g047(.A(G128), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n200), .A2(G143), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(KEYINPUT67), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT68), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n236), .A2(new_n237), .A3(new_n238), .A4(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(G128), .A3(new_n242), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n206), .A2(new_n209), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n235), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n191), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n189), .A2(G137), .ZN(new_n247));
  OAI21_X1  g061(.A(G131), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n197), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n214), .B(new_n228), .C1(new_n245), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT70), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n242), .A2(G128), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n241), .B1(new_n253), .B2(new_n236), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n244), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n235), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n249), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n259), .A2(new_n260), .A3(new_n214), .A4(new_n228), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n251), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n214), .ZN(new_n263));
  INV_X1    g077(.A(new_n228), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT75), .B1(new_n266), .B2(KEYINPUT28), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n250), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n251), .A2(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(new_n268), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n267), .B1(KEYINPUT75), .B2(new_n271), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT26), .B(G101), .Z(new_n273));
  NOR2_X1   g087(.A1(G237), .A2(G953), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G210), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n273), .B(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n198), .A2(new_n213), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n207), .A2(new_n210), .A3(KEYINPUT65), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT65), .B1(new_n207), .B2(new_n210), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n259), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n251), .A2(new_n261), .B1(new_n287), .B2(new_n264), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n269), .B(new_n278), .C1(new_n288), .C2(new_n268), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n214), .B(KEYINPUT30), .C1(new_n245), .C2(new_n249), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n282), .A2(new_n285), .B1(new_n257), .B2(new_n258), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n264), .B(new_n290), .C1(new_n291), .C2(KEYINPUT30), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n262), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n279), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n289), .A2(new_n280), .A3(new_n294), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n272), .A2(new_n281), .B1(new_n295), .B2(KEYINPUT74), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n289), .A2(new_n294), .A3(new_n297), .A4(new_n280), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n187), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n292), .A2(new_n262), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT31), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n278), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n287), .A2(new_n264), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n268), .B1(new_n262), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n269), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n279), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n292), .A2(new_n262), .A3(new_n304), .A4(new_n278), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT31), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n306), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n313), .A2(KEYINPUT32), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT32), .B1(new_n313), .B2(new_n314), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT73), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(KEYINPUT73), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n302), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G125), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT16), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT77), .B1(new_n321), .B2(G125), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(G140), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n325), .A2(new_n328), .B1(G125), .B2(new_n321), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n324), .B1(new_n329), .B2(new_n323), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G146), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(G140), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n322), .A2(new_n332), .A3(new_n200), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT23), .B1(new_n218), .B2(G128), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n336));
  INV_X1    g150(.A(G128), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G119), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n335), .A2(new_n338), .B1(new_n218), .B2(G128), .ZN(new_n339));
  INV_X1    g153(.A(G110), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(G119), .B(G128), .Z(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT24), .B(G110), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n334), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n331), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n200), .B(new_n324), .C1(new_n329), .C2(new_n323), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n331), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n342), .A2(new_n343), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n339), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n340), .B1(new_n339), .B2(new_n351), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n349), .A2(KEYINPUT78), .A3(new_n354), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n347), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G137), .ZN(new_n360));
  INV_X1    g174(.A(G953), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(G221), .A3(G234), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n360), .B(new_n362), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n363), .B(KEYINPUT79), .Z(new_n364));
  OAI21_X1  g178(.A(KEYINPUT80), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n358), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT78), .B1(new_n349), .B2(new_n354), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n346), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n369));
  INV_X1    g183(.A(new_n364), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n359), .A2(new_n363), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n365), .A2(new_n371), .A3(new_n299), .A4(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G217), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(G234), .B2(new_n299), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(G902), .ZN(new_n379));
  XOR2_X1   g193(.A(new_n379), .B(KEYINPUT81), .Z(new_n380));
  NAND4_X1  g194(.A1(new_n365), .A2(new_n371), .A3(new_n372), .A4(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT82), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n361), .A2(G952), .ZN(new_n385));
  NAND2_X1  g199(.A1(G234), .A2(G237), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g201(.A(KEYINPUT21), .B(G898), .Z(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(G902), .A3(G953), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n337), .A2(G143), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n189), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n204), .A2(G128), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n391), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G116), .B(G122), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n397), .A2(G107), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(G107), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n395), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n396), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n395), .B(G134), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n397), .A2(KEYINPUT14), .A3(G107), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(KEYINPUT14), .B(G107), .C1(new_n220), .C2(G122), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n398), .A2(new_n399), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n401), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT9), .B(G234), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n408), .A2(new_n376), .A3(G953), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n401), .B(new_n409), .C1(new_n404), .C2(new_n406), .ZN(new_n412));
  AOI21_X1  g226(.A(G902), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G113), .B(G122), .ZN(new_n417));
  INV_X1    g231(.A(G104), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G237), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(new_n361), .A3(G214), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n204), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n274), .A2(G143), .A3(G214), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n196), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT17), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n331), .A2(new_n348), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT89), .ZN(new_n427));
  INV_X1    g241(.A(new_n423), .ZN(new_n428));
  AOI21_X1  g242(.A(G143), .B1(new_n274), .B2(G214), .ZN(new_n429));
  OAI21_X1  g243(.A(G131), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n422), .A2(new_n196), .A3(new_n423), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n432), .A2(KEYINPUT17), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT89), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n331), .A2(new_n434), .A3(new_n348), .A4(new_n425), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n427), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n325), .A2(new_n328), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n322), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(G146), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT87), .B1(new_n329), .B2(new_n200), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n333), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n428), .A2(new_n429), .ZN(new_n443));
  NAND2_X1  g257(.A1(KEYINPUT18), .A2(G131), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n443), .A2(new_n444), .B1(new_n424), .B2(KEYINPUT18), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n419), .B1(new_n436), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n436), .A2(new_n419), .A3(new_n446), .ZN(new_n449));
  AOI21_X1  g263(.A(G902), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G475), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n390), .B(new_n416), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT19), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n322), .A2(new_n332), .A3(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n200), .B(new_n455), .C1(new_n329), .C2(new_n454), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n331), .A2(new_n432), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n446), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n419), .B1(new_n458), .B2(KEYINPUT88), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n446), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n449), .ZN(new_n463));
  NOR2_X1   g277(.A1(G475), .A2(G902), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n464), .B(KEYINPUT90), .Z(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n453), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  AOI211_X1 g281(.A(KEYINPUT20), .B(new_n465), .C1(new_n462), .C2(new_n449), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT91), .B1(new_n452), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n446), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n435), .A2(new_n433), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n471), .B1(new_n473), .B2(new_n427), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n474), .A2(new_n419), .B1(new_n461), .B2(new_n459), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT20), .B1(new_n475), .B2(new_n465), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n463), .A2(new_n453), .A3(new_n466), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n415), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n413), .B(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n436), .A2(new_n419), .A3(new_n446), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n299), .B1(new_n481), .B2(new_n447), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n480), .B1(new_n482), .B2(G475), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT91), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n478), .A2(new_n483), .A3(new_n484), .A4(new_n390), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n470), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G221), .B1(new_n408), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n489));
  INV_X1    g303(.A(G107), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(G104), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT3), .ZN(new_n492));
  INV_X1    g306(.A(G101), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT3), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n489), .A2(new_n494), .A3(new_n490), .A4(G104), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n490), .A2(G104), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n492), .A2(new_n493), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n418), .A2(G107), .ZN(new_n499));
  OAI21_X1  g313(.A(G101), .B1(new_n499), .B2(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G128), .B1(new_n206), .B2(new_n232), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n229), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(new_n235), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT10), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n496), .B1(new_n491), .B2(KEYINPUT3), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n493), .B1(new_n508), .B2(new_n495), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n511));
  AOI211_X1 g325(.A(KEYINPUT4), .B(new_n493), .C1(new_n508), .C2(new_n495), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n211), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n257), .A2(KEYINPUT10), .A3(new_n502), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n507), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n282), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n198), .A2(new_n213), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT84), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n520), .A2(new_n514), .A3(new_n507), .A4(new_n515), .ZN(new_n521));
  XNOR2_X1  g335(.A(G110), .B(G140), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n361), .A2(G227), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n522), .B(new_n523), .Z(new_n524));
  AND3_X1   g338(.A1(new_n517), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n505), .B1(new_n257), .B2(new_n502), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n282), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT12), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n529), .A3(new_n282), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n521), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n524), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n525), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(G469), .B1(new_n533), .B2(G902), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n517), .A2(new_n521), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n532), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n528), .A2(new_n521), .A3(new_n530), .A4(new_n524), .ZN(new_n537));
  AOI21_X1  g351(.A(G902), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT85), .B(G469), .Z(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n488), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G214), .B1(G237), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(new_n509), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n545), .A2(new_n228), .A3(new_n512), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT5), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(G113), .C1(KEYINPUT5), .C2(new_n219), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n224), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(new_n501), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT86), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n511), .A2(new_n264), .A3(new_n513), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT86), .ZN(new_n553));
  INV_X1    g367(.A(new_n550), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  XOR2_X1   g369(.A(G110), .B(G122), .Z(new_n556));
  NAND3_X1  g370(.A1(new_n551), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT6), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n551), .A2(new_n555), .A3(KEYINPUT6), .A4(new_n556), .ZN(new_n560));
  INV_X1    g374(.A(new_n556), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n552), .A2(new_n554), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n361), .A2(G224), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n245), .A2(new_n327), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n211), .A2(new_n327), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n564), .A3(new_n566), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G210), .B1(G237), .B2(G902), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT7), .B1(new_n565), .B2(new_n566), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n556), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n549), .A2(new_n501), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n554), .B2(new_n575), .ZN(new_n576));
  OR3_X1    g390(.A1(new_n567), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT7), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n562), .B1(new_n569), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n299), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(new_n572), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n572), .ZN(new_n583));
  INV_X1    g397(.A(new_n570), .ZN(new_n584));
  INV_X1    g398(.A(new_n562), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n557), .B2(new_n558), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n584), .B1(new_n586), .B2(new_n560), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n583), .B1(new_n587), .B2(new_n580), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n543), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n486), .A2(new_n541), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n320), .A2(new_n384), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  NAND2_X1  g406(.A1(new_n313), .A2(new_n299), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G472), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n313), .A2(new_n314), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n534), .A2(new_n540), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n487), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n383), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n482), .A2(G475), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n467), .B2(new_n468), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n411), .A2(new_n412), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(G478), .A3(new_n299), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n413), .A2(G478), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n601), .A2(KEYINPUT92), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n589), .A2(new_n390), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n599), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT34), .B(G104), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT93), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n614), .B(new_n616), .ZN(G6));
  INV_X1    g431(.A(KEYINPUT94), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n477), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n469), .B2(new_n618), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT95), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n416), .B1(new_n482), .B2(G475), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n390), .A4(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n476), .A2(new_n618), .A3(new_n477), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n468), .A2(KEYINPUT94), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n390), .A4(new_n622), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT95), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n623), .A2(new_n627), .A3(new_n589), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n599), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NAND2_X1  g445(.A1(new_n368), .A2(KEYINPUT96), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n359), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n370), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n375), .A2(new_n377), .B1(new_n637), .B2(new_n380), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n596), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n590), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT37), .B(G110), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT97), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n640), .B(new_n642), .ZN(G12));
  AOI21_X1  g457(.A(new_n572), .B1(new_n571), .B2(new_n581), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n587), .A2(new_n583), .A3(new_n580), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n542), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n638), .A2(new_n598), .A3(new_n646), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n320), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n387), .B(KEYINPUT99), .Z(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT98), .B(G900), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n650), .B1(new_n389), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT100), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n620), .A2(new_n622), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n648), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT101), .B(G128), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G30));
  NAND2_X1  g472(.A1(new_n637), .A2(new_n380), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n378), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n601), .A2(new_n480), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n660), .A2(new_n543), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n653), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n541), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n662), .B1(KEYINPUT40), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(KEYINPUT40), .B2(new_n665), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT32), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n595), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT73), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n313), .A2(KEYINPUT32), .A3(new_n314), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n318), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n293), .A2(new_n279), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n270), .A2(new_n278), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n299), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G472), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n582), .A2(new_n588), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n667), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  NOR2_X1   g498(.A1(new_n607), .A2(new_n653), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n648), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  INV_X1    g501(.A(G469), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n538), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n539), .ZN(new_n690));
  AOI211_X1 g504(.A(G902), .B(new_n690), .C1(new_n536), .C2(new_n537), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n689), .A2(new_n691), .A3(new_n488), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n320), .A2(new_n613), .A3(new_n384), .A4(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT41), .B(G113), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT104), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n693), .B(new_n695), .ZN(G15));
  NAND4_X1  g510(.A1(new_n320), .A2(new_n628), .A3(new_n384), .A4(new_n692), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n540), .B(new_n487), .C1(new_n688), .C2(new_n538), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n699), .B1(new_n646), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n589), .A2(new_n692), .A3(KEYINPUT105), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n638), .B1(new_n485), .B2(new_n470), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n320), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  INV_X1    g520(.A(new_n314), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n271), .A2(KEYINPUT75), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT75), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n270), .B2(new_n268), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT106), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n708), .A2(new_n713), .A3(new_n710), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n279), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n306), .A2(new_n312), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n707), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n594), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n646), .A2(new_n700), .ZN(new_n721));
  INV_X1    g535(.A(new_n390), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n661), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n720), .A2(new_n384), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NOR3_X1   g539(.A1(new_n718), .A2(new_n638), .A3(new_n719), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n703), .A3(new_n685), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  NOR2_X1   g542(.A1(new_n315), .A2(new_n316), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n383), .B1(new_n302), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n535), .B2(new_n532), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n732), .B(G469), .C1(new_n533), .C2(new_n731), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n688), .A2(new_n299), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n538), .B2(new_n539), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n488), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n730), .A2(KEYINPUT42), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n582), .A2(new_n588), .A3(new_n542), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n582), .A2(new_n588), .A3(KEYINPUT108), .A4(new_n542), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n685), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n301), .B1(new_n672), .B2(new_n318), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n740), .A2(new_n741), .A3(new_n736), .ZN(new_n747));
  INV_X1    g561(.A(new_n685), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n746), .A2(new_n747), .A3(new_n383), .A4(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n745), .B1(new_n749), .B2(KEYINPUT42), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n740), .A2(new_n741), .A3(new_n736), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n320), .A2(new_n751), .A3(new_n384), .A4(new_n685), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(KEYINPUT109), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n744), .B1(new_n750), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n196), .ZN(G33));
  NAND4_X1  g570(.A1(new_n320), .A2(new_n751), .A3(new_n384), .A4(new_n655), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  INV_X1    g572(.A(new_n742), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n601), .B1(new_n605), .B2(new_n604), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT43), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n596), .A3(new_n660), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n763), .B2(new_n762), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n531), .A2(new_n532), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT107), .B1(new_n766), .B2(new_n525), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n767), .A2(KEYINPUT45), .A3(new_n732), .ZN(new_n768));
  OAI21_X1  g582(.A(G469), .B1(new_n533), .B2(KEYINPUT45), .ZN(new_n769));
  OAI22_X1  g583(.A1(new_n768), .A2(new_n769), .B1(new_n688), .B2(new_n299), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n691), .B1(new_n770), .B2(new_n772), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n487), .A3(new_n664), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n765), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT111), .B(G137), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G39));
  NAND2_X1  g594(.A1(new_n776), .A2(new_n487), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT47), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT47), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n776), .A2(new_n783), .A3(new_n487), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n743), .A2(new_n320), .A3(new_n384), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  NOR2_X1   g601(.A1(new_n689), .A2(new_n691), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT49), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(new_n487), .A3(new_n542), .A4(new_n760), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n790), .A2(new_n678), .A3(new_n682), .A4(new_n383), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT112), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n646), .A2(new_n661), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n660), .A2(new_n653), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n678), .A2(new_n736), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n320), .B(new_n647), .C1(new_n655), .C2(new_n685), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n727), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(KEYINPUT52), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n752), .A2(KEYINPUT109), .A3(new_n753), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT109), .B1(new_n752), .B2(new_n753), .ZN(new_n802));
  OAI22_X1  g616(.A1(new_n801), .A2(new_n802), .B1(new_n743), .B2(new_n737), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n693), .A2(new_n697), .A3(new_n705), .A4(new_n724), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n708), .A2(new_n713), .A3(new_n710), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n713), .B1(new_n708), .B2(new_n710), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n805), .A2(new_n806), .A3(new_n278), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n314), .B1(new_n807), .B2(new_n716), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(new_n660), .A3(new_n594), .A4(new_n685), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT115), .B1(new_n809), .B2(new_n747), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n726), .A2(new_n751), .A3(new_n811), .A4(new_n685), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n483), .A2(new_n541), .A3(new_n620), .A4(new_n654), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n320), .A2(new_n660), .A3(new_n813), .A4(new_n742), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n810), .A2(new_n812), .A3(new_n757), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n601), .A2(new_n816), .A3(new_n606), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n816), .B1(new_n601), .B2(new_n606), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(new_n612), .A3(KEYINPUT114), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n607), .A2(KEYINPUT113), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n817), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n722), .B(new_n543), .C1(new_n582), .C2(new_n588), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n599), .B1(new_n821), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n478), .A2(new_n622), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n612), .A2(new_n828), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n599), .A2(new_n829), .B1(new_n590), .B2(new_n639), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(new_n830), .A3(new_n591), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n815), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n803), .A2(new_n804), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n800), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n803), .A2(new_n832), .A3(KEYINPUT116), .A4(new_n804), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT53), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n757), .A2(new_n810), .A3(new_n812), .A4(new_n814), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n827), .A2(new_n591), .A3(new_n830), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n804), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n834), .B1(new_n840), .B2(new_n755), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n798), .A2(new_n799), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n836), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT54), .B1(new_n837), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n798), .A2(KEYINPUT53), .A3(new_n799), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n833), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n843), .B2(new_n844), .ZN(new_n849));
  XNOR2_X1  g663(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n761), .A2(new_n649), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n384), .A3(new_n720), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n855), .A2(new_n542), .A3(new_n682), .A4(new_n700), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT50), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n759), .A2(new_n700), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n854), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n726), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n678), .A2(new_n383), .A3(new_n387), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n858), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n863), .A2(new_n601), .A3(new_n606), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n857), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n855), .A2(new_n759), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n782), .A2(new_n784), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n788), .A2(new_n488), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n865), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n870), .B(KEYINPUT118), .Z(new_n873));
  AOI21_X1  g687(.A(new_n868), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n866), .B1(new_n865), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n860), .A2(new_n730), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT48), .Z(new_n877));
  INV_X1    g691(.A(new_n703), .ZN(new_n878));
  OAI221_X1 g692(.A(new_n385), .B1(new_n855), .B2(new_n878), .C1(new_n611), .C2(new_n863), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n852), .A2(new_n872), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(G952), .A2(G953), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n792), .B1(new_n882), .B2(new_n883), .ZN(G75));
  NOR2_X1   g698(.A1(new_n563), .A2(new_n570), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n587), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT119), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT55), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(KEYINPUT56), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n887), .A2(KEYINPUT55), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(G210), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n849), .A2(new_n894), .A3(new_n299), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n895), .B2(KEYINPUT56), .ZN(new_n896));
  OAI211_X1 g710(.A(G210), .B(G902), .C1(new_n837), .C2(new_n848), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n898), .A3(new_n892), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n361), .A2(G952), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n896), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT121), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n896), .A2(new_n899), .A3(new_n904), .A4(new_n901), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n905), .ZN(G51));
  NAND2_X1  g720(.A1(new_n536), .A2(new_n537), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n849), .A2(new_n850), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n849), .A2(new_n850), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n734), .B(KEYINPUT57), .Z(new_n911));
  OAI21_X1  g725(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n849), .A2(new_n299), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n768), .A2(new_n769), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n900), .B1(new_n912), .B2(new_n915), .ZN(G54));
  AND2_X1   g730(.A1(KEYINPUT58), .A2(G475), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n913), .A2(new_n463), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n463), .B1(new_n913), .B2(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n900), .ZN(G60));
  INV_X1    g734(.A(new_n603), .ZN(new_n921));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT59), .Z(new_n923));
  NOR2_X1   g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n908), .B2(new_n909), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(KEYINPUT122), .B(new_n924), .C1(new_n908), .C2(new_n909), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n923), .B1(new_n846), .B2(new_n851), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n901), .B1(new_n930), .B2(new_n603), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(new_n843), .A2(new_n844), .ZN(new_n933));
  INV_X1    g747(.A(new_n848), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT60), .Z(new_n937));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n637), .A3(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n935), .A2(new_n937), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n365), .A2(new_n372), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n940), .A2(new_n371), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n901), .B(new_n938), .C1(new_n939), .C2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G66));
  NAND2_X1  g758(.A1(new_n388), .A2(G224), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(G953), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n804), .A2(new_n839), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(G953), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n586), .B(new_n560), .C1(G898), .C2(new_n361), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G69));
  AOI21_X1  g764(.A(new_n361), .B1(G227), .B2(G900), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n796), .A2(new_n727), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n778), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT124), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n730), .A2(new_n793), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n777), .A2(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n786), .A2(new_n757), .A3(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n955), .A2(new_n361), .A3(new_n803), .A4(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n290), .B1(new_n291), .B2(KEYINPUT30), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n455), .B1(new_n329), .B2(new_n454), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(G900), .B2(G953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n962), .B(KEYINPUT123), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n683), .A2(new_n727), .A3(new_n796), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n665), .B1(new_n820), .B2(new_n828), .ZN(new_n970));
  AND4_X1   g784(.A1(new_n320), .A2(new_n970), .A3(new_n384), .A4(new_n742), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n778), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n972), .A2(new_n786), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n966), .B1(new_n974), .B2(G953), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT125), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n965), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n976), .B1(new_n965), .B2(new_n975), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n952), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n965), .A2(new_n975), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT125), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n965), .A2(new_n975), .A3(new_n976), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n951), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n979), .A2(new_n983), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  INV_X1    g800(.A(new_n294), .ZN(new_n987));
  OAI221_X1 g801(.A(new_n986), .B1(new_n674), .B2(new_n987), .C1(new_n837), .C2(new_n845), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT127), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n955), .A2(new_n803), .A3(new_n947), .A4(new_n958), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n986), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n293), .A2(new_n278), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n900), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n969), .A2(new_n947), .A3(new_n973), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n995), .B2(new_n986), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n994), .A3(new_n986), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(new_n278), .A3(new_n293), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n993), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n989), .A2(new_n999), .ZN(G57));
endmodule


