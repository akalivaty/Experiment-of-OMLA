//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n203));
  INV_X1    g002(.A(G120gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G113gat), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G120gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT1), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G127gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G134gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n211));
  OR3_X1    g010(.A1(new_n203), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G148gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT76), .B1(new_n213), .B2(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215));
  INV_X1    g014(.A(G141gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(G148gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(G141gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n218), .A2(new_n219), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(KEYINPUT2), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT77), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT77), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n220), .A2(new_n226), .A3(KEYINPUT2), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n216), .A2(G148gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n230), .A2(new_n231), .B1(G155gat), .B2(G162gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT75), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n221), .B(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n223), .A2(new_n228), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G134gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G127gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n210), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n202), .A2(KEYINPUT67), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT68), .B1(new_n242), .B2(new_n208), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n210), .A2(new_n237), .A3(KEYINPUT67), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT67), .B1(new_n210), .B2(new_n237), .ZN(new_n245));
  OAI211_X1 g044(.A(KEYINPUT68), .B(new_n208), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n212), .B(new_n235), .C1(new_n243), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n218), .A2(new_n219), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n222), .A2(new_n220), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n228), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT78), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n230), .A2(new_n231), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n253), .A3(new_n220), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n252), .B1(new_n251), .B2(new_n254), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n203), .A2(new_n208), .A3(new_n211), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n208), .B1(new_n244), .B2(new_n245), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n261), .B2(new_n246), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n248), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G225gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT3), .B1(new_n255), .B2(new_n256), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n261), .A2(new_n246), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n212), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n235), .A2(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n267), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n268), .A2(new_n273), .A3(new_n235), .A4(new_n212), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n262), .B2(new_n235), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT80), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n248), .A2(KEYINPUT4), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT80), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n274), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n272), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(KEYINPUT39), .B(new_n266), .C1(new_n281), .C2(new_n264), .ZN(new_n282));
  XNOR2_X1  g081(.A(G1gat), .B(G29gat), .ZN(new_n283));
  INV_X1    g082(.A(G85gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT0), .B(G57gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n267), .A2(new_n269), .A3(new_n271), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n278), .A2(new_n279), .A3(new_n274), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n279), .B1(new_n278), .B2(new_n274), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT39), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n293), .A3(new_n265), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n282), .A2(KEYINPUT40), .A3(new_n288), .A4(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n296), .B1(new_n263), .B2(new_n265), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT79), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n274), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n262), .A2(KEYINPUT79), .A3(new_n273), .A4(new_n235), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n299), .A2(new_n300), .A3(new_n278), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n289), .A2(new_n264), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n297), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n265), .A2(KEYINPUT5), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n289), .B(new_n304), .C1(new_n290), .C2(new_n291), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n288), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n295), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n277), .A2(new_n280), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n264), .B1(new_n309), .B2(new_n289), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n287), .B1(new_n310), .B2(new_n293), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT40), .B1(new_n311), .B2(new_n282), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT26), .ZN(new_n317));
  NAND2_X1  g116(.A1(G183gat), .A2(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n320), .A2(KEYINPUT26), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n317), .B(new_n318), .C1(new_n321), .C2(new_n316), .ZN(new_n322));
  OR2_X1    g121(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n324));
  AOI21_X1  g123(.A(G190gat), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n325), .A2(KEYINPUT64), .A3(KEYINPUT28), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT64), .ZN(new_n327));
  INV_X1    g126(.A(G190gat), .ZN(new_n328));
  AND2_X1   g127(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT65), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT65), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n336), .B1(new_n323), .B2(new_n324), .ZN(new_n337));
  OAI211_X1 g136(.A(KEYINPUT28), .B(new_n328), .C1(new_n335), .C2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n322), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n318), .A2(KEYINPUT24), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT24), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(G183gat), .A3(G190gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G183gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n328), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n316), .B(new_n347), .ZN(new_n348));
  AND4_X1   g147(.A1(KEYINPUT25), .A2(new_n346), .A3(new_n348), .A4(new_n319), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n320), .B1(new_n343), .B2(new_n345), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT25), .B1(new_n350), .B2(new_n348), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n315), .B1(new_n339), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G197gat), .B(G204gat), .ZN(new_n354));
  INV_X1    g153(.A(G211gat), .ZN(new_n355));
  INV_X1    g154(.A(G218gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n354), .B1(KEYINPUT22), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n358), .B(new_n359), .Z(new_n360));
  INV_X1    g159(.A(new_n322), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT64), .B1(new_n325), .B2(KEYINPUT28), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n331), .A2(new_n327), .A3(new_n332), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n323), .A2(new_n336), .A3(new_n324), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT65), .B1(new_n329), .B2(new_n330), .ZN(new_n366));
  AOI211_X1 g165(.A(new_n332), .B(G190gat), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n361), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n346), .A2(new_n348), .A3(new_n319), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n350), .A2(KEYINPUT25), .A3(new_n348), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT29), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n353), .B(new_n360), .C1(new_n374), .C2(new_n315), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT72), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n338), .A2(new_n362), .A3(new_n363), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n378), .A2(new_n361), .B1(new_n371), .B2(new_n372), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n314), .B1(new_n379), .B2(KEYINPUT29), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n380), .A2(KEYINPUT72), .A3(new_n360), .A4(new_n353), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n358), .B(new_n359), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT71), .B1(new_n380), .B2(new_n353), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT71), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n373), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n388), .B2(new_n314), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n383), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT73), .B(G64gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(G92gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G8gat), .B(G36gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n382), .A2(KEYINPUT30), .A3(new_n390), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n353), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n385), .ZN(new_n398));
  INV_X1    g197(.A(new_n389), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n360), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n377), .A2(new_n381), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n390), .A2(new_n377), .A3(new_n381), .A4(new_n395), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT30), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT74), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT74), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n408), .A3(new_n405), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n403), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n313), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n360), .B1(new_n271), .B2(new_n387), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT3), .B1(new_n360), .B2(new_n387), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n415), .A2(new_n235), .ZN(new_n416));
  NAND2_X1  g215(.A1(G228gat), .A2(G233gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n412), .A2(new_n413), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n414), .A2(new_n416), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n415), .A2(new_n257), .ZN(new_n420));
  OAI211_X1 g219(.A(G228gat), .B(G233gat), .C1(new_n420), .C2(new_n412), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G22gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n424), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n419), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT31), .B(G50gat), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n425), .A2(new_n429), .A3(new_n427), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n404), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT37), .B1(new_n400), .B2(new_n401), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT37), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n390), .A2(new_n436), .A3(new_n377), .A4(new_n381), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n394), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n434), .B1(new_n438), .B2(KEYINPUT38), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n306), .A2(KEYINPUT6), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443));
  AOI211_X1 g242(.A(new_n443), .B(new_n288), .C1(new_n303), .C2(new_n305), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT84), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT81), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n303), .A2(new_n305), .A3(new_n288), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n447), .B1(new_n448), .B2(new_n306), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n303), .A2(new_n305), .A3(new_n288), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT6), .B1(new_n450), .B2(KEYINPUT81), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n439), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n360), .B1(new_n384), .B2(new_n389), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n454), .B(KEYINPUT37), .C1(new_n360), .C2(new_n397), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT38), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n455), .A2(new_n437), .A3(new_n456), .A4(new_n394), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(KEYINPUT83), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n411), .B(new_n433), .C1(new_n453), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n431), .A2(new_n432), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n444), .B1(new_n449), .B2(new_n451), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n460), .B1(new_n410), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT69), .B1(new_n386), .B2(new_n269), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n386), .A2(new_n269), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT69), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n379), .A2(new_n465), .A3(new_n262), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT32), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT34), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT34), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(KEYINPUT32), .A3(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n463), .A2(new_n468), .A3(new_n466), .A4(new_n464), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT70), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n477), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n473), .B1(new_n470), .B2(KEYINPUT32), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT32), .ZN(new_n481));
  AOI211_X1 g280(.A(new_n481), .B(KEYINPUT34), .C1(new_n467), .C2(new_n469), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n479), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n470), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G43gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n486), .B(new_n487), .Z(new_n488));
  NAND2_X1  g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n478), .A2(new_n483), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n478), .B2(new_n483), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n477), .B1(new_n472), .B2(new_n474), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n480), .A2(new_n482), .A3(new_n479), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n489), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n483), .A3(new_n490), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT36), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n459), .A2(new_n462), .A3(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n403), .A2(new_n407), .A3(new_n409), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n452), .A2(new_n440), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n433), .B1(new_n491), .B2(new_n492), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT35), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n460), .B1(new_n497), .B2(new_n498), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT35), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n446), .A2(new_n452), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n502), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n513), .A2(KEYINPUT89), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(KEYINPUT89), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT16), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(G1gat), .ZN(new_n518));
  INV_X1    g317(.A(G1gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(new_n519), .A3(new_n515), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G8gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT90), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n518), .B(new_n520), .C1(new_n523), .C2(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT87), .B(G29gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  AND2_X1   g328(.A1(KEYINPUT86), .A2(KEYINPUT14), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n528), .A2(G36gat), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(KEYINPUT86), .A2(KEYINPUT14), .ZN(new_n532));
  OR3_X1    g331(.A1(new_n530), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n531), .B(new_n533), .C1(KEYINPUT15), .C2(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n527), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT13), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT88), .B(KEYINPUT17), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n535), .A2(new_n536), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n535), .A2(new_n536), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(KEYINPUT17), .A3(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n543), .A2(new_n526), .A3(new_n525), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n527), .A2(new_n537), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n539), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT18), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT18), .A4(new_n539), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n541), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G169gat), .B(G197gat), .Z(new_n554));
  XNOR2_X1  g353(.A(G113gat), .B(G141gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT12), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n553), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n541), .A2(new_n551), .A3(new_n552), .A4(new_n559), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(KEYINPUT91), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n553), .A2(new_n564), .A3(new_n560), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n512), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n571));
  NAND2_X1  g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  OR2_X1    g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(G57gat), .B(G64gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT9), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n572), .B(new_n573), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT93), .ZN(new_n577));
  INV_X1    g376(.A(G64gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(G57gat), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT94), .B(G57gat), .Z(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(new_n578), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n572), .B1(new_n573), .B2(new_n575), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT21), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(new_n526), .A3(new_n525), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(new_n344), .ZN(new_n587));
  AND2_X1   g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n587), .A2(new_n588), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n571), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  INV_X1    g392(.A(new_n571), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n584), .A2(KEYINPUT21), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G211gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  XOR2_X1   g400(.A(G127gat), .B(G155gat), .Z(new_n602));
  OR3_X1    g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n600), .B2(new_n601), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n596), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n592), .A2(new_n595), .A3(new_n604), .A4(new_n603), .ZN(new_n607));
  AND2_X1   g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  INV_X1    g411(.A(G92gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(KEYINPUT8), .A2(new_n612), .B1(new_n284), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT7), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(new_n284), .B2(new_n613), .ZN(new_n616));
  NAND3_X1  g415(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G99gat), .B(G106gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT97), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n543), .A2(new_n625), .A3(new_n546), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n624), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n537), .A2(new_n629), .B1(KEYINPUT41), .B2(new_n608), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n543), .A2(new_n625), .A3(KEYINPUT98), .A4(new_n546), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n633), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n628), .A2(new_n630), .A3(new_n631), .A4(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n611), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n611), .A3(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n618), .A2(KEYINPUT99), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n584), .A2(new_n629), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n577), .A2(new_n583), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n624), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n584), .A2(new_n629), .A3(KEYINPUT10), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n642), .A2(new_n645), .ZN(new_n651));
  INV_X1    g450(.A(new_n649), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n650), .A2(new_n653), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n606), .A2(new_n607), .A3(new_n640), .A4(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n570), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n503), .B(KEYINPUT100), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g467(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n570), .A2(new_n664), .A3(new_n410), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n570), .A2(KEYINPUT102), .A3(new_n664), .A4(new_n410), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT16), .B(G8gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT103), .Z(new_n676));
  OAI21_X1  g475(.A(new_n669), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n675), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n665), .A2(KEYINPUT42), .A3(new_n410), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n674), .A2(G8gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(G1325gat));
  NAND2_X1  g480(.A1(new_n497), .A2(new_n498), .ZN(new_n682));
  AOI21_X1  g481(.A(G15gat), .B1(new_n665), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n500), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(G15gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT104), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n683), .B1(new_n665), .B2(new_n686), .ZN(G1326gat));
  NAND2_X1  g486(.A1(new_n665), .A2(new_n460), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NAND2_X1  g489(.A1(new_n606), .A2(new_n607), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(new_n640), .A3(new_n661), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n570), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n528), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n666), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n563), .A2(KEYINPUT105), .A3(new_n565), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT105), .B1(new_n563), .B2(new_n565), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n661), .B(KEYINPUT106), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n702), .A2(new_n692), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n462), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g507(.A(KEYINPUT108), .B(new_n460), .C1(new_n410), .C2(new_n461), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n459), .A2(new_n708), .A3(new_n500), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n511), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n634), .A2(new_n611), .A3(new_n636), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n637), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT107), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n512), .B2(new_n714), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(KEYINPUT107), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n706), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n666), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT109), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n724), .A3(new_n666), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n723), .A2(new_n528), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n696), .A2(new_n697), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n698), .A2(new_n726), .A3(new_n727), .ZN(G1328gat));
  NOR2_X1   g527(.A1(new_n502), .A2(G36gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n570), .A2(new_n693), .A3(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT46), .Z(new_n731));
  NAND2_X1  g530(.A1(new_n721), .A2(new_n410), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G36gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1329gat));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n720), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n735), .A2(G43gat), .A3(new_n684), .A4(new_n705), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n568), .A2(new_n569), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT92), .B1(new_n512), .B2(new_n567), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n682), .B(new_n693), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(G43gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI211_X1 g540(.A(KEYINPUT110), .B(KEYINPUT47), .C1(new_n736), .C2(new_n741), .ZN(new_n742));
  OR2_X1    g541(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n743));
  NAND2_X1  g542(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n744));
  AND4_X1   g543(.A1(new_n743), .A2(new_n736), .A3(new_n744), .A4(new_n741), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n742), .A2(new_n745), .ZN(G1330gat));
  AOI21_X1  g545(.A(new_n717), .B1(KEYINPUT107), .B2(new_n715), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n717), .A2(KEYINPUT107), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n460), .B(new_n705), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT112), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n751), .A3(new_n460), .A4(new_n705), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n752), .A3(G50gat), .ZN(new_n753));
  INV_X1    g552(.A(G50gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n460), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT111), .Z(new_n756));
  NAND2_X1  g555(.A1(new_n694), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n753), .A2(KEYINPUT48), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759));
  INV_X1    g558(.A(new_n757), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n754), .B1(new_n721), .B2(new_n460), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(G1331gat));
  AOI21_X1  g562(.A(new_n701), .B1(new_n710), .B2(new_n511), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n691), .A2(new_n714), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n764), .A2(new_n765), .A3(new_n704), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n666), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(new_n580), .ZN(G1332gat));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n410), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT49), .B(G64gat), .Z(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(G1333gat));
  NAND2_X1  g571(.A1(new_n766), .A2(new_n684), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G71gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n766), .A2(new_n682), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(G71gat), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g576(.A1(new_n766), .A2(new_n460), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT114), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT113), .B(G78gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1335gat));
  INV_X1    g580(.A(new_n666), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n782), .A2(G85gat), .A3(new_n662), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n692), .A2(new_n640), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n764), .A2(KEYINPUT51), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT51), .B1(new_n764), .B2(new_n785), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n764), .A2(KEYINPUT51), .A3(new_n785), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(KEYINPUT115), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT116), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n764), .A2(new_n785), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(KEYINPUT115), .A3(new_n790), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n786), .A2(new_n788), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n784), .B1(new_n792), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n692), .A2(new_n662), .A3(new_n701), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n802), .B1(new_n719), .B2(new_n720), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n284), .B1(new_n803), .B2(new_n666), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT117), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n797), .B1(new_n796), .B2(new_n798), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n783), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n803), .A2(new_n666), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G85gat), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n805), .A2(new_n812), .ZN(G1336gat));
  NAND2_X1  g612(.A1(new_n803), .A2(new_n410), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G92gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n789), .A2(new_n791), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n703), .A2(new_n502), .A3(G92gat), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n795), .A2(new_n790), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n814), .A2(G92gat), .B1(new_n821), .B2(new_n818), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n816), .B2(new_n822), .ZN(G1337gat));
  NOR2_X1   g622(.A1(new_n806), .A2(new_n807), .ZN(new_n824));
  INV_X1    g623(.A(G99gat), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n682), .A2(new_n825), .A3(new_n661), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n803), .A2(new_n684), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n824), .A2(new_n826), .B1(new_n827), .B2(new_n825), .ZN(G1338gat));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n803), .A2(new_n829), .A3(new_n460), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n460), .B(new_n801), .C1(new_n747), .C2(new_n748), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT118), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n832), .A3(G106gat), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n703), .A2(G106gat), .A3(new_n433), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT53), .B1(new_n817), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n831), .A2(G106gat), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n821), .A2(new_n834), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT53), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(G1339gat));
  NAND3_X1  g639(.A1(new_n646), .A2(new_n652), .A3(new_n647), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n652), .B1(new_n646), .B2(new_n647), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n659), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n845), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n660), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n699), .A2(new_n700), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n538), .A2(new_n540), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n539), .B1(new_n547), .B2(new_n548), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n558), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n562), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n661), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n640), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n845), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT55), .B1(new_n842), .B2(new_n845), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n861), .A2(new_n714), .A3(new_n660), .A4(new_n855), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n692), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n663), .A2(new_n701), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n505), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n666), .A2(new_n502), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n206), .A3(new_n701), .ZN(new_n872));
  OAI21_X1  g671(.A(G113gat), .B1(new_n870), .B2(new_n566), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1340gat));
  NAND3_X1  g673(.A1(new_n871), .A2(new_n204), .A3(new_n661), .ZN(new_n875));
  OAI21_X1  g674(.A(G120gat), .B1(new_n870), .B2(new_n703), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1341gat));
  NOR2_X1   g676(.A1(new_n870), .A2(new_n691), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(new_n209), .ZN(G1342gat));
  NAND3_X1  g678(.A1(new_n871), .A2(new_n236), .A3(new_n714), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n881));
  OAI21_X1  g680(.A(G134gat), .B1(new_n870), .B2(new_n640), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G1343gat));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n684), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n856), .B1(new_n566), .B2(new_n850), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n640), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n692), .B1(new_n887), .B2(new_n862), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n460), .B1(new_n888), .B2(new_n865), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT57), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n460), .B1(new_n863), .B2(new_n865), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n885), .B(new_n890), .C1(new_n891), .C2(KEYINPUT57), .ZN(new_n892));
  OAI21_X1  g691(.A(G141gat), .B1(new_n892), .B2(new_n566), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT58), .ZN(new_n894));
  INV_X1    g693(.A(new_n891), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n895), .A2(new_n216), .A3(new_n567), .A4(new_n885), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898));
  OAI21_X1  g697(.A(G141gat), .B1(new_n892), .B2(new_n702), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n896), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n900), .B2(KEYINPUT58), .ZN(new_n901));
  AOI211_X1 g700(.A(KEYINPUT119), .B(new_n894), .C1(new_n899), .C2(new_n896), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(G1344gat));
  NAND2_X1  g702(.A1(new_n895), .A2(new_n885), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n213), .A3(new_n661), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT121), .B1(new_n850), .B2(new_n640), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n861), .A2(new_n714), .A3(new_n909), .A4(new_n660), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n910), .A3(new_n855), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n887), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n887), .B2(new_n911), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(new_n692), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n664), .A2(KEYINPUT120), .A3(new_n566), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(new_n663), .B2(new_n567), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT123), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n887), .A2(new_n911), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT122), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n887), .A2(new_n911), .A3(new_n912), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n691), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n916), .A2(new_n918), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n920), .A2(new_n921), .A3(new_n460), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n929), .A2(new_n661), .A3(new_n885), .A4(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n907), .B1(new_n931), .B2(G148gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n907), .B1(new_n892), .B2(new_n662), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(new_n213), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n906), .B1(new_n932), .B2(new_n934), .ZN(G1345gat));
  INV_X1    g734(.A(G155gat), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n892), .A2(new_n936), .A3(new_n691), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n905), .A2(new_n692), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n936), .B2(new_n938), .ZN(G1346gat));
  INV_X1    g738(.A(G162gat), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n892), .A2(new_n940), .A3(new_n640), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n905), .A2(new_n714), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n940), .B2(new_n942), .ZN(G1347gat));
  NOR2_X1   g742(.A1(new_n666), .A2(new_n502), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n867), .A2(new_n944), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n945), .A2(G169gat), .A3(new_n702), .ZN(new_n946));
  OAI21_X1  g745(.A(G169gat), .B1(new_n945), .B2(new_n566), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1348gat));
  INV_X1    g747(.A(new_n945), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(G176gat), .A3(new_n704), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  AOI21_X1  g752(.A(G176gat), .B1(new_n949), .B2(new_n661), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G1349gat));
  OAI211_X1 g754(.A(new_n949), .B(new_n692), .C1(new_n337), .C2(new_n335), .ZN(new_n956));
  OAI21_X1  g755(.A(G183gat), .B1(new_n945), .B2(new_n691), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(KEYINPUT60), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT60), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n956), .A2(new_n960), .A3(new_n957), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(G1350gat));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n867), .A2(new_n714), .A3(new_n944), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n965), .A3(G190gat), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n965), .B1(new_n964), .B2(G190gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n968), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(KEYINPUT61), .A3(new_n966), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n969), .B(new_n971), .C1(G190gat), .C2(new_n964), .ZN(G1351gat));
  NOR3_X1   g771(.A1(new_n684), .A2(new_n666), .A3(new_n502), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n895), .A2(new_n973), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n974), .A2(G197gat), .A3(new_n702), .ZN(new_n975));
  XOR2_X1   g774(.A(new_n975), .B(KEYINPUT126), .Z(new_n976));
  NAND3_X1  g775(.A1(new_n929), .A2(new_n930), .A3(new_n973), .ZN(new_n977));
  OAI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n566), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1352gat));
  NAND4_X1  g778(.A1(new_n929), .A2(new_n704), .A3(new_n930), .A4(new_n973), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(G204gat), .A3(new_n983), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n974), .A2(G204gat), .A3(new_n662), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n986), .ZN(G1353gat));
  INV_X1    g786(.A(new_n974), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n988), .A2(new_n355), .A3(new_n692), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n929), .A2(new_n692), .A3(new_n930), .A4(new_n973), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT63), .B1(new_n990), .B2(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  NOR3_X1   g792(.A1(new_n977), .A2(new_n356), .A3(new_n640), .ZN(new_n994));
  AOI21_X1  g793(.A(G218gat), .B1(new_n988), .B2(new_n714), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n994), .A2(new_n995), .ZN(G1355gat));
endmodule


