//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G20), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT65), .B(G238), .Z(new_n220));
  OAI221_X1 g0020(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n215), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT66), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT67), .Z(new_n226));
  NAND2_X1  g0026(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n221), .A2(KEYINPUT66), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n210), .B1(new_n213), .B2(new_n217), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT68), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT72), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n248), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n211), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(new_n251), .B2(new_n252), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n202), .B1(new_n248), .B2(G20), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n202), .A2(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n203), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  INV_X1    g0060(.A(G20), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n259), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n214), .A2(KEYINPUT71), .A3(KEYINPUT8), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT8), .B(G58), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT71), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n262), .A2(G20), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n255), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n258), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT70), .A2(G1698), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT70), .A2(G1698), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT3), .B(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(G222), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(G223), .A3(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n278), .B(new_n279), .C1(new_n280), .C2(new_n277), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n212), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(KEYINPUT69), .A2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT69), .A2(G45), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n248), .A2(G274), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G45), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n212), .A2(new_n282), .B1(new_n293), .B2(new_n248), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n291), .B1(G226), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n285), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n273), .B1(new_n297), .B2(G169), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n297), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n285), .A2(G190), .A3(new_n295), .ZN(new_n301));
  XOR2_X1   g0101(.A(new_n301), .B(KEYINPUT74), .Z(new_n302));
  NAND2_X1  g0102(.A1(new_n273), .A2(KEYINPUT9), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(new_n258), .C1(new_n271), .C2(new_n272), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n303), .A2(new_n305), .B1(G200), .B2(new_n296), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n302), .A2(new_n309), .A3(new_n306), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n300), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT70), .ZN(new_n315));
  INV_X1    g0115(.A(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(KEYINPUT70), .A2(G1698), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(G226), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G232), .A2(G1698), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n314), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G97), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n284), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n294), .A2(G238), .B1(new_n289), .B2(new_n290), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n325), .B1(new_n324), .B2(new_n326), .ZN(new_n329));
  OAI21_X1  g0129(.A(G169), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n274), .A2(new_n275), .A3(new_n219), .ZN(new_n333));
  INV_X1    g0133(.A(new_n320), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n277), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n283), .B1(new_n335), .B2(new_n322), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n294), .A2(G238), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n289), .A2(new_n290), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT13), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n327), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n341), .A2(KEYINPUT76), .A3(KEYINPUT14), .A4(G169), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n327), .A2(KEYINPUT75), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT75), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n324), .A2(new_n344), .A3(new_n325), .A4(new_n326), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n329), .A2(new_n299), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n332), .A2(new_n342), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n248), .A2(G20), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n256), .A2(G68), .A3(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n270), .A2(G77), .B1(G20), .B2(new_n215), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n202), .B2(new_n263), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT11), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n352), .A2(new_n353), .A3(new_n255), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(new_n352), .B2(new_n255), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n350), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n251), .A2(new_n252), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(G68), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT12), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n348), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n341), .A2(G200), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n343), .A2(G190), .A3(new_n345), .A4(new_n340), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(new_n360), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n276), .A2(G232), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n366), .B(new_n277), .C1(new_n316), .C2(new_n220), .ZN(new_n367));
  INV_X1    g0167(.A(G107), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n283), .B1(new_n368), .B2(new_n314), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n291), .B1(G244), .B2(new_n294), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT73), .A4(new_n299), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n256), .A2(G77), .A3(new_n349), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT15), .B(G87), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n374), .A2(G20), .A3(new_n262), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n267), .A2(new_n263), .B1(new_n261), .B2(new_n280), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n373), .B1(G77), .B2(new_n357), .C1(new_n377), .C2(new_n272), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(G169), .B1(new_n370), .B2(new_n371), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT73), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n370), .A2(new_n371), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n380), .A2(new_n381), .B1(new_n382), .B2(G179), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n378), .B1(G200), .B2(new_n382), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n370), .A2(new_n371), .A3(G190), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n379), .A2(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n311), .A2(new_n362), .A3(new_n365), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT83), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n291), .B1(G232), .B2(new_n294), .ZN(new_n389));
  INV_X1    g0189(.A(G87), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n262), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n313), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT77), .B(G33), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT3), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n317), .A2(G223), .A3(new_n318), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G226), .A2(G1698), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n391), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT81), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n284), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT77), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(G33), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n262), .A2(KEYINPUT77), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT3), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n406), .A2(KEYINPUT81), .A3(new_n391), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n389), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G169), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT81), .B1(new_n406), .B2(new_n391), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n395), .A2(new_n398), .ZN(new_n412));
  INV_X1    g0212(.A(new_n391), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n400), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(new_n414), .A3(new_n284), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT82), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(new_n299), .A4(new_n389), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n261), .B(new_n392), .C1(new_n393), .C2(new_n394), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT7), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(KEYINPUT78), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n405), .A2(new_n261), .A3(new_n392), .A4(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(G68), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G58), .A2(G68), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(G20), .B1(new_n428), .B2(new_n201), .ZN(new_n429));
  INV_X1    g0229(.A(G159), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(KEYINPUT79), .C1(new_n430), .C2(new_n263), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT79), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n261), .B1(new_n216), .B2(new_n427), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n263), .A2(new_n430), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n426), .A2(new_n436), .A3(KEYINPUT16), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT16), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n431), .A2(new_n435), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n262), .A2(KEYINPUT77), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n402), .A2(G33), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n441), .A3(new_n394), .ZN(new_n442));
  AOI21_X1  g0242(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(KEYINPUT7), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n392), .A2(new_n443), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n421), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n215), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n438), .B1(new_n439), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n437), .A2(new_n255), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n267), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n265), .B1(new_n450), .B2(KEYINPUT71), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n253), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n269), .A2(new_n256), .A3(new_n349), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT80), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT80), .B1(new_n452), .B2(new_n453), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n299), .B(new_n389), .C1(new_n401), .C2(new_n407), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT82), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n418), .A2(new_n419), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n410), .A3(new_n417), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n449), .A2(new_n456), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT18), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G190), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n389), .C1(new_n401), .C2(new_n407), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(G200), .B1(new_n415), .B2(new_n389), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n456), .B(new_n449), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT17), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G200), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n408), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n465), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n462), .A2(new_n473), .A3(KEYINPUT17), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n460), .A2(new_n463), .A3(new_n470), .A4(new_n474), .ZN(new_n475));
  OR3_X1    g0275(.A1(new_n387), .A2(new_n388), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n388), .B1(new_n387), .B2(new_n475), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT86), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n248), .A2(G33), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n481), .B(KEYINPUT84), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n256), .A2(new_n482), .A3(G116), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n253), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n254), .A2(new_n211), .B1(G20), .B2(new_n484), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n261), .C1(G33), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT20), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT20), .B1(new_n487), .B2(new_n490), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n480), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n491), .B(new_n492), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(KEYINPUT86), .A3(new_n483), .A4(new_n485), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n292), .A2(G1), .ZN(new_n500));
  AND2_X1   g0300(.A1(KEYINPUT5), .A2(G41), .ZN(new_n501));
  NOR2_X1   g0301(.A1(KEYINPUT5), .A2(G41), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n503), .A2(new_n283), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G270), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n500), .B(G274), .C1(new_n502), .C2(new_n501), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n395), .A2(G264), .A3(G1698), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n395), .A2(G257), .A3(new_n276), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n314), .A2(G303), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n507), .B1(new_n511), .B2(new_n284), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n499), .A2(G179), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n284), .ZN(new_n514));
  INV_X1    g0314(.A(new_n507), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G200), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n496), .A2(new_n498), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(G190), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n409), .B1(new_n514), .B2(new_n515), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n521), .A2(new_n499), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n521), .B2(new_n499), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n513), .B(new_n520), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n394), .B1(new_n440), .B2(new_n441), .ZN(new_n526));
  OAI211_X1 g0326(.A(G244), .B(new_n276), .C1(new_n526), .C2(new_n313), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT4), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g0329(.A1(KEYINPUT4), .A2(G244), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n276), .A2(new_n277), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n277), .A2(G250), .A3(G1698), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n531), .A2(new_n532), .A3(new_n488), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(new_n284), .B1(G257), .B2(new_n504), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(G179), .A3(new_n506), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n504), .A2(G257), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n531), .A2(new_n532), .A3(new_n488), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n528), .B2(new_n527), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n506), .B(new_n537), .C1(new_n539), .C2(new_n283), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G169), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n443), .A2(KEYINPUT7), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n393), .B2(new_n394), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT7), .B1(new_n392), .B2(new_n443), .ZN(new_n545));
  OAI21_X1  g0345(.A(G107), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT6), .ZN(new_n547));
  AND2_X1   g0347(.A1(G97), .A2(G107), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G97), .A2(G107), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n368), .A2(KEYINPUT6), .A3(G97), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n263), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n552), .A2(G20), .B1(G77), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n272), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n256), .A2(new_n482), .A3(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n253), .A2(new_n489), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n542), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT24), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n261), .A2(G87), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(new_n314), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n440), .A2(new_n441), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n261), .A3(G116), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT23), .B1(new_n261), .B2(G107), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n368), .A3(G20), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n565), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n563), .A2(new_n390), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n261), .B(new_n574), .C1(new_n526), .C2(new_n313), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n562), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n484), .B1(new_n440), .B2(new_n441), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n571), .B1(new_n577), .B2(new_n261), .ZN(new_n578));
  AND4_X1   g0378(.A1(new_n562), .A2(new_n575), .A3(new_n578), .A4(new_n565), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n255), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n503), .A2(new_n283), .A3(G264), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n506), .ZN(new_n582));
  OAI211_X1 g0382(.A(G257), .B(G1698), .C1(new_n526), .C2(new_n313), .ZN(new_n583));
  OAI211_X1 g0383(.A(G250), .B(new_n276), .C1(new_n526), .C2(new_n313), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n566), .A2(G294), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n582), .B1(new_n586), .B2(new_n284), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G190), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n256), .A2(new_n482), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n368), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT25), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n357), .B2(G107), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n590), .A2(G107), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n580), .A2(new_n588), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n587), .A2(new_n471), .ZN(new_n596));
  OR2_X1    g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n374), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n357), .A2(new_n598), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n395), .A2(new_n261), .A3(G68), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT19), .B1(new_n270), .B2(G97), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT19), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n261), .B1(new_n322), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n549), .A2(new_n390), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n599), .B(new_n601), .C1(new_n608), .C2(new_n272), .ZN(new_n609));
  OAI211_X1 g0409(.A(G244), .B(G1698), .C1(new_n526), .C2(new_n313), .ZN(new_n610));
  OAI211_X1 g0410(.A(G238), .B(new_n276), .C1(new_n526), .C2(new_n313), .ZN(new_n611));
  INV_X1    g0411(.A(new_n577), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n284), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n290), .A2(G45), .ZN(new_n615));
  OAI21_X1  g0415(.A(G250), .B1(new_n292), .B2(G1), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n615), .B1(new_n284), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n614), .A2(new_n299), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n613), .B2(new_n284), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n609), .B(new_n619), .C1(G169), .C2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n614), .A2(G190), .A3(new_n618), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n272), .B1(new_n602), .B2(new_n607), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n589), .A2(new_n390), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n623), .A2(new_n624), .A3(new_n600), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n622), .B(new_n625), .C1(new_n471), .C2(new_n620), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n535), .A2(new_n464), .A3(new_n506), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n540), .A2(new_n471), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT85), .B1(new_n555), .B2(new_n558), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n552), .A2(G20), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n553), .A2(G77), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n368), .B1(new_n444), .B2(new_n446), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n255), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n558), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT85), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n631), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n630), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n561), .A2(new_n597), .A3(new_n627), .A4(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n580), .A2(new_n594), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n299), .B(new_n582), .C1(new_n586), .C2(new_n284), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n586), .A2(new_n284), .ZN(new_n645));
  INV_X1    g0445(.A(new_n582), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G169), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT87), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n647), .A2(KEYINPUT87), .A3(G169), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n643), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR4_X1   g0452(.A1(new_n479), .A2(new_n525), .A3(new_n642), .A4(new_n652), .ZN(G372));
  AND3_X1   g0453(.A1(new_n363), .A2(new_n364), .A3(new_n360), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n379), .A2(new_n383), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n470), .B(new_n474), .C1(new_n361), .C2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n460), .A2(new_n463), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n657), .A2(new_n659), .B1(new_n308), .B2(new_n310), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n300), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT88), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n621), .A2(new_n626), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT26), .B1(new_n561), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n640), .B1(new_n541), .B2(new_n536), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n627), .A3(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n664), .A2(new_n667), .A3(new_n621), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n621), .B(new_n626), .C1(new_n595), .C2(new_n596), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n631), .A2(new_n639), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n628), .B2(new_n629), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n559), .B1(new_n536), .B2(new_n541), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n513), .B1(new_n523), .B2(new_n524), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n652), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n478), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n662), .A2(new_n677), .ZN(G369));
  XNOR2_X1  g0478(.A(KEYINPUT90), .B(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n525), .ZN(new_n680));
  INV_X1    g0480(.A(G13), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n681), .A2(G1), .A3(G20), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT89), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n683), .A2(new_n684), .A3(KEYINPUT27), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n683), .B2(KEYINPUT27), .ZN(new_n686));
  OAI221_X1 g0486(.A(G213), .B1(KEYINPUT27), .B2(new_n683), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n680), .B1(new_n518), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n674), .A2(new_n499), .A3(new_n689), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n679), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n580), .A2(new_n594), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n689), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n652), .B1(new_n597), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n649), .B1(new_n587), .B2(new_n409), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n299), .B2(new_n647), .ZN(new_n698));
  INV_X1    g0498(.A(new_n651), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n694), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n689), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n674), .A2(new_n690), .ZN(new_n704));
  OAI22_X1  g0504(.A1(new_n696), .A2(new_n704), .B1(new_n700), .B2(new_n689), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n703), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n208), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n606), .A2(G116), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n709), .A2(new_n248), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n217), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n709), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  AOI21_X1  g0515(.A(new_n689), .B1(new_n668), .B2(new_n675), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n716), .A2(KEYINPUT29), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n523), .A2(new_n524), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT92), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(new_n513), .A4(new_n700), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT92), .B1(new_n674), .B2(new_n652), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(new_n673), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n627), .A2(new_n666), .A3(new_n672), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n621), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n666), .B1(new_n665), .B2(new_n627), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n689), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT29), .ZN(new_n728));
  INV_X1    g0528(.A(new_n679), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n690), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n535), .A2(new_n620), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(KEYINPUT30), .A3(new_n512), .A4(new_n644), .ZN(new_n733));
  AOI21_X1  g0533(.A(G179), .B1(new_n614), .B2(new_n618), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n734), .A2(new_n516), .A3(new_n647), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n644), .A2(new_n535), .A3(new_n512), .A4(new_n620), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n735), .A2(new_n540), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT91), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n733), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n736), .A2(new_n737), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n540), .A2(new_n734), .A3(new_n516), .A4(new_n647), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n741), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n731), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n673), .A2(new_n680), .A3(new_n700), .A4(new_n690), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n733), .A2(new_n741), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n689), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n730), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n744), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n717), .A2(new_n728), .B1(new_n729), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n715), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(new_n709), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n681), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n248), .B1(new_n753), .B2(G45), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n693), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n691), .A2(new_n679), .A3(new_n692), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n691), .A2(new_n692), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n708), .A2(new_n314), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G355), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G116), .B2(new_n208), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n708), .A2(new_n395), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n286), .A2(new_n288), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n768), .B1(new_n713), .B2(new_n770), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n243), .A2(new_n292), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n766), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n211), .B1(G20), .B2(new_n409), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n762), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n756), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n261), .A2(G179), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT94), .Z(new_n780));
  NAND3_X1  g0580(.A1(new_n299), .A2(new_n471), .A3(KEYINPUT93), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT93), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(G179), .B2(G200), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n464), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n261), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n780), .A2(G303), .B1(new_n786), .B2(G294), .ZN(new_n787));
  NAND2_X1  g0587(.A1(G20), .A2(G179), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n788), .A2(G190), .A3(G200), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n314), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n778), .A2(new_n464), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n792), .B1(G283), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(G20), .A2(G179), .A3(G190), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n471), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n797), .A2(G322), .B1(new_n798), .B2(G326), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n788), .A2(new_n471), .A3(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n801), .B1(KEYINPUT95), .B2(new_n803), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n803), .A2(KEYINPUT95), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n261), .B(G190), .C1(new_n781), .C2(new_n783), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(G329), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n787), .A2(new_n795), .A3(new_n799), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(G159), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT32), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n277), .B1(new_n790), .B2(new_n280), .C1(new_n215), .C2(new_n801), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n793), .A2(new_n368), .B1(new_n779), .B2(new_n390), .ZN(new_n812));
  INV_X1    g0612(.A(new_n798), .ZN(new_n813));
  INV_X1    g0613(.A(new_n797), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n202), .A2(new_n813), .B1(new_n814), .B2(new_n214), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n811), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n489), .B2(new_n785), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n808), .B1(new_n810), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n777), .B1(new_n818), .B2(new_n774), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n763), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n759), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n689), .A2(new_n378), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n377), .A2(new_n272), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n280), .B2(new_n253), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n382), .A2(G200), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n826), .A2(new_n827), .A3(new_n373), .A4(new_n385), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n824), .B1(new_n655), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n823), .B1(new_n379), .B2(new_n383), .ZN(new_n830));
  OAI21_X1  g0630(.A(KEYINPUT100), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n830), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT100), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(new_n386), .C2(new_n824), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n716), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n749), .A2(new_n729), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n756), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  INV_X1    g0639(.A(new_n774), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n761), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n756), .B1(G77), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT96), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G150), .A2(new_n800), .B1(new_n789), .B2(G159), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n797), .A2(G143), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n813), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT34), .Z(new_n848));
  OAI21_X1  g0648(.A(new_n395), .B1(new_n215), .B2(new_n793), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G132), .B2(new_n806), .ZN(new_n850));
  INV_X1    g0650(.A(new_n780), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n214), .B2(new_n785), .C1(new_n851), .C2(new_n202), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n848), .B1(new_n852), .B2(KEYINPUT98), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n852), .A2(KEYINPUT98), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G116), .A2(new_n789), .B1(new_n800), .B2(G283), .ZN(new_n855));
  INV_X1    g0655(.A(G303), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n855), .B1(new_n813), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT97), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n851), .A2(new_n368), .B1(new_n489), .B2(new_n785), .ZN(new_n859));
  INV_X1    g0659(.A(new_n806), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(new_n791), .ZN(new_n861));
  INV_X1    g0661(.A(G294), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n314), .B1(new_n793), .B2(new_n390), .C1(new_n862), .C2(new_n814), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n859), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n853), .A2(new_n854), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n843), .B1(new_n865), .B2(new_n840), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT99), .Z(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n761), .B2(new_n835), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n839), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(G384));
  AOI211_X1 g0670(.A(new_n484), .B(new_n213), .C1(new_n552), .C2(KEYINPUT35), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(KEYINPUT35), .B2(new_n552), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT36), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n427), .A2(G77), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n217), .A2(new_n874), .B1(G50), .B2(new_n215), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(G1), .A3(new_n681), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT101), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n437), .A2(new_n255), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT16), .B1(new_n426), .B2(new_n436), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n456), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT103), .ZN(new_n883));
  INV_X1    g0683(.A(new_n687), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT103), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n885), .B(new_n456), .C1(new_n880), .C2(new_n881), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n883), .A2(new_n886), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n887), .B(new_n468), .C1(new_n888), .C2(new_n461), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n457), .A2(new_n459), .A3(new_n410), .A4(new_n417), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT104), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n687), .B1(new_n449), .B2(new_n456), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n468), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n890), .A2(new_n891), .ZN(new_n898));
  AOI22_X1  g0698(.A1(KEYINPUT37), .A2(new_n889), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n887), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n475), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n879), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n418), .A2(KEYINPUT104), .A3(new_n457), .A4(new_n459), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n893), .B1(new_n473), .B2(new_n462), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n905), .A2(new_n898), .A3(new_n895), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n746), .A2(new_n731), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n745), .A2(new_n748), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n360), .A2(new_n690), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n365), .B(new_n914), .C1(new_n348), .C2(new_n360), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT102), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n347), .A2(new_n343), .A3(new_n345), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n341), .A2(G169), .B1(KEYINPUT76), .B2(KEYINPUT14), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n409), .B(new_n331), .C1(new_n340), .C2(new_n327), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n916), .B(new_n913), .C1(new_n920), .C2(new_n654), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n348), .A2(new_n365), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n916), .B1(new_n923), .B2(new_n913), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n835), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT106), .B1(new_n912), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n831), .A2(new_n834), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n915), .A2(new_n921), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n923), .A2(new_n913), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT102), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n927), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT106), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n745), .A2(new_n748), .A3(new_n911), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n910), .A2(new_n926), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n931), .A2(KEYINPUT40), .A3(new_n933), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n470), .A2(new_n474), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n893), .B1(new_n658), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n906), .A2(new_n890), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT37), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n940), .A2(KEYINPUT105), .B1(new_n907), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT105), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n475), .A2(new_n944), .A3(new_n893), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT38), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n899), .A2(new_n902), .A3(new_n879), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n938), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n937), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n479), .A2(new_n912), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n729), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n655), .A2(new_n689), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n716), .B2(new_n835), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n922), .A2(new_n924), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n957), .A2(new_n910), .B1(new_n658), .B2(new_n687), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT39), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n946), .B2(new_n947), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n362), .A2(new_n689), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n903), .A2(new_n909), .A3(KEYINPUT39), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n478), .A2(new_n717), .A3(new_n728), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n662), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n964), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n953), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n248), .B2(new_n753), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n953), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n878), .B1(new_n969), .B2(new_n970), .ZN(G367));
  INV_X1    g0771(.A(new_n704), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n561), .B(new_n641), .C1(new_n640), .C2(new_n690), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n665), .A2(new_n689), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n702), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT42), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT42), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n672), .B1(new_n975), .B2(new_n652), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n977), .B(new_n978), .C1(new_n689), .C2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n690), .A2(new_n625), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT107), .Z(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n627), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n621), .B2(new_n982), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n980), .A2(KEYINPUT43), .A3(new_n984), .ZN(new_n989));
  INV_X1    g0789(.A(new_n703), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n975), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n988), .A2(new_n989), .B1(KEYINPUT108), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(KEYINPUT108), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n709), .B(KEYINPUT41), .Z(new_n996));
  XNOR2_X1  g0796(.A(new_n702), .B(new_n972), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(new_n693), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n750), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(KEYINPUT110), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT110), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n975), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n705), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n705), .A2(new_n1004), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n703), .B1(new_n1011), .B2(KEYINPUT109), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT109), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1010), .A2(new_n1013), .A3(new_n990), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1001), .A2(new_n1003), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n996), .B1(new_n1015), .B2(new_n750), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n754), .B(KEYINPUT111), .Z(new_n1017));
  OAI211_X1 g0817(.A(new_n994), .B(new_n995), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n235), .A2(new_n768), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n775), .B1(new_n208), .B2(new_n374), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n756), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n277), .B1(new_n790), .B2(new_n202), .C1(new_n430), .C2(new_n801), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G137), .B2(new_n806), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n793), .A2(new_n280), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n814), .A2(new_n260), .B1(new_n779), .B2(new_n214), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G143), .C2(new_n798), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1023), .B(new_n1026), .C1(new_n215), .C2(new_n785), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT113), .Z(new_n1028));
  NAND3_X1  g0828(.A1(new_n780), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT112), .ZN(new_n1030));
  INV_X1    g0830(.A(G317), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n860), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n779), .ZN(new_n1033));
  AOI21_X1  g0833(.A(KEYINPUT46), .B1(new_n1033), .B2(G116), .ZN(new_n1034));
  INV_X1    g0834(.A(G283), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n801), .A2(new_n862), .B1(new_n790), .B2(new_n1035), .ZN(new_n1036));
  NOR4_X1   g0836(.A1(new_n1032), .A2(new_n395), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n793), .A2(new_n489), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G311), .B2(new_n798), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n856), .B2(new_n814), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G107), .B2(new_n786), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1030), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1028), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT47), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1021), .B1(new_n1044), .B2(new_n774), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n762), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1045), .B1(new_n1046), .B2(new_n984), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1018), .A2(new_n1047), .ZN(G387));
  NOR2_X1   g0848(.A1(new_n702), .A2(new_n1046), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n764), .A2(new_n711), .B1(new_n368), .B2(new_n708), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n450), .A2(new_n202), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT50), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  AOI211_X1 g0853(.A(G45), .B(new_n711), .C1(G68), .C2(G77), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n768), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(KEYINPUT114), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT114), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1055), .A2(new_n1058), .B1(new_n239), .B2(new_n770), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1050), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n776), .B1(new_n1060), .B2(KEYINPUT115), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(KEYINPUT115), .B2(new_n1060), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n756), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1033), .A2(G77), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n813), .B2(new_n430), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1038), .B(new_n1065), .C1(G50), .C2(new_n797), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n806), .A2(G150), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n395), .B1(new_n215), .B2(new_n790), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n269), .B2(new_n800), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n786), .A2(new_n598), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n806), .A2(G326), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n395), .B1(G116), .B2(new_n794), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G303), .A2(new_n789), .B1(new_n800), .B2(G311), .ZN(new_n1074));
  INV_X1    g0874(.A(G322), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1074), .B1(new_n814), .B2(new_n1031), .C1(new_n1075), .C2(new_n813), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n1035), .B2(new_n785), .C1(new_n862), .C2(new_n779), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT116), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT49), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1072), .B(new_n1073), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1071), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1049), .B(new_n1063), .C1(new_n774), .C2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n998), .B2(new_n1017), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n999), .A2(new_n709), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n998), .A2(new_n750), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(G393));
  INV_X1    g0891(.A(KEYINPUT117), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1011), .A2(new_n1092), .A3(new_n703), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT117), .B1(new_n1010), .B2(new_n990), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1010), .A2(new_n990), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1015), .B(new_n709), .C1(new_n1096), .C2(new_n1000), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1004), .A2(new_n762), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n768), .A2(new_n246), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n775), .B1(new_n208), .B2(new_n489), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n756), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n314), .B1(new_n790), .B2(new_n862), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n793), .A2(new_n368), .B1(new_n779), .B2(new_n1035), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(G303), .C2(new_n800), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n484), .B2(new_n785), .C1(new_n1075), .C2(new_n860), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n797), .A2(G311), .B1(new_n798), .B2(G317), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT52), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1033), .A2(G68), .B1(new_n794), .B2(G87), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n806), .A2(G143), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n450), .A2(new_n789), .B1(new_n800), .B2(G50), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1108), .A2(new_n395), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n786), .A2(G77), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n797), .A2(G159), .B1(new_n798), .B2(G150), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1113), .A2(KEYINPUT51), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(KEYINPUT51), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1105), .A2(new_n1107), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1101), .B1(new_n1117), .B2(new_n774), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1096), .A2(new_n1017), .B1(new_n1098), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1097), .A2(new_n1119), .ZN(G390));
  INV_X1    g0920(.A(new_n961), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n955), .B2(new_n956), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n940), .A2(KEYINPUT105), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n942), .A2(new_n907), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n945), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n879), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT39), .B1(new_n1126), .B2(new_n909), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n903), .A2(new_n909), .A3(KEYINPUT39), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n909), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n954), .B1(new_n727), .B2(new_n835), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1130), .B(new_n1121), .C1(new_n956), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n956), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1133), .A2(new_n749), .A3(new_n729), .A4(new_n835), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1129), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n931), .A2(G330), .A3(new_n933), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n933), .A2(G330), .A3(new_n835), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n956), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT118), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n912), .A2(new_n925), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n749), .A2(new_n729), .A3(new_n835), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1143), .A2(G330), .B1(new_n1144), .B2(new_n956), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1142), .B1(new_n1145), .B2(new_n955), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n956), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1136), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n674), .A2(new_n652), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1149), .A2(new_n642), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n664), .A2(new_n667), .A3(new_n621), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n835), .B(new_n690), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n954), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1148), .A2(KEYINPUT118), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1141), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n478), .A2(G330), .A3(new_n933), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n965), .A2(new_n1157), .A3(new_n662), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1135), .A2(new_n1137), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT118), .B1(new_n1148), .B2(new_n1154), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1142), .B(new_n955), .C1(new_n1147), .C2(new_n1136), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1140), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1136), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n961), .B1(new_n1154), .B2(new_n1133), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n960), .B2(new_n962), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1121), .B1(new_n946), .B2(new_n947), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n727), .A2(new_n835), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n956), .B1(new_n1167), .B2(new_n1153), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1163), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1129), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n965), .A2(new_n1157), .A3(new_n662), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1162), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1159), .A2(new_n709), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1170), .A2(new_n1171), .A3(new_n1017), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n760), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n756), .B1(new_n269), .B2(new_n841), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n314), .B1(new_n790), .B2(new_n489), .C1(new_n368), .C2(new_n801), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G294), .B2(new_n806), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n814), .A2(new_n484), .B1(new_n793), .B2(new_n215), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G283), .B2(new_n798), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n780), .A2(G87), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1112), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n806), .A2(G125), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1033), .A2(G150), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1184), .B1(KEYINPUT53), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(KEYINPUT53), .B2(new_n1185), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT54), .B(G143), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n277), .B1(new_n790), .B2(new_n1188), .C1(new_n846), .C2(new_n801), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G50), .B2(new_n794), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1187), .B(new_n1190), .C1(new_n430), .C2(new_n785), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n797), .A2(G132), .B1(new_n798), .B2(G128), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT119), .Z(new_n1193));
  OAI21_X1  g0993(.A(new_n1183), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1177), .B1(new_n1194), .B2(new_n774), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1176), .A2(new_n1195), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1175), .A2(new_n1196), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1174), .A2(KEYINPUT120), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT120), .B1(new_n1174), .B2(new_n1197), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(G378));
  NAND2_X1  g1000(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1172), .B1(new_n1201), .B2(new_n1156), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT122), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT122), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1173), .A2(new_n1204), .A3(new_n1172), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n964), .ZN(new_n1207));
  INV_X1    g1007(.A(G330), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1130), .B2(new_n938), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n884), .A2(new_n273), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n311), .B(new_n1210), .Z(new_n1211));
  XNOR2_X1  g1011(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1211), .B(new_n1212), .Z(new_n1213));
  AND3_X1   g1013(.A1(new_n937), .A2(new_n1209), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n937), .B2(new_n1209), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1207), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1211), .B(new_n1212), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n931), .A2(new_n933), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(KEYINPUT106), .A2(new_n1218), .B1(new_n903), .B2(new_n909), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT40), .B1(new_n1219), .B2(new_n934), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n948), .A2(G330), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1217), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n937), .A2(new_n1209), .A3(new_n1213), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n964), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1216), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT57), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1222), .A2(new_n964), .A3(new_n1223), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n964), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT123), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT123), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1216), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1228), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n752), .B1(new_n1234), .B2(new_n1206), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1017), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1216), .B2(new_n1224), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n756), .B1(G50), .B2(new_n841), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1217), .A2(new_n761), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n395), .A2(G41), .ZN(new_n1240));
  AOI211_X1 g1040(.A(G50), .B(new_n1240), .C1(new_n262), .C2(new_n287), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n793), .A2(new_n214), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n368), .A2(new_n814), .B1(new_n813), .B2(new_n484), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(G68), .C2(new_n786), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1064), .B1(new_n489), .B2(new_n801), .C1(new_n374), .C2(new_n790), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1240), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1244), .B(new_n1247), .C1(new_n1035), .C2(new_n860), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT58), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1241), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(G132), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n801), .A2(new_n1251), .B1(new_n790), .B2(new_n846), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1188), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(new_n1033), .B2(new_n1253), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n797), .A2(G128), .B1(new_n798), .B2(G125), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1254), .B(new_n1255), .C1(new_n260), .C2(new_n785), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(KEYINPUT59), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(KEYINPUT59), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n262), .B(new_n287), .C1(new_n793), .C2(new_n430), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G124), .B2(new_n806), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n1250), .B1(new_n1249), .B2(new_n1248), .C1(new_n1257), .C2(new_n1261), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1238), .B(new_n1239), .C1(new_n774), .C2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT121), .B1(new_n1237), .B2(new_n1263), .ZN(new_n1264));
  OR3_X1    g1064(.A1(new_n1237), .A2(KEYINPUT121), .A3(new_n1263), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1227), .A2(new_n1235), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(G375));
  NAND2_X1  g1067(.A1(new_n956), .A2(new_n760), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n756), .B1(G68), .B2(new_n841), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n813), .A2(new_n1251), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1242), .B(new_n1270), .C1(G137), .C2(new_n797), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n806), .A2(G128), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1253), .A2(new_n800), .B1(new_n789), .B2(G150), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1271), .A2(new_n395), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n851), .A2(new_n430), .B1(new_n202), .B2(new_n785), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1070), .B1(new_n851), .B2(new_n489), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n314), .B1(new_n801), .B2(new_n484), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(G107), .B2(new_n789), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n797), .A2(G283), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1024), .B1(G294), .B2(new_n798), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n806), .A2(G303), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n1274), .A2(new_n1275), .B1(new_n1276), .B2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1269), .B1(new_n1283), .B2(new_n774), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1162), .A2(new_n1017), .B1(new_n1268), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1162), .A2(new_n1172), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n996), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1162), .A2(new_n1172), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1285), .B1(new_n1288), .B2(new_n1289), .ZN(G381));
  AND2_X1   g1090(.A1(new_n1174), .A2(new_n1197), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1266), .A2(new_n1291), .ZN(new_n1292));
  OR2_X1    g1092(.A1(G393), .A2(G396), .ZN(new_n1293));
  OR4_X1    g1093(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1293), .ZN(new_n1294));
  OR3_X1    g1094(.A1(new_n1292), .A2(new_n1294), .A3(G381), .ZN(G407));
  OAI211_X1 g1095(.A(G407), .B(G213), .C1(G343), .C2(new_n1292), .ZN(G409));
  AOI21_X1  g1096(.A(new_n996), .B1(new_n1216), .B2(new_n1224), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1173), .A2(new_n1204), .A3(new_n1172), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1204), .B1(new_n1173), .B2(new_n1172), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT124), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT124), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1206), .A2(new_n1302), .A3(new_n1297), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1263), .B1(new_n1304), .B2(new_n1017), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1301), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1291), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1265), .A2(new_n1264), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1232), .B1(new_n1216), .B2(new_n1224), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1230), .A2(KEYINPUT123), .ZN(new_n1311));
  OAI21_X1  g1111(.A(KEYINPUT57), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n709), .B1(new_n1309), .B2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G378), .B(new_n1308), .C1(new_n1313), .C2(new_n1226), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1307), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n688), .A2(G213), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1289), .B1(KEYINPUT60), .B2(new_n1286), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1156), .A2(KEYINPUT60), .A3(new_n1158), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n709), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1285), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  OR2_X1    g1120(.A1(new_n1320), .A2(new_n869), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n869), .ZN(new_n1322));
  AND2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1315), .A2(new_n1316), .A3(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT126), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1325), .A3(KEYINPUT62), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1316), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(G2897), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1321), .A2(new_n1322), .A3(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1329), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT61), .B1(new_n1327), .B2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1328), .B1(new_n1307), .B2(new_n1314), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(new_n1323), .A3(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1326), .A2(new_n1333), .A3(new_n1336), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(G393), .B(new_n821), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1018), .A2(G390), .A3(new_n1047), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(G390), .B1(new_n1018), .B2(new_n1047), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1339), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1342), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1344), .A2(new_n1338), .A3(new_n1340), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1337), .A2(new_n1346), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1321), .A2(KEYINPUT63), .A3(new_n1322), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1315), .A2(new_n1316), .A3(new_n1348), .ZN(new_n1349));
  AND2_X1   g1149(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(KEYINPUT63), .B1(new_n1334), .B2(new_n1323), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(KEYINPUT125), .B1(new_n1353), .B2(new_n1333), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT63), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1324), .A2(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1346), .B1(new_n1334), .B2(new_n1348), .ZN(new_n1357));
  AND4_X1   g1157(.A1(KEYINPUT125), .A2(new_n1333), .A3(new_n1356), .A4(new_n1357), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1347), .B1(new_n1354), .B2(new_n1358), .ZN(G405));
  INV_X1    g1159(.A(new_n1291), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1314), .B1(new_n1266), .B2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(KEYINPUT127), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1323), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT127), .ZN(new_n1364));
  OAI211_X1 g1164(.A(new_n1364), .B(new_n1314), .C1(new_n1266), .C2(new_n1360), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1362), .A2(new_n1363), .A3(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1366), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1363), .B1(new_n1362), .B2(new_n1365), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1346), .B1(new_n1367), .B2(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1368), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1370), .A2(new_n1350), .A3(new_n1366), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1369), .A2(new_n1371), .ZN(G402));
endmodule


