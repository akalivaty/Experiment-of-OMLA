//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n865, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(KEYINPUT78), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(KEYINPUT78), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n211), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n213), .A2(new_n208), .A3(new_n207), .A4(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT79), .B(KEYINPUT29), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G226gat), .A2(G233gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  AND2_X1   g020(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT70), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(KEYINPUT28), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI221_X1 g026(.A(new_n221), .B1(new_n225), .B2(KEYINPUT28), .C1(new_n222), .C2(new_n223), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(G169gat), .ZN(new_n231));
  INV_X1    g030(.A(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT71), .B1(new_n233), .B2(KEYINPUT26), .ZN(new_n234));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT68), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(G169gat), .A3(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(KEYINPUT26), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n231), .A4(new_n232), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n234), .A2(new_n239), .A3(new_n240), .A4(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n230), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT72), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT72), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n229), .A2(new_n247), .A3(new_n244), .A4(new_n230), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT23), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(G176gat), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n252), .B2(new_n231), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT24), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n230), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n256));
  INV_X1    g055(.A(G183gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n221), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n260));
  NAND2_X1  g059(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n233), .A3(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n253), .A2(new_n259), .A3(new_n262), .A4(new_n239), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT69), .ZN(new_n264));
  AND2_X1   g063(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n265));
  NOR2_X1   g064(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n267), .A2(new_n233), .B1(new_n236), .B2(new_n238), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n268), .A2(new_n269), .A3(new_n253), .A4(new_n259), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n273), .A2(new_n255), .A3(new_n258), .A4(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n231), .A2(KEYINPUT66), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n231), .A2(KEYINPUT66), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n252), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n268), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n271), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n220), .B1(new_n249), .B2(new_n282), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n264), .A2(new_n270), .B1(new_n279), .B2(new_n280), .ZN(new_n284));
  INV_X1    g083(.A(new_n245), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n284), .A2(new_n285), .A3(new_n219), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n216), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n249), .A2(G226gat), .A3(new_n282), .A4(G233gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n289), .B(new_n219), .C1(new_n284), .C2(new_n285), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n290), .A3(new_n215), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT37), .ZN(new_n293));
  AOI211_X1 g092(.A(KEYINPUT38), .B(new_n205), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n215), .B1(new_n283), .B2(new_n286), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT91), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n288), .A2(new_n216), .A3(new_n290), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT91), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n298), .B(new_n215), .C1(new_n283), .C2(new_n286), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT37), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303));
  INV_X1    g102(.A(G155gat), .ZN(new_n304));
  INV_X1    g103(.A(G162gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  INV_X1    g106(.A(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G141gat), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G148gat), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n306), .A2(new_n307), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n310), .A2(G148gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n308), .A2(G141gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n303), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G155gat), .B(G162gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT81), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT2), .B1(new_n309), .B2(new_n311), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT81), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n320), .A2(new_n321), .A3(new_n317), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n313), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(KEYINPUT82), .A3(KEYINPUT3), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT81), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n321), .B1(new_n320), .B2(new_n317), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n312), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G127gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G134gat), .ZN(new_n332));
  INV_X1    g131(.A(G134gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G127gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(KEYINPUT73), .A3(G134gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G113gat), .B(G120gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n336), .B(new_n337), .C1(KEYINPUT1), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n338), .ZN(new_n340));
  XOR2_X1   g139(.A(KEYINPUT74), .B(KEYINPUT1), .Z(new_n341));
  XNOR2_X1  g140(.A(G127gat), .B(G134gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n329), .B(new_n313), .C1(new_n319), .C2(new_n322), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n324), .A2(new_n330), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n339), .B2(new_n343), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n328), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(KEYINPUT5), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n328), .A2(KEYINPUT4), .A3(new_n339), .A4(new_n343), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n346), .A2(new_n352), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  OAI22_X1  g156(.A1(new_n323), .A2(new_n344), .B1(new_n351), .B2(new_n354), .ZN(new_n358));
  OAI211_X1 g157(.A(KEYINPUT4), .B(new_n328), .C1(new_n347), .C2(new_n349), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n346), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n328), .B(new_n344), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT5), .B1(new_n362), .B2(new_n353), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n357), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(G57gat), .B(G85gat), .Z(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n369), .B(KEYINPUT90), .Z(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n357), .B(new_n369), .C1(new_n361), .C2(new_n363), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n369), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n364), .A2(KEYINPUT6), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n292), .A2(new_n205), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n302), .A2(new_n375), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n287), .A2(new_n380), .A3(new_n291), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n287), .B2(new_n291), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT37), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n205), .B1(new_n292), .B2(new_n293), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT92), .B1(new_n385), .B2(KEYINPUT38), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT38), .ZN(new_n388));
  AOI211_X1 g187(.A(new_n387), .B(new_n388), .C1(new_n383), .C2(new_n384), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n379), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT85), .B(G50gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G78gat), .B(G106gat), .Z(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G228gat), .ZN(new_n396));
  INV_X1    g195(.A(G233gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n323), .A2(new_n215), .A3(new_n218), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT86), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n323), .A2(KEYINPUT3), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n399), .B2(new_n401), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n217), .B1(new_n328), .B2(new_n329), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT87), .B1(new_n405), .B2(new_n215), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n345), .A2(new_n218), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT87), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n216), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n398), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT3), .B1(new_n215), .B2(new_n289), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(new_n328), .ZN(new_n413));
  INV_X1    g212(.A(new_n398), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT88), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n407), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n405), .A2(KEYINPUT88), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(new_n216), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n411), .A2(G22gat), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G22gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n399), .A2(new_n401), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT86), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n424), .A2(new_n409), .A3(new_n406), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n414), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n415), .A2(new_n419), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n422), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n395), .B1(new_n421), .B2(new_n429), .ZN(new_n430));
  AND4_X1   g229(.A1(KEYINPUT89), .A2(new_n427), .A3(new_n422), .A4(new_n428), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(G22gat), .B1(new_n411), .B2(new_n420), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n427), .A2(new_n422), .A3(new_n428), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n395), .A2(KEYINPUT89), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n430), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n360), .B(KEYINPUT5), .C1(new_n353), .C2(new_n362), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n370), .B1(new_n439), .B2(new_n357), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n346), .A2(new_n352), .A3(new_n356), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n354), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n362), .A2(new_n353), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(KEYINPUT39), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT39), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n445), .A3(new_n354), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n370), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT40), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n440), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n204), .B1(new_n381), .B2(new_n382), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(KEYINPUT30), .A3(new_n378), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n378), .A2(KEYINPUT30), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n444), .A2(KEYINPUT40), .A3(new_n370), .A4(new_n446), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n449), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT93), .B1(new_n390), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n374), .A2(new_n373), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n369), .B1(new_n439), .B2(new_n357), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n377), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n451), .A2(new_n452), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n433), .A2(new_n434), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n431), .B1(new_n461), .B2(new_n395), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n459), .A2(new_n460), .B1(new_n462), .B2(new_n436), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT36), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT77), .B(KEYINPUT34), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n249), .A2(new_n282), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n347), .A2(new_n349), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT76), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  INV_X1    g268(.A(new_n467), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT76), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n470), .A2(new_n249), .A3(new_n471), .A4(new_n282), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G227gat), .A2(G233gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT33), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G15gat), .B(G43gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(G71gat), .B(G99gat), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n477), .B(new_n478), .Z(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n465), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n473), .A2(new_n475), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n468), .A2(new_n472), .A3(new_n474), .A4(new_n469), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(KEYINPUT32), .A3(new_n484), .ZN(new_n485));
  OR3_X1    g284(.A1(new_n473), .A2(KEYINPUT32), .A3(new_n475), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n476), .A2(new_n465), .A3(new_n480), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n482), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n476), .ZN(new_n490));
  INV_X1    g289(.A(new_n465), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(new_n479), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n492), .A2(new_n481), .B1(new_n486), .B2(new_n485), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n464), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n487), .B1(new_n482), .B2(new_n488), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n492), .A2(new_n481), .A3(new_n486), .A4(new_n485), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(KEYINPUT36), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n463), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n377), .B1(new_n457), .B2(new_n440), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n301), .B2(new_n294), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n292), .A2(KEYINPUT80), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n287), .A2(new_n380), .A3(new_n291), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n293), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n384), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT38), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n387), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n385), .A2(KEYINPUT92), .A3(KEYINPUT38), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n500), .A2(new_n506), .A3(new_n378), .A4(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n451), .A2(new_n452), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n447), .A2(new_n448), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n510), .A2(new_n372), .A3(new_n453), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n437), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n508), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n456), .A2(new_n498), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n489), .A2(new_n493), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n460), .A2(new_n499), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n438), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n489), .A2(new_n493), .A3(new_n437), .ZN(new_n520));
  INV_X1    g319(.A(new_n459), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n509), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G57gat), .B(G64gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT99), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT9), .ZN(new_n527));
  XOR2_X1   g326(.A(G71gat), .B(G78gat), .Z(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G71gat), .ZN(new_n530));
  INV_X1    g329(.A(G78gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT9), .ZN(new_n532));
  NAND2_X1  g331(.A1(G71gat), .A2(G78gat), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(new_n525), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT100), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n529), .A2(KEYINPUT100), .A3(new_n536), .ZN(new_n540));
  NAND2_X1  g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  INV_X1    g341(.A(G99gat), .ZN(new_n543));
  INV_X1    g342(.A(G106gat), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT8), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n542), .B(new_n545), .C1(G85gat), .C2(G92gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(G99gat), .B(G106gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n539), .A2(new_n540), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT10), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n547), .A2(KEYINPUT105), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n546), .B(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n537), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n556), .A2(KEYINPUT106), .A3(KEYINPUT10), .A4(new_n548), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT100), .B1(new_n529), .B2(new_n536), .ZN(new_n558));
  AOI211_X1 g357(.A(new_n538), .B(new_n535), .C1(new_n527), .C2(new_n528), .ZN(new_n559));
  OAI211_X1 g358(.A(KEYINPUT10), .B(new_n548), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT106), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G230gat), .A2(G233gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n554), .ZN(new_n566));
  INV_X1    g365(.A(new_n564), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT107), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT107), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n565), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G120gat), .B(G148gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n565), .A2(new_n577), .A3(new_n569), .A4(new_n571), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT108), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT109), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n578), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n576), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n579), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT109), .ZN(new_n585));
  INV_X1    g384(.A(new_n576), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G1gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(G15gat), .B(G22gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n592), .B2(KEYINPUT96), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT96), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n594), .A3(G1gat), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n593), .B(new_n595), .C1(KEYINPUT16), .C2(new_n592), .ZN(new_n596));
  INV_X1    g395(.A(G8gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n591), .A2(G1gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(KEYINPUT97), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n596), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G43gat), .B(G50gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT15), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(G29gat), .ZN(new_n604));
  INV_X1    g403(.A(G36gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT14), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT14), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(G29gat), .B2(G36gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g410(.A1(G29gat), .A2(G36gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n612), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n603), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n601), .A2(KEYINPUT15), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n616), .A2(new_n610), .A3(new_n602), .A4(new_n612), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n618), .B(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n619), .B(new_n620), .C1(new_n622), .C2(new_n600), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n618), .B(KEYINPUT17), .ZN(new_n626));
  INV_X1    g425(.A(new_n600), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n628), .A2(KEYINPUT18), .A3(new_n619), .A4(new_n620), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n620), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n619), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n600), .A2(new_n618), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n625), .A2(new_n629), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G113gat), .B(G141gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G197gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT11), .B(G169gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XOR2_X1   g439(.A(new_n640), .B(KEYINPUT94), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n625), .A2(new_n629), .A3(new_n640), .A4(new_n634), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n589), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G183gat), .B(G211gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(new_n331), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n600), .B1(new_n556), .B2(KEYINPUT21), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n558), .A2(new_n559), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT21), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(G231gat), .A2(G233gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n652), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n655), .A2(new_n656), .ZN(new_n661));
  INV_X1    g460(.A(new_n652), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(new_n657), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n660), .B2(new_n663), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n651), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n667), .ZN(new_n669));
  INV_X1    g468(.A(new_n651), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n665), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G155gat), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G190gat), .B(G218gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(new_n305), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n626), .A2(new_n549), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n548), .A2(new_n618), .ZN(new_n683));
  NAND3_X1  g482(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G134gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n682), .A2(new_n333), .A3(new_n683), .A4(new_n684), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n686), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n690), .B1(new_n686), .B2(new_n691), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n681), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n694), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(new_n680), .A3(new_n692), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n678), .A2(new_n699), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n524), .A2(new_n649), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n521), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G1gat), .ZN(G1324gat));
  NAND4_X1  g502(.A1(new_n524), .A2(new_n649), .A3(new_n700), .A4(new_n509), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT16), .B(G8gat), .ZN(new_n706));
  OR3_X1    g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n704), .B(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n705), .B1(new_n709), .B2(G8gat), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n706), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT111), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n707), .B(new_n714), .C1(new_n710), .C2(new_n711), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1325gat));
  AOI21_X1  g515(.A(G15gat), .B1(new_n701), .B2(new_n516), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n494), .A2(new_n497), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n719), .A2(G15gat), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n717), .B1(new_n701), .B2(new_n720), .ZN(G1326gat));
  NAND2_X1  g520(.A1(new_n701), .A2(new_n437), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT43), .B(G22gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1327gat));
  NAND2_X1  g523(.A1(new_n524), .A2(new_n699), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n649), .A2(new_n678), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n604), .A3(new_n521), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n725), .A2(KEYINPUT113), .A3(KEYINPUT44), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n698), .B1(new_n515), .B2(new_n523), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n695), .A2(new_n697), .A3(KEYINPUT115), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT115), .B1(new_n695), .B2(new_n697), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n515), .A2(new_n740), .A3(new_n523), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n515), .B2(new_n523), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n734), .B(new_n739), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n459), .B(new_n726), .C1(new_n736), .C2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n730), .B1(new_n744), .B2(new_n604), .ZN(G1328gat));
  NAND3_X1  g544(.A1(new_n727), .A2(new_n605), .A3(new_n509), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT46), .Z(new_n747));
  AOI211_X1 g546(.A(new_n460), .B(new_n726), .C1(new_n736), .C2(new_n743), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n605), .ZN(G1329gat));
  AOI21_X1  g548(.A(KEYINPUT113), .B1(new_n725), .B2(KEYINPUT44), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n733), .A2(new_n732), .A3(new_n734), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n743), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n726), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n752), .A2(G43gat), .A3(new_n719), .A4(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n727), .A2(new_n516), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(G43gat), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT47), .ZN(G1330gat));
  NOR4_X1   g556(.A1(new_n725), .A2(G50gat), .A3(new_n438), .A4(new_n726), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n752), .A2(new_n437), .A3(new_n753), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(G50gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g560(.A1(new_n741), .A2(new_n742), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n676), .A2(new_n648), .A3(new_n677), .A4(new_n698), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n589), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n521), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n770));
  NAND2_X1  g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n767), .A2(new_n770), .A3(new_n509), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n762), .A2(new_n764), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n774), .A2(new_n589), .A3(new_n509), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT116), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n772), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n773), .B1(new_n772), .B2(new_n776), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(G1333gat));
  NAND3_X1  g578(.A1(new_n767), .A2(G71gat), .A3(new_n719), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n516), .B(KEYINPUT117), .Z(new_n781));
  OAI21_X1  g580(.A(new_n530), .B1(new_n766), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT50), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n780), .A2(new_n785), .A3(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1334gat));
  NOR2_X1   g586(.A1(new_n766), .A2(new_n438), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT118), .B(G78gat), .Z(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1335gat));
  AND2_X1   g589(.A1(new_n676), .A2(new_n677), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n647), .ZN(new_n792));
  AND4_X1   g591(.A1(KEYINPUT51), .A2(new_n524), .A3(new_n699), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT51), .B1(new_n733), .B2(new_n792), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n795), .A2(new_n589), .ZN(new_n796));
  AOI21_X1  g595(.A(G85gat), .B1(new_n796), .B2(new_n521), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n792), .A2(new_n589), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n736), .B2(new_n743), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n521), .A2(G85gat), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n797), .B1(new_n799), .B2(new_n801), .ZN(G1336gat));
  NOR2_X1   g601(.A1(new_n460), .A2(G92gat), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n795), .A2(new_n589), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n799), .A2(new_n509), .ZN(new_n807));
  INV_X1    g606(.A(G92gat), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n805), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n799), .B2(new_n509), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT52), .B1(new_n810), .B2(new_n804), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1337gat));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n543), .A3(new_n516), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n799), .A2(new_n719), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n543), .B2(new_n814), .ZN(G1338gat));
  AOI21_X1  g614(.A(new_n544), .B1(new_n799), .B2(new_n437), .ZN(new_n816));
  INV_X1    g615(.A(new_n589), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(G106gat), .A3(new_n438), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT119), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n795), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT53), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n798), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n752), .A2(new_n437), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G106gat), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n818), .B1(new_n793), .B2(new_n794), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT120), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830));
  AOI211_X1 g629(.A(new_n830), .B(new_n827), .C1(new_n823), .C2(G106gat), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n821), .B1(new_n829), .B2(new_n831), .ZN(G1339gat));
  OR2_X1    g631(.A1(new_n737), .A2(new_n738), .ZN(new_n833));
  INV_X1    g632(.A(new_n639), .ZN(new_n834));
  OR3_X1    g633(.A1(new_n632), .A2(new_n633), .A3(new_n631), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n620), .B1(new_n628), .B2(new_n619), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n645), .B2(new_n646), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n583), .B2(new_n588), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n555), .A2(new_n557), .A3(new_n562), .A4(new_n567), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n565), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n563), .A2(new_n844), .A3(new_n564), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n575), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n841), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n565), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n848), .A2(KEYINPUT55), .A3(new_n575), .A4(new_n845), .ZN(new_n849));
  AND4_X1   g648(.A1(new_n578), .A2(new_n647), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n833), .B1(new_n840), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n839), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n847), .A2(new_n578), .A3(new_n849), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n739), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n791), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n764), .A2(new_n589), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n509), .A2(new_n459), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n520), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n647), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n589), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g663(.A1(new_n859), .A2(new_n678), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(new_n331), .ZN(G1342gat));
  NOR2_X1   g665(.A1(new_n859), .A2(new_n698), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n333), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n869), .B(new_n870), .C1(new_n333), .C2(new_n867), .ZN(G1343gat));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n850), .B1(new_n589), .B2(new_n852), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n854), .B1(new_n873), .B2(new_n699), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n856), .B1(new_n874), .B2(new_n678), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT57), .B1(new_n875), .B2(new_n438), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n877), .B(new_n437), .C1(new_n855), .C2(new_n856), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n718), .A2(new_n858), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n876), .A2(new_n647), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n872), .B1(new_n881), .B2(G141gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n437), .B1(new_n855), .B2(new_n856), .ZN(new_n883));
  NOR4_X1   g682(.A1(new_n883), .A2(G141gat), .A3(new_n648), .A4(new_n879), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n881), .B2(G141gat), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n882), .A2(new_n885), .A3(KEYINPUT58), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  AOI221_X4 g686(.A(new_n884), .B1(new_n872), .B2(new_n887), .C1(new_n881), .C2(G141gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n886), .A2(new_n888), .ZN(G1344gat));
  INV_X1    g688(.A(new_n883), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n890), .A2(new_n308), .A3(new_n589), .A4(new_n880), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n878), .A3(new_n880), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT59), .B(new_n308), .C1(new_n893), .C2(new_n589), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n873), .A2(new_n699), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n853), .A2(new_n699), .A3(new_n852), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n678), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n589), .B2(new_n764), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n438), .A2(KEYINPUT57), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n899), .A2(new_n900), .B1(new_n883), .B2(KEYINPUT57), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n589), .A3(new_n880), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n895), .B1(new_n902), .B2(G148gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n891), .B1(new_n894), .B2(new_n903), .ZN(G1345gat));
  NAND2_X1  g703(.A1(new_n791), .A2(G155gat), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT122), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n791), .A3(new_n880), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n893), .A2(new_n906), .B1(new_n907), .B2(new_n304), .ZN(G1346gat));
  OAI21_X1  g707(.A(G162gat), .B1(new_n892), .B2(new_n833), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n890), .A2(new_n305), .A3(new_n699), .A4(new_n880), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n855), .A2(new_n856), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(new_n521), .A3(new_n460), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n520), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n647), .B1(new_n276), .B2(new_n277), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n460), .A2(new_n521), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n438), .B(new_n916), .C1(new_n855), .C2(new_n856), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n917), .A2(new_n648), .A3(new_n781), .ZN(new_n918));
  OAI22_X1  g717(.A1(new_n914), .A2(new_n915), .B1(new_n918), .B2(new_n231), .ZN(G1348gat));
  INV_X1    g718(.A(new_n914), .ZN(new_n920));
  AOI21_X1  g719(.A(G176gat), .B1(new_n920), .B2(new_n589), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n917), .A2(new_n781), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(G176gat), .A3(new_n589), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(KEYINPUT123), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(KEYINPUT123), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(G1349gat));
  OR2_X1    g725(.A1(new_n222), .A2(new_n223), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n913), .A2(new_n791), .A3(new_n927), .A4(new_n520), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n917), .A2(new_n678), .A3(new_n781), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n257), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n931), .A2(KEYINPUT60), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(KEYINPUT60), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n929), .A2(new_n257), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n935), .A2(new_n931), .A3(KEYINPUT60), .A4(new_n928), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n934), .A2(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n221), .A3(new_n739), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n699), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(G190gat), .ZN(new_n941));
  AOI211_X1 g740(.A(KEYINPUT61), .B(new_n221), .C1(new_n922), .C2(new_n699), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1351gat));
  NAND2_X1  g742(.A1(new_n899), .A2(new_n900), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n883), .A2(KEYINPUT57), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n944), .A2(new_n945), .A3(new_n718), .A4(new_n916), .ZN(new_n946));
  OAI21_X1  g745(.A(G197gat), .B1(new_n946), .B2(new_n648), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n912), .A2(new_n521), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n718), .A2(new_n437), .A3(new_n509), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT125), .Z(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n648), .A2(G197gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(G1352gat));
  AND3_X1   g752(.A1(new_n944), .A2(new_n945), .A3(new_n916), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n954), .A2(KEYINPUT126), .A3(new_n589), .A4(new_n718), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n956), .B1(new_n946), .B2(new_n817), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n955), .A2(G204gat), .A3(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(G204gat), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n948), .A2(new_n959), .A3(new_n589), .A4(new_n950), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT62), .Z(new_n961));
  NAND2_X1  g760(.A1(new_n958), .A2(new_n961), .ZN(G1353gat));
  OR3_X1    g761(.A1(new_n951), .A2(G211gat), .A3(new_n678), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n901), .A2(new_n791), .A3(new_n718), .A4(new_n916), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  INV_X1    g767(.A(new_n946), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n699), .A2(G218gat), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT127), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n948), .A2(new_n739), .A3(new_n950), .ZN(new_n972));
  INV_X1    g771(.A(G218gat), .ZN(new_n973));
  AOI22_X1  g772(.A1(new_n969), .A2(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G1355gat));
endmodule


