//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n462), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT65), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n471), .B(G125), .C1(new_n463), .C2(new_n464), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n468), .B1(new_n474), .B2(G2105), .ZN(G160));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n462), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n463), .A2(new_n464), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n482), .B1(G136), .B2(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n463), .B2(new_n464), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n476), .A2(new_n477), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(new_n496), .A3(new_n492), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n490), .B1(new_n494), .B2(new_n497), .ZN(G164));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI21_X1  g085(.A(G543), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n504), .A2(new_n513), .ZN(G166));
  NAND3_X1  g089(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n515));
  AND3_X1   g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT7), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT66), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n515), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G89), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n509), .A2(new_n525), .B1(new_n511), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G168));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n509), .A2(new_n529), .B1(new_n511), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(G64), .B1(new_n506), .B2(new_n505), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n503), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  AOI22_X1  g110(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n503), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  INV_X1    g113(.A(G43), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n509), .A2(new_n538), .B1(new_n511), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT67), .Z(G188));
  OR2_X1    g122(.A1(KEYINPUT6), .A2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(KEYINPUT6), .A2(G651), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n499), .A2(new_n500), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G91), .ZN(new_n551));
  INV_X1    g126(.A(G65), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n499), .B2(new_n500), .ZN(new_n553));
  INV_X1    g128(.A(G78), .ZN(new_n554));
  INV_X1    g129(.A(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n555), .B1(new_n548), .B2(new_n549), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G53), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n558), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  NOR3_X1   g138(.A1(new_n511), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n551), .B(new_n557), .C1(new_n563), .C2(new_n564), .ZN(G299));
  NAND2_X1  g140(.A1(new_n559), .A2(G52), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n548), .A2(new_n549), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n501), .A2(new_n567), .A3(G90), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n532), .A2(new_n533), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n566), .B(new_n568), .C1(new_n569), .C2(new_n503), .ZN(G301));
  NAND3_X1  g145(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n517), .A2(KEYINPUT66), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(new_n521), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n559), .A2(G51), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n501), .A2(new_n567), .A3(G89), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n575), .A2(new_n515), .A3(new_n576), .A4(new_n577), .ZN(G286));
  INV_X1    g153(.A(G166), .ZN(G303));
  INV_X1    g154(.A(KEYINPUT69), .ZN(new_n580));
  NOR3_X1   g155(.A1(new_n506), .A2(new_n505), .A3(G74), .ZN(new_n581));
  INV_X1    g156(.A(G49), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n581), .A2(new_n503), .B1(new_n511), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n509), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n580), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n550), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n559), .A2(G49), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n587), .A2(KEYINPUT69), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n586), .A2(new_n590), .ZN(G288));
  OAI21_X1  g166(.A(G61), .B1(new_n506), .B2(new_n505), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n550), .A2(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n559), .A2(G48), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n559), .A2(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI221_X1 g176(.A(new_n599), .B1(new_n600), .B2(new_n509), .C1(new_n601), .C2(new_n503), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  AND2_X1   g178(.A1(KEYINPUT70), .A2(KEYINPUT10), .ZN(new_n604));
  NOR2_X1   g179(.A1(KEYINPUT70), .A2(KEYINPUT10), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n509), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n499), .B2(new_n500), .ZN(new_n611));
  AND2_X1   g186(.A1(G79), .A2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n559), .A2(G54), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n501), .A2(new_n567), .A3(new_n606), .A4(G92), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n609), .A2(new_n613), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n603), .B1(new_n617), .B2(G868), .ZN(G321));
  XOR2_X1   g193(.A(G321), .B(KEYINPUT71), .Z(G284));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n617), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(KEYINPUT72), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(KEYINPUT72), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n628), .B(new_n629), .C1(G868), .C2(new_n541), .ZN(G323));
  XOR2_X1   g205(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n631));
  XNOR2_X1  g206(.A(G323), .B(new_n631), .ZN(G282));
  NAND2_X1  g207(.A1(new_n495), .A2(new_n466), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n478), .A2(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n462), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  INV_X1    g216(.A(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n495), .A2(new_n462), .ZN(new_n643));
  OAI221_X1 g218(.A(new_n639), .B1(new_n640), .B2(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n637), .A2(new_n638), .A3(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n656), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n648), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n647), .A3(new_n661), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n664), .A2(new_n666), .A3(G14), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2072), .B(G2078), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT77), .B(KEYINPUT18), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n671), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT17), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n675), .B1(new_n676), .B2(new_n670), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(new_n676), .B2(new_n670), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n670), .A2(KEYINPUT78), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n670), .A2(KEYINPUT78), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n679), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n669), .A2(new_n671), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n674), .B1(new_n678), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2096), .B(G2100), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(KEYINPUT80), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT79), .B(KEYINPUT19), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n689), .A2(KEYINPUT80), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n687), .A2(new_n688), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n689), .A2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(new_n698), .B(new_n697), .S(new_n693), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT81), .ZN(new_n701));
  XOR2_X1   g276(.A(G1981), .B(G1986), .Z(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n701), .B(new_n706), .ZN(G229));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G166), .B2(new_n708), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G1971), .Z(new_n711));
  NOR2_X1   g286(.A1(G6), .A2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G305), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(G16), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n717));
  MUX2_X1   g292(.A(G23), .B(new_n717), .S(G16), .Z(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT33), .B(G1976), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n711), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G25), .ZN(new_n725));
  OR2_X1    g300(.A1(G95), .A2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT82), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n484), .A2(G131), .B1(G119), .B2(new_n478), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n724), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT35), .B(G1991), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT83), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n732), .B(new_n734), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n708), .A2(G24), .ZN(new_n736));
  INV_X1    g311(.A(G290), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n708), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1986), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n722), .A2(new_n723), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(KEYINPUT36), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT36), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n722), .A2(new_n743), .A3(new_n723), .A4(new_n740), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n724), .A2(G26), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT87), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n478), .A2(G128), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n462), .A2(G116), .ZN(new_n750));
  OAI21_X1  g325(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n751));
  INV_X1    g326(.A(G140), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n749), .B1(new_n750), .B2(new_n751), .C1(new_n752), .C2(new_n643), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT86), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n748), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT88), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G2067), .ZN(new_n758));
  NOR2_X1   g333(.A1(G29), .A2(G35), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G162), .B2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G2090), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n724), .A2(G33), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT25), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G139), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n643), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n495), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(new_n462), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT89), .ZN(new_n773));
  OR3_X1    g348(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n770), .B2(new_n772), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n765), .B1(new_n777), .B2(new_n724), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n778), .A2(G2072), .B1(new_n762), .B2(new_n763), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n758), .A2(new_n764), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G171), .A2(new_n708), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G5), .B2(new_n708), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  NAND2_X1  g360(.A1(G164), .A2(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G27), .B2(G29), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n784), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n785), .B2(new_n787), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n778), .A2(G2072), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT31), .B(G11), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT93), .ZN(new_n792));
  INV_X1    g367(.A(G28), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT30), .ZN(new_n794));
  AOI21_X1  g369(.A(G29), .B1(new_n793), .B2(KEYINPUT30), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n796), .B1(new_n724), .B2(new_n644), .C1(new_n782), .C2(new_n783), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n724), .A2(G32), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT26), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n478), .A2(G129), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n466), .A2(G105), .ZN(new_n803));
  INV_X1    g378(.A(G141), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n643), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n798), .B1(new_n806), .B2(new_n724), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT27), .B(G1996), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n797), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n708), .A2(G4), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n617), .B2(new_n708), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT84), .B(G1348), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n789), .A2(new_n790), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n708), .A2(G21), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G168), .B2(new_n708), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT92), .B(G1966), .Z(new_n818));
  XOR2_X1   g393(.A(new_n817), .B(new_n818), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n708), .A2(G20), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT95), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT23), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n621), .B2(new_n708), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT96), .B(G1956), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n819), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(KEYINPUT24), .A2(G34), .ZN(new_n826));
  NOR2_X1   g401(.A1(KEYINPUT24), .A2(G34), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n724), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT90), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G160), .B2(G29), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT91), .B(G2084), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(G16), .A2(G19), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n541), .B2(G16), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT85), .B(G1341), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n823), .A2(new_n824), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n825), .A2(new_n832), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n757), .A2(G2067), .ZN(new_n839));
  NOR4_X1   g414(.A1(new_n780), .A2(new_n815), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n745), .A2(new_n840), .ZN(G311));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n745), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n745), .B2(new_n840), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(G150));
  AND2_X1   g420(.A1(G80), .A2(G543), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n501), .B2(G67), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(new_n503), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  INV_X1    g424(.A(G55), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n509), .A2(new_n849), .B1(new_n511), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n624), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n536), .A2(new_n503), .ZN(new_n860));
  INV_X1    g435(.A(new_n540), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n860), .A2(new_n848), .A3(new_n861), .A4(new_n852), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n847), .A2(new_n503), .ZN(new_n863));
  OAI22_X1  g438(.A1(new_n537), .A2(new_n540), .B1(new_n863), .B2(new_n851), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n859), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  INV_X1    g443(.A(G860), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n867), .B2(KEYINPUT39), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n856), .B1(new_n868), .B2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(KEYINPUT100), .B(G37), .ZN(new_n872));
  INV_X1    g447(.A(new_n806), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n776), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n776), .A2(new_n873), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n730), .B(new_n634), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n777), .A2(new_n806), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(new_n874), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n494), .A2(new_n497), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n486), .A2(new_n489), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n755), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n753), .B(KEYINPUT86), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(G164), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n484), .A2(G142), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n478), .A2(G130), .ZN(new_n889));
  OR2_X1    g464(.A1(G106), .A2(G2105), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n890), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n885), .A2(new_n887), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n885), .B2(new_n887), .ZN(new_n895));
  OAI22_X1  g470(.A1(new_n878), .A2(new_n881), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n880), .A2(new_n874), .A3(new_n879), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n893), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(G160), .B(new_n644), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G162), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(new_n896), .B2(new_n900), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n872), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g483(.A(G868), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n853), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(G166), .A2(new_n717), .ZN(new_n911));
  INV_X1    g486(.A(new_n583), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n912), .B(new_n587), .C1(new_n504), .C2(new_n513), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n713), .A2(G290), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n713), .A2(G290), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n737), .A2(G305), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n919), .A2(new_n911), .A3(new_n915), .A4(new_n913), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n918), .A2(KEYINPUT42), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT42), .B1(new_n918), .B2(new_n920), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n865), .B(new_n626), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n609), .A2(new_n615), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n613), .A2(new_n614), .ZN(new_n927));
  NAND3_X1  g502(.A1(G299), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n559), .A2(new_n558), .A3(new_n562), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT9), .B1(new_n511), .B2(new_n561), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n506), .A2(new_n505), .ZN(new_n932));
  OAI22_X1  g507(.A1(new_n932), .A2(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n933), .A2(G651), .B1(new_n550), .B2(G91), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n616), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT41), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT101), .B1(new_n621), .B2(new_n616), .ZN(new_n939));
  XOR2_X1   g514(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(G299), .B(new_n616), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n939), .B(new_n941), .C1(new_n942), .C2(KEYINPUT101), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n925), .A2(new_n938), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n936), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n947), .B2(new_n939), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT101), .B1(new_n928), .B2(new_n935), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n617), .B2(G299), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n949), .A2(KEYINPUT102), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n944), .B1(new_n925), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n922), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n918), .A2(KEYINPUT42), .A3(new_n920), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT104), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n923), .B1(new_n921), .B2(new_n922), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n958), .B(new_n944), .C1(new_n952), .C2(new_n925), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n924), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n910), .B1(new_n960), .B2(new_n909), .ZN(G331));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n962));
  XNOR2_X1  g537(.A(G331), .B(new_n962), .ZN(G295));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(G168), .B2(G301), .ZN(new_n966));
  NAND3_X1  g541(.A1(G171), .A2(G286), .A3(KEYINPUT107), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n969));
  NAND3_X1  g544(.A1(G168), .A2(new_n969), .A3(G301), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT106), .B1(G171), .B2(G286), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n862), .A2(new_n864), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n968), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n968), .B2(new_n972), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n943), .B(new_n938), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n968), .A2(new_n972), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n865), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n949), .A2(new_n950), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n968), .A2(new_n972), .A3(new_n973), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n976), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n918), .A2(new_n920), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n978), .A2(new_n980), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n940), .B1(new_n949), .B2(new_n950), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n928), .A2(KEYINPUT41), .A3(new_n935), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT109), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n980), .B(new_n978), .C1(new_n948), .C2(new_n951), .ZN(new_n990));
  INV_X1    g565(.A(new_n983), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n984), .A2(new_n992), .A3(new_n872), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT110), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n984), .A2(new_n992), .A3(new_n995), .A4(new_n872), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n964), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n976), .A2(new_n991), .A3(new_n981), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n999));
  INV_X1    g574(.A(G37), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1001), .A2(new_n984), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n999), .B1(new_n998), .B2(new_n1000), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT43), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT44), .B1(new_n997), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1001), .A2(new_n984), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT43), .B1(new_n1007), .B2(new_n1003), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n984), .A2(new_n992), .A3(new_n964), .A4(new_n872), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1006), .A2(new_n1012), .ZN(G397));
  NAND3_X1  g588(.A1(new_n465), .A2(new_n467), .A3(G40), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT111), .B(G1384), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(G164), .B2(new_n1017), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n1014), .B(new_n1018), .C1(G2105), .C2(new_n474), .ZN(new_n1019));
  INV_X1    g594(.A(G2067), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n755), .B(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n806), .B(G1996), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n731), .A2(new_n734), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n731), .A2(new_n734), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(G290), .B(G1986), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1019), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1015), .B1(G164), .B2(G1384), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n884), .A2(KEYINPUT45), .A3(new_n1016), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1014), .B1(new_n474), .B2(G2105), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n785), .A4(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n1035));
  INV_X1    g610(.A(G1384), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n884), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1037), .A3(new_n1030), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n783), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n884), .A2(KEYINPUT45), .A3(new_n1036), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n785), .A2(KEYINPUT53), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1028), .A2(new_n1040), .A3(new_n1030), .A4(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1033), .A2(new_n1039), .A3(G301), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT124), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1031), .A2(new_n1032), .B1(new_n1038), .B2(new_n783), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT124), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1046), .A2(new_n1047), .A3(G301), .A4(new_n1043), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n468), .A2(KEYINPUT123), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n468), .A2(KEYINPUT123), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1042), .A2(G40), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n474), .A2(G2105), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1018), .A2(new_n1054), .A3(new_n1029), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1046), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1050), .B1(new_n1057), .B2(G171), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1049), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT125), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1049), .A2(new_n1058), .A3(KEYINPUT125), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n1064));
  INV_X1    g639(.A(G1956), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1038), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(G299), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n1070));
  OR2_X1    g645(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1071));
  NAND2_X1  g646(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n934), .A2(new_n931), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1064), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1038), .A2(new_n813), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1384), .B1(new_n882), .B2(new_n883), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1030), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1020), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n616), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1075), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1076), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1066), .A2(new_n1075), .A3(new_n1068), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1087), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n1084), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1030), .B1(new_n1078), .B2(KEYINPUT45), .ZN(new_n1092));
  NOR3_X1   g667(.A1(G164), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1092), .A2(new_n1093), .A3(G1996), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1095));
  XOR2_X1   g670(.A(new_n1095), .B(G1341), .Z(new_n1096));
  NOR2_X1   g671(.A1(new_n1080), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n541), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT59), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1077), .A2(new_n1081), .A3(new_n616), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT60), .B1(new_n1102), .B2(new_n1082), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1038), .A2(new_n813), .B1(new_n1080), .B2(new_n1020), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1098), .A2(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1091), .A2(new_n1101), .A3(new_n1103), .A4(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1087), .A2(KEYINPUT61), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1076), .A2(new_n1109), .A3(new_n1085), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1088), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(G301), .B1(new_n1046), .B2(new_n1043), .ZN(new_n1112));
  AND4_X1   g687(.A1(G301), .A2(new_n1033), .A3(new_n1056), .A4(new_n1039), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1050), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G8), .ZN(new_n1115));
  NOR2_X1   g690(.A1(G168), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT51), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1034), .A2(new_n1037), .A3(new_n1030), .ZN(new_n1121));
  INV_X1    g696(.A(G2084), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1028), .A2(new_n1030), .A3(new_n1040), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1121), .A2(new_n1122), .B1(new_n1123), .B2(new_n818), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1117), .B(new_n1120), .C1(new_n1124), .C2(new_n1115), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n818), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1034), .A2(new_n1037), .A3(new_n1122), .A4(new_n1030), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(G8), .B(new_n1119), .C1(new_n1128), .C2(G286), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1116), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT112), .B(G1971), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1034), .A2(new_n1037), .A3(new_n763), .A4(new_n1030), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT55), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(G166), .B2(new_n1115), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1135), .A2(G8), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT113), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1115), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(KEYINPUT113), .A3(new_n1139), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n912), .A2(G1976), .A3(new_n587), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1079), .A2(G8), .A3(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT114), .B(G1976), .Z(new_n1148));
  NAND3_X1  g723(.A1(new_n586), .A2(new_n590), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT52), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1115), .B1(new_n1030), .B2(new_n1078), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1150), .B1(new_n1153), .B2(new_n1146), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(G86), .ZN(new_n1156));
  INV_X1    g731(.A(G48), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n509), .A2(new_n1156), .B1(new_n511), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n503), .B1(new_n592), .B2(new_n593), .ZN(new_n1159));
  OAI21_X1  g734(.A(G1981), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(G1981), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n595), .A2(new_n596), .A3(new_n1161), .A4(new_n597), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT115), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1160), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT49), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT49), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1164), .A2(new_n1168), .A3(new_n1165), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1167), .A2(new_n1153), .A3(new_n1169), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1155), .B(new_n1170), .C1(new_n1139), .C2(new_n1143), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  AND4_X1   g747(.A1(new_n1114), .A2(new_n1131), .A3(new_n1145), .A4(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1063), .A2(new_n1111), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1131), .A2(KEYINPUT62), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1171), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1125), .A2(new_n1129), .A3(new_n1177), .A4(new_n1130), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1175), .A2(new_n1176), .A3(new_n1112), .A4(new_n1178), .ZN(new_n1179));
  AND4_X1   g754(.A1(new_n1142), .A2(new_n1144), .A3(new_n1170), .A4(new_n1155), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1181));
  NOR2_X1   g756(.A1(G288), .A2(G1976), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1115), .B(new_n1080), .C1(new_n1183), .C2(new_n1162), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1124), .A2(new_n1115), .A3(G286), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n1176), .B2(new_n1186), .ZN(new_n1187));
  AND4_X1   g762(.A1(KEYINPUT63), .A2(new_n1172), .A3(new_n1145), .A4(new_n1186), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1179), .B(new_n1185), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1027), .B1(new_n1174), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(G1996), .ZN(new_n1191));
  AOI21_X1  g766(.A(KEYINPUT46), .B1(new_n1019), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1021), .A2(new_n806), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1192), .B1(new_n1193), .B2(new_n1019), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1019), .A2(KEYINPUT46), .A3(new_n1191), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1195), .A2(KEYINPUT126), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1195), .A2(KEYINPUT126), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1198), .B(KEYINPUT47), .Z(new_n1199));
  NAND2_X1  g774(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1200));
  OAI22_X1  g775(.A1(new_n1200), .A2(new_n1023), .B1(G2067), .B2(new_n755), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1019), .ZN(new_n1202));
  INV_X1    g777(.A(G1986), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1019), .A2(new_n1203), .A3(new_n737), .ZN(new_n1204));
  XOR2_X1   g779(.A(new_n1204), .B(KEYINPUT48), .Z(new_n1205));
  AND2_X1   g780(.A1(new_n1025), .A2(new_n1019), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1202), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1199), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1190), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g784(.A1(new_n460), .A2(G227), .ZN(new_n1211));
  NAND3_X1  g785(.A1(new_n667), .A2(KEYINPUT127), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g786(.A(KEYINPUT127), .B1(new_n667), .B2(new_n1211), .ZN(new_n1213));
  NOR2_X1   g787(.A1(new_n1213), .A2(G229), .ZN(new_n1214));
  NAND4_X1  g788(.A1(new_n1010), .A2(new_n907), .A3(new_n1212), .A4(new_n1214), .ZN(G225));
  INV_X1    g789(.A(G225), .ZN(G308));
endmodule


