//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n450, new_n453, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n591, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1125, new_n1126, new_n1127;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n456), .A2(new_n460), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(G101), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n468), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n475), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n483), .A2(new_n468), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n473), .A2(G126), .A3(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n480), .A2(new_n482), .A3(G138), .A4(new_n468), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n473), .A2(KEYINPUT4), .A3(G138), .A4(new_n468), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n498));
  AND4_X1   g073(.A1(new_n492), .A2(new_n495), .A3(new_n496), .A4(new_n498), .ZN(G164));
  XOR2_X1   g074(.A(KEYINPUT5), .B(G543), .Z(new_n500));
  INV_X1    g075(.A(G62), .ZN(new_n501));
  OR3_X1    g076(.A1(new_n500), .A2(KEYINPUT70), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT70), .B1(new_n500), .B2(new_n501), .ZN(new_n503));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n504), .B(KEYINPUT71), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G651), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n511), .A2(G543), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n514), .A2(G88), .B1(new_n515), .B2(G50), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n511), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n511), .A2(G89), .ZN(new_n523));
  NAND2_X1  g098(.A1(G63), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n500), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n522), .A2(new_n525), .ZN(G168));
  INV_X1    g101(.A(G52), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n527), .A2(new_n520), .B1(new_n513), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OR3_X1    g108(.A1(new_n529), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n530), .B1(new_n529), .B2(new_n533), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(new_n514), .A2(G81), .B1(new_n515), .B2(G43), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  XOR2_X1   g114(.A(new_n539), .B(KEYINPUT73), .Z(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  XNOR2_X1  g122(.A(new_n500), .B(KEYINPUT74), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT75), .B(G65), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(G78), .A2(G543), .ZN(new_n551));
  OAI21_X1  g126(.A(G651), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n520), .A2(KEYINPUT9), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT9), .B1(new_n520), .B2(new_n555), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n556), .A2(new_n557), .B1(G91), .B2(new_n514), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND2_X1  g137(.A1(new_n514), .A2(G87), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n515), .A2(G49), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  AOI22_X1  g141(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n532), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(KEYINPUT77), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n514), .A2(G86), .B1(new_n515), .B2(G48), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(KEYINPUT77), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G305));
  AOI22_X1  g147(.A1(new_n514), .A2(G85), .B1(new_n515), .B2(G47), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(new_n532), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n575), .A2(KEYINPUT78), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(KEYINPUT78), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(G290));
  NAND2_X1  g153(.A1(new_n514), .A2(G92), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT10), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(G54), .B2(new_n515), .ZN(new_n581));
  INV_X1    g156(.A(G66), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n548), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g158(.A1(G79), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(G868), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(G868), .B2(G171), .ZN(G284));
  XOR2_X1   g163(.A(G284), .B(KEYINPUT79), .Z(G321));
  NAND2_X1  g164(.A1(G286), .A2(G868), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n554), .A2(new_n558), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(G868), .ZN(G297));
  OAI21_X1  g167(.A(new_n590), .B1(new_n591), .B2(G868), .ZN(G280));
  INV_X1    g168(.A(new_n586), .ZN(new_n594));
  INV_X1    g169(.A(G559), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(G860), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT80), .ZN(G148));
  NAND2_X1  g172(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n541), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n484), .A2(G2104), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT12), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT13), .ZN(new_n605));
  INV_X1    g180(.A(G2100), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n484), .A2(G135), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n486), .A2(G123), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n468), .A2(G111), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(G2096), .Z(new_n614));
  NAND3_X1  g189(.A1(new_n607), .A2(new_n608), .A3(new_n614), .ZN(G156));
  XNOR2_X1  g190(.A(KEYINPUT15), .B(G2435), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT83), .B(G2438), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(G2427), .B(G2430), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(KEYINPUT14), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(G1341), .B(G1348), .Z(new_n623));
  XNOR2_X1  g198(.A(G2443), .B(G2446), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n622), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2451), .B(G2454), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(G14), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(new_n626), .ZN(G401));
  XOR2_X1   g206(.A(G2067), .B(G2678), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT84), .ZN(new_n633));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n635), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT17), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT18), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g216(.A1(G2072), .A2(G2078), .ZN(new_n642));
  OAI22_X1  g217(.A1(new_n636), .A2(new_n640), .B1(new_n444), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2096), .B(G2100), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(G227));
  XOR2_X1   g221(.A(G1971), .B(G1976), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT19), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1956), .B(G2474), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1961), .B(G1966), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NOR3_X1   g227(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n648), .A2(new_n651), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT20), .Z(new_n655));
  AOI211_X1 g230(.A(new_n653), .B(new_n655), .C1(new_n648), .C2(new_n652), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1991), .B(G1996), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1981), .B(G1986), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G229));
  INV_X1    g237(.A(G29), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G27), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT93), .Z(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(G164), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2078), .ZN(new_n667));
  INV_X1    g242(.A(G34), .ZN(new_n668));
  AOI21_X1  g243(.A(G29), .B1(new_n668), .B2(KEYINPUT24), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(KEYINPUT24), .B2(new_n668), .ZN(new_n670));
  INV_X1    g245(.A(G125), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n477), .B1(new_n483), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G2105), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n484), .A2(G137), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(new_n674), .A3(new_n471), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n670), .B1(new_n675), .B2(new_n663), .ZN(new_n676));
  INV_X1    g251(.A(G2084), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NOR2_X1   g254(.A1(G168), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n679), .B2(G21), .ZN(new_n681));
  INV_X1    g256(.A(G1966), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT25), .Z(new_n685));
  INV_X1    g260(.A(G139), .ZN(new_n686));
  AOI22_X1  g261(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n687));
  OAI221_X1 g262(.A(new_n685), .B1(new_n474), .B2(new_n686), .C1(new_n687), .C2(new_n468), .ZN(new_n688));
  MUX2_X1   g263(.A(G33), .B(new_n688), .S(G29), .Z(new_n689));
  AOI211_X1 g264(.A(new_n667), .B(new_n683), .C1(G2072), .C2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G1961), .ZN(new_n691));
  NOR2_X1   g266(.A1(G5), .A2(G16), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT92), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G301), .B2(new_n679), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT27), .B(G1996), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n663), .A2(G32), .ZN(new_n698));
  NAND3_X1  g273(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT26), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G129), .B2(new_n486), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n698), .B1(new_n704), .B2(new_n663), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT88), .ZN(new_n706));
  OAI221_X1 g281(.A(new_n690), .B1(new_n691), .B2(new_n694), .C1(new_n697), .C2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n679), .A2(G4), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n594), .B2(new_n679), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1348), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n681), .A2(new_n682), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n689), .A2(G2072), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT31), .B(G11), .Z(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT91), .Z(new_n714));
  INV_X1    g289(.A(G28), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(KEYINPUT30), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT30), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n663), .B1(new_n717), .B2(G28), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n714), .B1(new_n716), .B2(new_n718), .C1(new_n613), .C2(new_n663), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n676), .A2(new_n677), .ZN(new_n720));
  NOR4_X1   g295(.A1(new_n711), .A2(new_n712), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n663), .A2(G26), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT28), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n486), .A2(G128), .ZN(new_n724));
  INV_X1    g299(.A(G140), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n474), .ZN(new_n726));
  OAI21_X1  g301(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n727));
  INV_X1    g302(.A(G116), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G2105), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT87), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n723), .B1(new_n731), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2067), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n663), .A2(G35), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT94), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G162), .B2(new_n663), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT29), .B(G2090), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n721), .A2(new_n733), .A3(new_n738), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n707), .A2(new_n710), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n679), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT23), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n591), .B2(new_n679), .ZN(new_n743));
  INV_X1    g318(.A(G1956), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n706), .A2(new_n697), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT90), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n679), .A2(G19), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n541), .B2(new_n679), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1341), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n691), .B2(new_n694), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n740), .A2(new_n745), .A3(new_n747), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT95), .ZN(new_n753));
  XOR2_X1   g328(.A(G288), .B(KEYINPUT86), .Z(new_n754));
  MUX2_X1   g329(.A(G23), .B(new_n754), .S(G16), .Z(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT33), .B(G1976), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n679), .A2(G22), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G166), .B2(new_n679), .ZN(new_n759));
  INV_X1    g334(.A(G1971), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  MUX2_X1   g336(.A(G6), .B(G305), .S(G16), .Z(new_n762));
  XOR2_X1   g337(.A(KEYINPUT32), .B(G1981), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n757), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(KEYINPUT34), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(KEYINPUT34), .ZN(new_n767));
  OR2_X1    g342(.A1(G95), .A2(G2105), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n768), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT85), .Z(new_n770));
  AOI22_X1  g345(.A1(G119), .A2(new_n486), .B1(new_n484), .B2(G131), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G25), .B(new_n772), .S(G29), .Z(new_n773));
  XOR2_X1   g348(.A(KEYINPUT35), .B(G1991), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(G16), .A2(G24), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G290), .B2(new_n679), .ZN(new_n777));
  INV_X1    g352(.A(G1986), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n778), .B2(new_n777), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n766), .A2(new_n767), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT36), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n753), .A2(new_n782), .ZN(G150));
  INV_X1    g358(.A(G150), .ZN(G311));
  NAND2_X1  g359(.A1(new_n514), .A2(G93), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT96), .B(G55), .Z(new_n787));
  OAI221_X1 g362(.A(new_n785), .B1(new_n532), .B2(new_n786), .C1(new_n520), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n540), .A2(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n539), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT38), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n594), .A2(G559), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(KEYINPUT39), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(KEYINPUT39), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n795), .A2(new_n796), .A3(G860), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n788), .A2(G860), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT37), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n797), .A2(new_n799), .ZN(G145));
  AND2_X1   g375(.A1(new_n492), .A2(new_n498), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n495), .A2(new_n496), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n495), .B2(new_n496), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT100), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g382(.A(KEYINPUT100), .B(new_n801), .C1(new_n803), .C2(new_n804), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n731), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(new_n704), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n809), .B(new_n731), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(new_n703), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n688), .A2(KEYINPUT101), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n816), .A2(KEYINPUT101), .A3(new_n688), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n772), .B(new_n604), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n484), .A2(G142), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n486), .A2(G130), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n468), .A2(G118), .ZN(new_n821));
  OAI21_X1  g396(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n819), .B(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n818), .B(new_n823), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n688), .A2(KEYINPUT101), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n812), .A2(new_n814), .A3(new_n825), .A4(new_n815), .ZN(new_n826));
  AND3_X1   g401(.A1(new_n817), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n824), .B1(new_n817), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n675), .B(new_n490), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n613), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n831), .B(new_n832), .Z(new_n833));
  AOI21_X1  g408(.A(G37), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT102), .ZN(new_n835));
  INV_X1    g410(.A(new_n829), .ZN(new_n836));
  INV_X1    g411(.A(new_n833), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n835), .B(new_n837), .C1(new_n827), .C2(new_n828), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n834), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT103), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(new_n834), .C1(new_n838), .C2(new_n840), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n842), .A2(KEYINPUT40), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT40), .B1(new_n842), .B2(new_n844), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(G395));
  NOR2_X1   g422(.A1(new_n788), .A2(G868), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n598), .B(KEYINPUT104), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n791), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n591), .A2(new_n586), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n594), .A2(G299), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n594), .A2(KEYINPUT105), .A3(G299), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(KEYINPUT41), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n851), .A2(new_n857), .A3(new_n853), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n850), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n754), .B(G166), .ZN(new_n860));
  XOR2_X1   g435(.A(G290), .B(G305), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT42), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n854), .A2(new_n855), .ZN(new_n864));
  OAI221_X1 g439(.A(new_n859), .B1(KEYINPUT106), .B2(new_n863), .C1(new_n850), .C2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(KEYINPUT106), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n865), .B(new_n866), .Z(new_n867));
  AOI21_X1  g442(.A(new_n848), .B1(new_n867), .B2(G868), .ZN(G295));
  AOI21_X1  g443(.A(new_n848), .B1(new_n867), .B2(G868), .ZN(G331));
  NAND2_X1  g444(.A1(new_n856), .A2(new_n858), .ZN(new_n870));
  NAND2_X1  g445(.A1(G301), .A2(KEYINPUT107), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT107), .ZN(new_n873));
  AOI21_X1  g448(.A(G286), .B1(G171), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n876), .A3(new_n871), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n791), .ZN(new_n883));
  INV_X1    g458(.A(new_n791), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n884), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n870), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n864), .A3(new_n885), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n889), .B2(new_n862), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n857), .B1(new_n883), .B2(new_n885), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n851), .A2(new_n853), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n862), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n864), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n891), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n890), .A2(KEYINPUT43), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n862), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n887), .A2(new_n897), .A3(new_n888), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT43), .B1(new_n890), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT44), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n888), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n883), .A2(new_n885), .B1(new_n856), .B2(new_n858), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n862), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n898), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT43), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n890), .A2(new_n908), .A3(new_n895), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n906), .B1(new_n905), .B2(KEYINPUT43), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n900), .B1(new_n912), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g488(.A1(new_n495), .A2(new_n496), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT99), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n495), .A2(new_n496), .A3(new_n802), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT100), .B1(new_n917), .B2(new_n801), .ZN(new_n918));
  INV_X1    g493(.A(new_n808), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G1384), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT45), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n923));
  INV_X1    g498(.A(G40), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n675), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(G160), .A2(KEYINPUT110), .A3(G40), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G2067), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n731), .B(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n703), .B(G1996), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n770), .A2(new_n774), .A3(new_n771), .ZN(new_n934));
  INV_X1    g509(.A(new_n774), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n772), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(G290), .B(G1986), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n928), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G8), .ZN(new_n940));
  AOI21_X1  g515(.A(G1384), .B1(new_n917), .B2(new_n801), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(KEYINPUT45), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n801), .A2(new_n495), .A3(new_n496), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n921), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n925), .B(new_n926), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n682), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT50), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n944), .A2(KEYINPUT50), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n949), .A2(new_n927), .A3(new_n677), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n940), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT51), .B1(new_n952), .B2(KEYINPUT124), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(G168), .A3(new_n951), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(G8), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(G8), .ZN(new_n956));
  AOI21_X1  g531(.A(G168), .B1(new_n947), .B2(new_n951), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n955), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G301), .B1(new_n959), .B2(KEYINPUT62), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n920), .A2(KEYINPUT112), .A3(KEYINPUT45), .A4(new_n921), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n807), .A2(KEYINPUT45), .A3(new_n921), .A4(new_n808), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n944), .B2(new_n945), .ZN(new_n968));
  AOI211_X1 g543(.A(KEYINPUT111), .B(KEYINPUT45), .C1(new_n943), .C2(new_n921), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n927), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n961), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  AOI211_X1 g547(.A(KEYINPUT113), .B(new_n970), .C1(new_n962), .C2(new_n965), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n443), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n949), .A2(new_n927), .A3(new_n950), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n974), .A2(new_n975), .B1(new_n691), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n978));
  OR3_X1    g553(.A1(new_n942), .A2(new_n946), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n960), .B(new_n980), .C1(KEYINPUT62), .C2(new_n959), .ZN(new_n981));
  XOR2_X1   g556(.A(G171), .B(KEYINPUT54), .Z(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NOR4_X1   g558(.A1(new_n922), .A2(new_n924), .A3(new_n675), .A4(new_n978), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n982), .B1(new_n984), .B2(new_n966), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n977), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n986), .A3(new_n959), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n970), .B1(new_n962), .B2(new_n965), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(new_n442), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n925), .A2(new_n926), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n943), .A2(new_n948), .A3(new_n921), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(KEYINPUT118), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(KEYINPUT118), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n805), .A2(new_n921), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n744), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n991), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n554), .A2(new_n1002), .A3(new_n558), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n554), .B2(new_n558), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n992), .A2(new_n997), .A3(G2067), .ZN(new_n1008));
  INV_X1    g583(.A(G1348), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n976), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(new_n586), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT122), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1006), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT61), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1001), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1005), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n594), .B1(new_n1010), .B2(KEYINPUT60), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1010), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT123), .B1(new_n1010), .B2(KEYINPUT60), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n976), .A2(new_n1009), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1008), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT60), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n586), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(KEYINPUT60), .A3(new_n1023), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT123), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1010), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1021), .A2(new_n1031), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1001), .A2(new_n1005), .A3(KEYINPUT61), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1017), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n966), .A2(new_n971), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(G1996), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT58), .B(G1341), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n927), .B2(new_n941), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n541), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT59), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1013), .B1(new_n1034), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n981), .B1(new_n987), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G166), .A2(new_n940), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT55), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n972), .A2(new_n973), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT114), .B(G2090), .ZN(new_n1047));
  INV_X1    g622(.A(new_n999), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1046), .A2(new_n760), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1045), .B1(new_n1049), .B2(new_n940), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1044), .B(KEYINPUT115), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n972), .A2(new_n973), .A3(G1971), .ZN(new_n1052));
  INV_X1    g627(.A(new_n976), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1047), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(G8), .B(new_n1051), .C1(new_n1052), .C2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(G305), .A2(G1981), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n570), .A2(KEYINPUT117), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n570), .A2(KEYINPUT117), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1058), .B(new_n1059), .C1(new_n532), .C2(new_n567), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1057), .B1(new_n1060), .B2(G1981), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n940), .B1(new_n927), .B2(new_n941), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1976), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1063), .B1(new_n1066), .B2(new_n754), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT52), .ZN(new_n1069));
  NOR2_X1   g644(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1067), .A2(new_n1069), .B1(G288), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1072));
  AND4_X1   g647(.A1(new_n1050), .A2(new_n1056), .A3(new_n1065), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1042), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(G288), .A2(G1976), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1065), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1063), .B1(new_n1076), .B2(new_n1057), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1072), .A2(new_n1065), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1077), .B1(new_n1056), .B2(new_n1078), .ZN(new_n1079));
  AND4_X1   g654(.A1(G168), .A2(new_n1072), .A3(new_n1065), .A4(new_n952), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1035), .A2(KEYINPUT113), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n988), .A2(new_n961), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n760), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1048), .A2(new_n1047), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n940), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1056), .B(new_n1080), .C1(new_n1044), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1050), .A2(KEYINPUT119), .A3(new_n1056), .A4(new_n1080), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1045), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(KEYINPUT63), .A3(new_n1056), .A4(new_n1080), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1079), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1074), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g672(.A(KEYINPUT120), .B(new_n1079), .C1(new_n1091), .C2(new_n1094), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n939), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1996), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT46), .B1(new_n928), .B2(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n928), .A2(KEYINPUT46), .A3(new_n1100), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n930), .A2(new_n704), .ZN(new_n1103));
  AOI211_X1 g678(.A(new_n1101), .B(new_n1102), .C1(new_n928), .C2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(KEYINPUT126), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1105), .A2(KEYINPUT47), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(KEYINPUT47), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n937), .A2(new_n928), .ZN(new_n1108));
  NOR2_X1   g683(.A1(G290), .A2(G1986), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n928), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT48), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1111), .B2(new_n1110), .ZN(new_n1113));
  INV_X1    g688(.A(new_n933), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n934), .B(KEYINPUT125), .ZN(new_n1115));
  OAI22_X1  g690(.A1(new_n1114), .A2(new_n1115), .B1(G2067), .B2(new_n731), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(new_n928), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1106), .A2(new_n1107), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT127), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1106), .A2(new_n1107), .A3(KEYINPUT127), .A4(new_n1117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1099), .A2(new_n1122), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g698(.A1(new_n842), .A2(new_n844), .ZN(new_n1125));
  NOR4_X1   g699(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1126));
  OAI21_X1  g700(.A(new_n1126), .B1(new_n910), .B2(new_n911), .ZN(new_n1127));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1127), .ZN(G308));
  OR2_X1    g702(.A1(new_n1125), .A2(new_n1127), .ZN(G225));
endmodule


