

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595;

  XOR2_X1 U325 ( .A(n438), .B(KEYINPUT47), .Z(n293) );
  NAND2_X1 U326 ( .A1(n442), .A2(n299), .ZN(n298) );
  NOR2_X1 U327 ( .A1(n574), .A2(n300), .ZN(n299) );
  INV_X1 U328 ( .A(KEYINPUT80), .ZN(n294) );
  INV_X1 U329 ( .A(KEYINPUT48), .ZN(n296) );
  XNOR2_X1 U330 ( .A(n301), .B(KEYINPUT55), .ZN(n459) );
  NOR2_X1 U331 ( .A1(n579), .A2(n476), .ZN(n301) );
  NAND2_X1 U332 ( .A1(n302), .A2(n510), .ZN(n579) );
  XNOR2_X1 U333 ( .A(n297), .B(n296), .ZN(n543) );
  NAND2_X1 U334 ( .A1(n298), .A2(n293), .ZN(n297) );
  NOR2_X1 U335 ( .A1(n588), .A2(n593), .ZN(n440) );
  XNOR2_X1 U336 ( .A(n557), .B(n439), .ZN(n593) );
  INV_X1 U337 ( .A(n441), .ZN(n300) );
  XNOR2_X1 U338 ( .A(n572), .B(n294), .ZN(n557) );
  XNOR2_X1 U339 ( .A(n375), .B(n295), .ZN(n572) );
  INV_X1 U340 ( .A(n452), .ZN(n295) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n366) );
  XNOR2_X1 U342 ( .A(n458), .B(n457), .ZN(n302) );
  XNOR2_X1 U343 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U344 ( .A(n449), .B(n448), .ZN(n450) );
  OR2_X1 U345 ( .A1(n485), .A2(n459), .ZN(n460) );
  XNOR2_X1 U346 ( .A(n484), .B(n483), .ZN(n517) );
  XOR2_X1 U347 ( .A(n444), .B(n443), .Z(n303) );
  XNOR2_X1 U348 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U349 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n457) );
  XNOR2_X1 U350 ( .A(n384), .B(n383), .ZN(n386) );
  XNOR2_X1 U351 ( .A(n390), .B(n361), .ZN(n365) );
  XOR2_X1 U352 ( .A(G176GAT), .B(G64GAT), .Z(n453) );
  XNOR2_X1 U353 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U354 ( .A(n451), .B(n450), .ZN(n455) );
  XNOR2_X1 U355 ( .A(n396), .B(n395), .ZN(n441) );
  INV_X1 U356 ( .A(G190GAT), .ZN(n489) );
  XNOR2_X1 U357 ( .A(n460), .B(KEYINPUT123), .ZN(n577) );
  INV_X1 U358 ( .A(G43GAT), .ZN(n486) );
  BUF_X1 U359 ( .A(n464), .Z(n534) );
  XNOR2_X1 U360 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U361 ( .A(n486), .B(KEYINPUT40), .ZN(n487) );
  XNOR2_X1 U362 ( .A(n492), .B(n491), .ZN(G1351GAT) );
  XNOR2_X1 U363 ( .A(n488), .B(n487), .ZN(G1330GAT) );
  XOR2_X1 U364 ( .A(KEYINPUT19), .B(KEYINPUT89), .Z(n305) );
  XNOR2_X1 U365 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n304) );
  XNOR2_X1 U366 ( .A(n305), .B(n304), .ZN(n447) );
  XOR2_X1 U367 ( .A(G120GAT), .B(G71GAT), .Z(n376) );
  XOR2_X1 U368 ( .A(n447), .B(n376), .Z(n307) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G134GAT), .ZN(n306) );
  XNOR2_X1 U370 ( .A(n307), .B(n306), .ZN(n312) );
  XNOR2_X1 U371 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n308) );
  XNOR2_X1 U372 ( .A(n308), .B(G127GAT), .ZN(n352) );
  XOR2_X1 U373 ( .A(n352), .B(G169GAT), .Z(n310) );
  NAND2_X1 U374 ( .A1(G227GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U375 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U376 ( .A(n312), .B(n311), .Z(n320) );
  XOR2_X1 U377 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n314) );
  XNOR2_X1 U378 ( .A(G190GAT), .B(G99GAT), .ZN(n313) );
  XNOR2_X1 U379 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U380 ( .A(G176GAT), .B(G183GAT), .Z(n316) );
  XNOR2_X1 U381 ( .A(G15GAT), .B(KEYINPUT90), .ZN(n315) );
  XNOR2_X1 U382 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U383 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n485) );
  XOR2_X1 U385 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n322) );
  XNOR2_X1 U386 ( .A(G162GAT), .B(G106GAT), .ZN(n321) );
  XNOR2_X1 U387 ( .A(n322), .B(n321), .ZN(n327) );
  XNOR2_X1 U388 ( .A(G78GAT), .B(KEYINPUT75), .ZN(n323) );
  XNOR2_X1 U389 ( .A(n323), .B(G148GAT), .ZN(n392) );
  XOR2_X1 U390 ( .A(n392), .B(G218GAT), .Z(n325) );
  XOR2_X1 U391 ( .A(G141GAT), .B(G22GAT), .Z(n409) );
  XNOR2_X1 U392 ( .A(G50GAT), .B(n409), .ZN(n324) );
  XNOR2_X1 U393 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U394 ( .A(n327), .B(n326), .ZN(n338) );
  XOR2_X1 U395 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n329) );
  NAND2_X1 U396 ( .A1(G228GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U397 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U398 ( .A(n330), .B(KEYINPUT24), .Z(n336) );
  XOR2_X1 U399 ( .A(G204GAT), .B(G211GAT), .Z(n332) );
  XNOR2_X1 U400 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n331) );
  XNOR2_X1 U401 ( .A(n332), .B(n331), .ZN(n444) );
  XOR2_X1 U402 ( .A(G155GAT), .B(KEYINPUT3), .Z(n334) );
  XNOR2_X1 U403 ( .A(KEYINPUT2), .B(KEYINPUT93), .ZN(n333) );
  XNOR2_X1 U404 ( .A(n334), .B(n333), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n444), .B(n350), .ZN(n335) );
  XNOR2_X1 U406 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U407 ( .A(n338), .B(n337), .ZN(n476) );
  XOR2_X1 U408 ( .A(KEYINPUT95), .B(KEYINPUT1), .Z(n340) );
  XNOR2_X1 U409 ( .A(KEYINPUT94), .B(G57GAT), .ZN(n339) );
  XNOR2_X1 U410 ( .A(n340), .B(n339), .ZN(n347) );
  XOR2_X1 U411 ( .A(KEYINPUT5), .B(G148GAT), .Z(n342) );
  XNOR2_X1 U412 ( .A(G141GAT), .B(G120GAT), .ZN(n341) );
  XNOR2_X1 U413 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U414 ( .A(n343), .B(G85GAT), .Z(n345) );
  XOR2_X1 U415 ( .A(G134GAT), .B(G162GAT), .Z(n360) );
  XNOR2_X1 U416 ( .A(G29GAT), .B(n360), .ZN(n344) );
  XNOR2_X1 U417 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U418 ( .A(n347), .B(n346), .ZN(n356) );
  XOR2_X1 U419 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n349) );
  NAND2_X1 U420 ( .A1(G225GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U421 ( .A(n349), .B(n348), .ZN(n351) );
  XOR2_X1 U422 ( .A(n351), .B(n350), .Z(n354) );
  XNOR2_X1 U423 ( .A(G1GAT), .B(n352), .ZN(n353) );
  XNOR2_X1 U424 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U425 ( .A(n356), .B(n355), .ZN(n510) );
  XOR2_X1 U426 ( .A(KEYINPUT76), .B(G85GAT), .Z(n358) );
  XNOR2_X1 U427 ( .A(G99GAT), .B(G106GAT), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n358), .B(n357), .ZN(n390) );
  XOR2_X1 U429 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n359) );
  XOR2_X1 U430 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n363) );
  NAND2_X1 U431 ( .A1(G232GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U432 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U433 ( .A(n365), .B(n364), .Z(n371) );
  XNOR2_X1 U434 ( .A(n366), .B(G29GAT), .ZN(n367) );
  XOR2_X1 U435 ( .A(n367), .B(KEYINPUT7), .Z(n369) );
  XNOR2_X1 U436 ( .A(G50GAT), .B(KEYINPUT69), .ZN(n368) );
  XNOR2_X1 U437 ( .A(n369), .B(n368), .ZN(n410) );
  XNOR2_X1 U438 ( .A(n410), .B(KEYINPUT78), .ZN(n370) );
  XNOR2_X1 U439 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U440 ( .A(KEYINPUT79), .B(G92GAT), .Z(n373) );
  XNOR2_X1 U441 ( .A(G190GAT), .B(G218GAT), .ZN(n372) );
  XNOR2_X1 U442 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U443 ( .A(G36GAT), .B(n374), .Z(n452) );
  XOR2_X1 U444 ( .A(G92GAT), .B(n453), .Z(n378) );
  XNOR2_X1 U445 ( .A(n376), .B(G204GAT), .ZN(n377) );
  XNOR2_X1 U446 ( .A(n378), .B(n377), .ZN(n384) );
  XOR2_X1 U447 ( .A(KEYINPUT77), .B(KEYINPUT33), .Z(n380) );
  XNOR2_X1 U448 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n379) );
  XNOR2_X1 U449 ( .A(n380), .B(n379), .ZN(n382) );
  AND2_X1 U450 ( .A1(G230GAT), .A2(G233GAT), .ZN(n381) );
  INV_X1 U451 ( .A(KEYINPUT32), .ZN(n385) );
  NAND2_X1 U452 ( .A1(n386), .A2(n385), .ZN(n389) );
  INV_X1 U453 ( .A(n386), .ZN(n387) );
  NAND2_X1 U454 ( .A1(n387), .A2(KEYINPUT32), .ZN(n388) );
  NAND2_X1 U455 ( .A1(n389), .A2(n388), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n390), .B(KEYINPUT74), .ZN(n394) );
  XNOR2_X1 U457 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n391), .B(KEYINPUT13), .ZN(n431) );
  XOR2_X1 U459 ( .A(n392), .B(n431), .Z(n393) );
  XNOR2_X1 U460 ( .A(n441), .B(KEYINPUT41), .ZN(n565) );
  XOR2_X1 U461 ( .A(KEYINPUT68), .B(G197GAT), .Z(n398) );
  XOR2_X1 U462 ( .A(G169GAT), .B(G8GAT), .Z(n443) );
  XOR2_X1 U463 ( .A(G15GAT), .B(G1GAT), .Z(n423) );
  XNOR2_X1 U464 ( .A(n443), .B(n423), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U466 ( .A(n399), .B(G113GAT), .Z(n404) );
  XOR2_X1 U467 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n401) );
  XNOR2_X1 U468 ( .A(KEYINPUT66), .B(KEYINPUT29), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n402), .B(G36GAT), .ZN(n403) );
  XNOR2_X1 U471 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U472 ( .A(KEYINPUT65), .B(KEYINPUT70), .Z(n406) );
  NAND2_X1 U473 ( .A1(G229GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U475 ( .A(n408), .B(n407), .Z(n412) );
  XNOR2_X1 U476 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n581) );
  INV_X1 U478 ( .A(n581), .ZN(n413) );
  AND2_X1 U479 ( .A1(n565), .A2(n413), .ZN(n414) );
  XNOR2_X1 U480 ( .A(n414), .B(KEYINPUT46), .ZN(n436) );
  XOR2_X1 U481 ( .A(KEYINPUT12), .B(KEYINPUT86), .Z(n416) );
  XNOR2_X1 U482 ( .A(G8GAT), .B(G64GAT), .ZN(n415) );
  XNOR2_X1 U483 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U484 ( .A(G78GAT), .B(G155GAT), .Z(n418) );
  XNOR2_X1 U485 ( .A(G22GAT), .B(G211GAT), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n420), .B(n419), .ZN(n435) );
  XOR2_X1 U488 ( .A(KEYINPUT85), .B(KEYINPUT14), .Z(n422) );
  XNOR2_X1 U489 ( .A(KEYINPUT82), .B(KEYINPUT15), .ZN(n421) );
  XNOR2_X1 U490 ( .A(n422), .B(n421), .ZN(n427) );
  XOR2_X1 U491 ( .A(G183GAT), .B(KEYINPUT81), .Z(n448) );
  XOR2_X1 U492 ( .A(n448), .B(G71GAT), .Z(n425) );
  XNOR2_X1 U493 ( .A(n423), .B(G127GAT), .ZN(n424) );
  XNOR2_X1 U494 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U495 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U496 ( .A1(G231GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U497 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U498 ( .A(n430), .B(KEYINPUT83), .Z(n433) );
  XNOR2_X1 U499 ( .A(n431), .B(KEYINPUT84), .ZN(n432) );
  XNOR2_X1 U500 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U501 ( .A(n435), .B(n434), .ZN(n576) );
  NOR2_X1 U502 ( .A1(n436), .A2(n576), .ZN(n437) );
  NAND2_X1 U503 ( .A1(n572), .A2(n437), .ZN(n438) );
  XNOR2_X1 U504 ( .A(n581), .B(KEYINPUT71), .ZN(n574) );
  INV_X1 U505 ( .A(KEYINPUT36), .ZN(n439) );
  INV_X1 U506 ( .A(n576), .ZN(n588) );
  XNOR2_X1 U507 ( .A(n440), .B(KEYINPUT45), .ZN(n442) );
  NAND2_X1 U508 ( .A1(G226GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U509 ( .A(n303), .B(n445), .ZN(n446) );
  XOR2_X1 U510 ( .A(n446), .B(KEYINPUT97), .Z(n451) );
  XNOR2_X1 U511 ( .A(n447), .B(KEYINPUT96), .ZN(n449) );
  XOR2_X1 U512 ( .A(n453), .B(n452), .Z(n454) );
  XNOR2_X1 U513 ( .A(n455), .B(n454), .ZN(n464) );
  XNOR2_X1 U514 ( .A(n534), .B(KEYINPUT121), .ZN(n456) );
  NOR2_X1 U515 ( .A1(n543), .A2(n456), .ZN(n458) );
  NAND2_X1 U516 ( .A1(n577), .A2(n565), .ZN(n463) );
  XOR2_X1 U517 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(G176GAT), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  INV_X1 U520 ( .A(KEYINPUT38), .ZN(n484) );
  NAND2_X1 U521 ( .A1(n574), .A2(n441), .ZN(n497) );
  INV_X1 U522 ( .A(n485), .ZN(n546) );
  NAND2_X1 U523 ( .A1(n464), .A2(n546), .ZN(n465) );
  XNOR2_X1 U524 ( .A(KEYINPUT99), .B(n465), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n476), .A2(n466), .ZN(n467) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(n467), .Z(n468) );
  XNOR2_X1 U527 ( .A(KEYINPUT100), .B(n468), .ZN(n472) );
  XOR2_X1 U528 ( .A(n534), .B(KEYINPUT27), .Z(n475) );
  NAND2_X1 U529 ( .A1(n476), .A2(n485), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT26), .ZN(n580) );
  NOR2_X1 U531 ( .A1(n475), .A2(n580), .ZN(n470) );
  XNOR2_X1 U532 ( .A(KEYINPUT98), .B(n470), .ZN(n471) );
  NOR2_X1 U533 ( .A1(n472), .A2(n471), .ZN(n473) );
  XNOR2_X1 U534 ( .A(KEYINPUT101), .B(n473), .ZN(n474) );
  NAND2_X1 U535 ( .A1(n474), .A2(n510), .ZN(n479) );
  OR2_X1 U536 ( .A1(n510), .A2(n475), .ZN(n544) );
  XNOR2_X1 U537 ( .A(n476), .B(KEYINPUT28), .ZN(n537) );
  NOR2_X1 U538 ( .A1(n544), .A2(n537), .ZN(n477) );
  NAND2_X1 U539 ( .A1(n485), .A2(n477), .ZN(n478) );
  NAND2_X1 U540 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n480), .B(KEYINPUT102), .ZN(n495) );
  NAND2_X1 U542 ( .A1(n495), .A2(n588), .ZN(n481) );
  NOR2_X1 U543 ( .A1(n593), .A2(n481), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n482), .B(KEYINPUT37), .ZN(n530) );
  NOR2_X1 U545 ( .A1(n497), .A2(n530), .ZN(n483) );
  NOR2_X1 U546 ( .A1(n485), .A2(n517), .ZN(n488) );
  NAND2_X1 U547 ( .A1(n577), .A2(n557), .ZN(n492) );
  XOR2_X1 U548 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n490) );
  INV_X1 U549 ( .A(n510), .ZN(n532) );
  OR2_X1 U550 ( .A1(n557), .A2(n588), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n493), .B(KEYINPUT87), .ZN(n494) );
  XNOR2_X1 U552 ( .A(KEYINPUT16), .B(n494), .ZN(n496) );
  NAND2_X1 U553 ( .A1(n496), .A2(n495), .ZN(n520) );
  NOR2_X1 U554 ( .A1(n497), .A2(n520), .ZN(n507) );
  NAND2_X1 U555 ( .A1(n532), .A2(n507), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n498), .B(KEYINPUT103), .ZN(n499) );
  XOR2_X1 U557 ( .A(n499), .B(KEYINPUT104), .Z(n501) );
  XNOR2_X1 U558 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n501), .B(n500), .ZN(G1324GAT) );
  XOR2_X1 U560 ( .A(G8GAT), .B(KEYINPUT105), .Z(n503) );
  NAND2_X1 U561 ( .A1(n507), .A2(n534), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(G1325GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT106), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U564 ( .A1(n507), .A2(n546), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U566 ( .A(G15GAT), .B(n506), .ZN(G1326GAT) );
  XOR2_X1 U567 ( .A(G22GAT), .B(KEYINPUT107), .Z(n509) );
  NAND2_X1 U568 ( .A1(n507), .A2(n537), .ZN(n508) );
  XNOR2_X1 U569 ( .A(n509), .B(n508), .ZN(G1327GAT) );
  XNOR2_X1 U570 ( .A(KEYINPUT108), .B(KEYINPUT39), .ZN(n512) );
  NOR2_X1 U571 ( .A1(n510), .A2(n517), .ZN(n511) );
  XNOR2_X1 U572 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U573 ( .A(G29GAT), .B(n513), .ZN(G1328GAT) );
  INV_X1 U574 ( .A(n534), .ZN(n514) );
  NOR2_X1 U575 ( .A1(n517), .A2(n514), .ZN(n516) );
  XNOR2_X1 U576 ( .A(G36GAT), .B(KEYINPUT109), .ZN(n515) );
  XNOR2_X1 U577 ( .A(n516), .B(n515), .ZN(G1329GAT) );
  INV_X1 U578 ( .A(n537), .ZN(n547) );
  NOR2_X1 U579 ( .A1(n547), .A2(n517), .ZN(n518) );
  XOR2_X1 U580 ( .A(G50GAT), .B(n518), .Z(G1331GAT) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n522) );
  NAND2_X1 U582 ( .A1(n565), .A2(n581), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(KEYINPUT110), .ZN(n531) );
  NOR2_X1 U584 ( .A1(n531), .A2(n520), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n527), .A2(n532), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(G1332GAT) );
  XOR2_X1 U587 ( .A(G64GAT), .B(KEYINPUT111), .Z(n524) );
  NAND2_X1 U588 ( .A1(n527), .A2(n534), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(G1333GAT) );
  NAND2_X1 U590 ( .A1(n546), .A2(n527), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(KEYINPUT112), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G71GAT), .B(n526), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(G78GAT), .B(KEYINPUT43), .Z(n529) );
  NAND2_X1 U594 ( .A1(n527), .A2(n537), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(G1335GAT) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n538), .A2(n532), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G85GAT), .B(n533), .ZN(G1336GAT) );
  NAND2_X1 U599 ( .A1(n538), .A2(n534), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n535), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U601 ( .A1(n546), .A2(n538), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(KEYINPUT114), .ZN(n542) );
  XOR2_X1 U604 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n540) );
  NAND2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1339GAT) );
  NOR2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n545), .B(KEYINPUT115), .ZN(n562) );
  NAND2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U611 ( .A1(n562), .A2(n548), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n574), .A2(n558), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n549), .B(KEYINPUT116), .ZN(n550) );
  XNOR2_X1 U614 ( .A(G113GAT), .B(n550), .ZN(G1340GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n552) );
  NAND2_X1 U616 ( .A1(n558), .A2(n565), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n554) );
  XOR2_X1 U618 ( .A(G120GAT), .B(KEYINPUT117), .Z(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1341GAT) );
  NAND2_X1 U620 ( .A1(n558), .A2(n576), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(KEYINPUT50), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G127GAT), .B(n556), .ZN(G1342GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n560) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(G134GAT), .B(n561), .Z(G1343GAT) );
  NOR2_X1 U627 ( .A1(n580), .A2(n562), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT120), .B(n563), .Z(n571) );
  NOR2_X1 U629 ( .A1(n581), .A2(n571), .ZN(n564) );
  XOR2_X1 U630 ( .A(G141GAT), .B(n564), .Z(G1344GAT) );
  INV_X1 U631 ( .A(n565), .ZN(n566) );
  NOR2_X1 U632 ( .A1(n571), .A2(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G148GAT), .B(n569), .ZN(G1345GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n588), .ZN(n570) );
  XOR2_X1 U637 ( .A(G155GAT), .B(n570), .Z(G1346GAT) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(G162GAT), .B(n573), .Z(G1347GAT) );
  NAND2_X1 U640 ( .A1(n574), .A2(n577), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G183GAT), .ZN(G1350GAT) );
  OR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n592) );
  NOR2_X1 U645 ( .A1(n581), .A2(n592), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n584), .ZN(G1352GAT) );
  NOR2_X1 U649 ( .A1(n441), .A2(n592), .ZN(n586) );
  XNOR2_X1 U650 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(G204GAT), .B(n587), .Z(G1353GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n592), .ZN(n590) );
  XNOR2_X1 U654 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U656 ( .A(G211GAT), .B(n591), .ZN(G1354GAT) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(n594), .Z(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

