//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G107), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT75), .B1(new_n187), .B2(G104), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT75), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G104), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G101), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT76), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n196), .A3(G101), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n190), .A2(G107), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n187), .A2(KEYINPUT3), .A3(G104), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT3), .B1(new_n187), .B2(G104), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n198), .B(new_n199), .C1(new_n200), .C2(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT74), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT74), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n187), .A2(G104), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n190), .B2(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n187), .A2(KEYINPUT3), .A3(G104), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n204), .B1(new_n209), .B2(new_n198), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n195), .B(new_n197), .C1(new_n203), .C2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT82), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G116), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n214), .B2(KEYINPUT5), .ZN(new_n215));
  INV_X1    g029(.A(G116), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G119), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n217), .A3(KEYINPUT5), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT5), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n219), .A2(new_n213), .A3(KEYINPUT82), .A4(G116), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n215), .A2(new_n218), .A3(G113), .A4(new_n220), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n221), .A2(KEYINPUT83), .ZN(new_n222));
  XNOR2_X1  g036(.A(G116), .B(G119), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT2), .A2(G113), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n226), .A2(new_n227), .B1(KEYINPUT2), .B2(G113), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n221), .A2(KEYINPUT83), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n211), .A2(new_n222), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n227), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT2), .A2(G113), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n223), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n221), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT84), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n193), .A2(new_n196), .A3(G101), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n196), .B1(new_n193), .B2(G101), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n202), .A2(KEYINPUT74), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n209), .A2(new_n204), .A3(new_n198), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n221), .A2(new_n233), .A3(KEYINPUT84), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n236), .A2(new_n239), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(G110), .B(G122), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT8), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n230), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G224), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT7), .B1(new_n248), .B2(G953), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  OR2_X1    g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G143), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n251), .B(new_n252), .C1(new_n254), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n253), .A2(G146), .ZN(new_n259));
  AND2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n250), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G125), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n252), .A2(new_n251), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n258), .A2(new_n259), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT64), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n262), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n253), .A2(G128), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G128), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n255), .A2(new_n268), .B1(new_n256), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(G143), .B(G146), .ZN(new_n272));
  INV_X1    g086(.A(new_n270), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n263), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n249), .B1(new_n267), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n252), .A2(new_n251), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n261), .B1(new_n279), .B2(new_n272), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT64), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n257), .A2(new_n250), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(G125), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n249), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n276), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n247), .A2(new_n286), .A3(KEYINPUT85), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT85), .B1(new_n247), .B2(new_n286), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n228), .B(new_n223), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(G101), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n203), .A2(new_n210), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT4), .B1(new_n209), .B2(new_n198), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n289), .B(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n239), .A2(new_n222), .A3(new_n229), .A4(new_n242), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n245), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n287), .A2(new_n288), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT86), .B1(new_n299), .B2(G902), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n295), .A2(new_n296), .ZN(new_n301));
  INV_X1    g115(.A(new_n245), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT6), .A3(new_n297), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT6), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(new_n305), .A3(new_n302), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n267), .A2(new_n277), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n248), .A2(G953), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n304), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n247), .A2(new_n286), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT85), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n297), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n311), .B(new_n312), .C1(new_n316), .C2(new_n287), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n300), .A2(new_n310), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G210), .B1(G237), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT87), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n300), .A2(new_n317), .A3(new_n319), .A4(new_n310), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G214), .B1(G237), .B2(G902), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n323), .A2(new_n322), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT99), .ZN(new_n328));
  INV_X1    g142(.A(G237), .ZN(new_n329));
  INV_X1    g143(.A(G953), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G214), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n253), .ZN(new_n332));
  NOR2_X1   g146(.A1(G237), .A2(G953), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(G143), .A3(G214), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT18), .ZN(new_n335));
  INV_X1    g149(.A(G131), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n332), .B(new_n334), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(G125), .A2(G140), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(G125), .A2(G140), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n255), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n263), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(G146), .A3(new_n338), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n335), .B(new_n336), .C1(new_n332), .C2(new_n334), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT88), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n332), .A2(new_n334), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(KEYINPUT18), .A3(G131), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT88), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n337), .A4(new_n345), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT92), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(G131), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT17), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n349), .A2(KEYINPUT92), .A3(KEYINPUT17), .A4(G131), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n332), .A2(new_n336), .A3(new_n334), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n357), .B(new_n358), .C1(KEYINPUT17), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT16), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n343), .B2(new_n338), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n263), .A2(KEYINPUT16), .A3(G140), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n255), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT16), .B1(new_n339), .B2(new_n340), .ZN(new_n366));
  INV_X1    g180(.A(new_n364), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G146), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT91), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT91), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n371), .A3(new_n368), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n353), .B1(new_n361), .B2(new_n373), .ZN(new_n374));
  XOR2_X1   g188(.A(G113), .B(G122), .Z(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT90), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(new_n190), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n377), .B(new_n353), .C1(new_n361), .C2(new_n373), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(KEYINPUT94), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT94), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n374), .A2(new_n382), .A3(new_n378), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n312), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G475), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT89), .B1(new_n339), .B2(new_n340), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT19), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n360), .B(new_n368), .C1(new_n387), .C2(G146), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n353), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n378), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n380), .ZN(new_n391));
  NOR2_X1   g205(.A1(G475), .A2(G902), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(KEYINPUT93), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT20), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT20), .ZN(new_n396));
  AOI211_X1 g210(.A(new_n396), .B(new_n393), .C1(new_n390), .C2(new_n380), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n385), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G478), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT15), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT13), .ZN(new_n402));
  INV_X1    g216(.A(G128), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(G143), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT95), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n268), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n253), .A2(G128), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT95), .A3(new_n402), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT96), .B1(new_n407), .B2(new_n402), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT96), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n410), .A2(new_n253), .A3(KEYINPUT13), .A4(G128), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n406), .A2(new_n408), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G134), .ZN(new_n413));
  XNOR2_X1  g227(.A(G128), .B(G143), .ZN(new_n414));
  INV_X1    g228(.A(G134), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G116), .B(G122), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(new_n187), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n414), .B(new_n415), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n187), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT14), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n216), .A2(KEYINPUT14), .A3(G122), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(G107), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n420), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT9), .B(G234), .ZN(new_n428));
  INV_X1    g242(.A(G217), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n428), .A2(new_n429), .A3(G953), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n419), .A2(new_n426), .A3(new_n430), .ZN(new_n433));
  AOI21_X1  g247(.A(G902), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT97), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT97), .ZN(new_n436));
  AOI211_X1 g250(.A(new_n436), .B(G902), .C1(new_n432), .C2(new_n433), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n401), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(G234), .A2(G237), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n439), .A2(G952), .A3(new_n330), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT21), .B(G898), .Z(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(G902), .A3(G953), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n444), .B(KEYINPUT98), .Z(new_n445));
  INV_X1    g259(.A(new_n433), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n430), .B1(new_n419), .B2(new_n426), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n312), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n401), .B1(new_n448), .B2(new_n436), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n438), .A2(new_n445), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n328), .B1(new_n399), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n401), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n436), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n434), .A2(KEYINPUT97), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n445), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n456), .A2(new_n457), .A3(new_n449), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n458), .A2(KEYINPUT99), .A3(new_n385), .A4(new_n398), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G221), .B1(new_n428), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(G110), .B(G140), .Z(new_n464));
  AND2_X1   g278(.A1(new_n330), .A2(G227), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT11), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n415), .B2(G137), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT65), .ZN(new_n470));
  INV_X1    g284(.A(G137), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(G134), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(KEYINPUT11), .A3(G134), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n415), .A2(KEYINPUT65), .A3(G137), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n469), .A2(new_n472), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n475), .A2(G131), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(G131), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n274), .A2(KEYINPUT77), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT77), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n272), .A2(new_n480), .A3(new_n273), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n271), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n239), .A2(new_n242), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT10), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n275), .A2(KEYINPUT10), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n294), .B1(new_n241), .B2(new_n240), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n281), .A2(new_n292), .A3(new_n282), .ZN(new_n488));
  OAI22_X1  g302(.A1(new_n211), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT80), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n211), .A2(new_n486), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n483), .A2(new_n484), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n487), .A2(new_n488), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT80), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n478), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n497));
  INV_X1    g311(.A(new_n478), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n467), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT81), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(KEYINPUT81), .B(new_n467), .C1(new_n496), .C2(new_n499), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n499), .A2(new_n467), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n271), .A2(new_n274), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n211), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n478), .B1(new_n506), .B2(new_n483), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n509), .B(KEYINPUT79), .C1(KEYINPUT12), .C2(new_n507), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT79), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n511), .A3(new_n508), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n504), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n502), .A2(new_n503), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G469), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n312), .ZN(new_n516));
  INV_X1    g330(.A(new_n499), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n517), .A3(new_n512), .ZN(new_n518));
  INV_X1    g332(.A(new_n496), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n518), .A2(new_n467), .B1(new_n519), .B2(new_n504), .ZN(new_n520));
  OAI21_X1  g334(.A(G469), .B1(new_n520), .B2(G902), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n463), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT73), .ZN(new_n523));
  XNOR2_X1  g337(.A(G119), .B(G128), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT24), .B(G110), .Z(new_n525));
  AOI22_X1  g339(.A1(new_n365), .A2(new_n368), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n213), .A2(G128), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT23), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(G119), .B2(new_n403), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n213), .A2(KEYINPUT23), .A3(G128), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT69), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n533), .B(new_n527), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n534), .A3(G110), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n526), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT71), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT70), .B(G110), .Z(new_n538));
  OAI22_X1  g352(.A1(new_n531), .A2(new_n538), .B1(new_n524), .B2(new_n525), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n341), .A3(new_n368), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n536), .B2(new_n540), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n330), .A2(G221), .A3(G234), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT22), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(G137), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n541), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n536), .A2(new_n540), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n545), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n312), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT25), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n523), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(KEYINPUT72), .A3(new_n551), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT72), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n547), .A2(KEYINPUT71), .ZN(new_n555));
  INV_X1    g369(.A(new_n545), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(G902), .B1(new_n558), .B2(new_n548), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n554), .B1(new_n559), .B2(KEYINPUT25), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(KEYINPUT73), .A3(KEYINPUT25), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n552), .A2(new_n553), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n429), .B1(G234), .B2(new_n312), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n558), .A2(new_n548), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n563), .A2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT32), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT67), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n281), .B(new_n282), .C1(new_n476), .C2(new_n477), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT30), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n415), .A2(G137), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n471), .A2(G134), .ZN(new_n574));
  OAI21_X1  g388(.A(G131), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n275), .B(new_n575), .C1(G131), .C2(new_n475), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n571), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n572), .B1(new_n571), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n289), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n228), .B(new_n223), .Z(new_n580));
  NAND3_X1  g394(.A1(new_n571), .A2(new_n580), .A3(new_n576), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n333), .A2(G210), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n579), .A2(KEYINPUT31), .A3(new_n581), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n312), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n571), .A2(new_n580), .A3(new_n576), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n580), .B1(new_n571), .B2(new_n576), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT28), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT28), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n581), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n585), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT31), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n579), .A2(new_n581), .A3(new_n585), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n587), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(G472), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n570), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n586), .A2(new_n312), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n571), .A2(new_n576), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n289), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n591), .B1(new_n602), .B2(new_n581), .ZN(new_n603));
  INV_X1    g417(.A(new_n592), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n594), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT31), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n596), .ZN(new_n607));
  AND4_X1   g421(.A1(new_n570), .A2(new_n600), .A3(new_n607), .A4(new_n598), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n569), .B1(new_n599), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n600), .A2(new_n607), .A3(new_n598), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT29), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n590), .A2(new_n585), .A3(new_n592), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n579), .A2(new_n581), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n612), .B(new_n613), .C1(new_n615), .C2(new_n585), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n590), .A2(KEYINPUT29), .A3(new_n585), .A4(new_n592), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n617), .A2(KEYINPUT68), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(KEYINPUT68), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n616), .A2(new_n618), .A3(new_n312), .A4(new_n619), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n611), .A2(KEYINPUT32), .B1(new_n620), .B2(G472), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n568), .B1(new_n609), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n327), .A2(new_n461), .A3(new_n522), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  NOR2_X1   g438(.A1(new_n568), .A2(new_n463), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n610), .B(KEYINPUT67), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n600), .A2(new_n607), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(G472), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n516), .A2(new_n521), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n325), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n321), .B2(new_n323), .ZN(new_n633));
  INV_X1    g447(.A(new_n399), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n432), .A2(new_n433), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT100), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT33), .B1(new_n635), .B2(KEYINPUT100), .ZN(new_n639));
  OAI211_X1 g453(.A(G478), .B(new_n312), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n448), .A2(new_n400), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n634), .A2(new_n642), .A3(new_n457), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n631), .A2(new_n633), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n190), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n644), .B(new_n646), .ZN(G6));
  NAND2_X1  g461(.A1(new_n438), .A2(new_n450), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n634), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n457), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n631), .A2(new_n633), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n555), .A2(new_n557), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n556), .A2(KEYINPUT36), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n655), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n566), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n654), .B1(new_n564), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n659), .ZN(new_n661));
  AOI211_X1 g475(.A(KEYINPUT102), .B(new_n661), .C1(new_n562), .C2(new_n563), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n460), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n626), .ZN(new_n664));
  INV_X1    g478(.A(new_n628), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n327), .A2(new_n663), .A3(new_n522), .A4(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT37), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G110), .ZN(G12));
  INV_X1    g483(.A(new_n563), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT72), .B1(new_n550), .B2(new_n551), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n559), .A2(new_n554), .A3(KEYINPUT25), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND4_X1   g487(.A1(KEYINPUT73), .A2(new_n565), .A3(KEYINPUT25), .A4(new_n312), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT73), .B1(new_n559), .B2(KEYINPUT25), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n670), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT102), .B1(new_n677), .B2(new_n661), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT103), .B(G900), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(new_n443), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n441), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n634), .A2(new_n648), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n564), .A2(new_n654), .A3(new_n659), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n633), .A2(new_n678), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n609), .A2(new_n621), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n522), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n403), .ZN(G30));
  NAND2_X1  g502(.A1(new_n324), .A2(new_n326), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT38), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n660), .A2(new_n662), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n610), .A2(new_n569), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n626), .B2(new_n569), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n594), .B1(new_n588), .B2(new_n589), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n596), .A2(G472), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(G472), .A2(G902), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n694), .A2(KEYINPUT105), .A3(new_n699), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n681), .B(KEYINPUT39), .Z(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n706));
  NAND3_X1  g520(.A1(new_n522), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n702), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n706), .B1(new_n522), .B2(new_n705), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n399), .A2(new_n648), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n692), .A2(new_n325), .A3(new_n708), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  INV_X1    g527(.A(new_n681), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n634), .A2(new_n642), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n633), .A2(new_n678), .A3(new_n683), .A4(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n686), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n255), .ZN(G48));
  AND3_X1   g532(.A1(new_n514), .A2(new_n515), .A3(new_n312), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n515), .B1(new_n514), .B2(new_n312), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n719), .A2(new_n720), .A3(new_n463), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n721), .A2(new_n622), .A3(new_n633), .A4(new_n643), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n721), .A2(new_n622), .A3(new_n633), .A4(new_n650), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND4_X1  g540(.A1(new_n663), .A2(new_n685), .A3(new_n633), .A4(new_n721), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  NAND3_X1  g542(.A1(new_n628), .A2(KEYINPUT107), .A3(new_n610), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n627), .A2(new_n730), .A3(G472), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n562), .A2(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n732), .A2(new_n445), .A3(new_n733), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n632), .B(new_n710), .C1(new_n321), .C2(new_n323), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n721), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  NAND2_X1  g551(.A1(new_n514), .A2(new_n312), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(G469), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n462), .A3(new_n516), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n321), .A2(new_n323), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n325), .ZN(new_n742));
  INV_X1    g556(.A(new_n715), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT108), .B1(new_n691), .B2(new_n732), .ZN(new_n745));
  AND4_X1   g559(.A1(KEYINPUT108), .A2(new_n678), .A3(new_n683), .A4(new_n732), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  AOI21_X1  g562(.A(new_n632), .B1(new_n324), .B2(new_n326), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n522), .A3(new_n622), .A4(new_n715), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n610), .A2(new_n569), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n621), .A2(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n754), .A2(KEYINPUT42), .A3(new_n733), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n749), .A3(new_n522), .A4(new_n715), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G131), .ZN(G33));
  NAND4_X1  g572(.A1(new_n749), .A2(new_n522), .A3(new_n622), .A4(new_n682), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  INV_X1    g574(.A(new_n749), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n518), .A2(new_n467), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n496), .A2(new_n499), .A3(new_n467), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n520), .A2(KEYINPUT45), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(G469), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(G469), .A2(G902), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n719), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n768), .A2(KEYINPUT46), .A3(new_n769), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n462), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n762), .B1(new_n775), .B2(new_n704), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n463), .B1(new_n772), .B2(new_n773), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(KEYINPUT110), .A3(new_n705), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n761), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT43), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n642), .B2(new_n399), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n642), .A2(new_n399), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT43), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n666), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n691), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT44), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n779), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n775), .B2(KEYINPUT47), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n777), .A2(KEYINPUT111), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n775), .A2(KEYINPUT112), .A3(KEYINPUT47), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n777), .B2(new_n791), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n743), .A2(new_n685), .A3(new_n733), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n793), .A2(new_n797), .A3(new_n749), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  NOR2_X1   g614(.A1(new_n719), .A2(new_n720), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n782), .B1(new_n802), .B2(KEYINPUT49), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n632), .B(new_n803), .C1(KEYINPUT49), .C2(new_n802), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n702), .A2(new_n703), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n625), .A3(new_n690), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n522), .A2(new_n685), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n399), .A2(new_n648), .A3(new_n714), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n691), .A3(new_n749), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n745), .A2(new_n746), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n749), .A2(new_n522), .A3(new_n715), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n759), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n749), .A2(new_n522), .A3(new_n715), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n815), .A2(new_n755), .B1(new_n750), .B2(new_n751), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n686), .B1(new_n684), .B2(new_n716), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n678), .A2(new_n683), .A3(new_n732), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n691), .A2(KEYINPUT108), .A3(new_n732), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n818), .B1(new_n823), .B2(new_n744), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n714), .A2(KEYINPUT115), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n630), .A2(new_n463), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n564), .A2(new_n659), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n694), .B2(new_n699), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n714), .A2(KEYINPUT115), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n826), .A2(new_n828), .A3(new_n735), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n633), .A2(new_n678), .A3(new_n683), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n809), .B(new_n832), .C1(new_n682), .C2(new_n715), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n747), .A2(new_n830), .A3(new_n833), .A4(KEYINPUT52), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n817), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n722), .A2(new_n736), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(KEYINPUT113), .A3(new_n725), .A4(new_n727), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n727), .A2(new_n722), .A3(new_n725), .A4(new_n736), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n327), .A2(KEYINPUT114), .A3(new_n643), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n324), .A2(new_n326), .A3(new_n643), .A4(new_n325), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n843), .A2(new_n631), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n631), .A2(new_n327), .A3(new_n650), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n623), .A4(new_n667), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n842), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n808), .B1(new_n836), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n823), .A2(new_n815), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n757), .A2(new_n759), .A3(new_n811), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n747), .A2(new_n833), .A3(new_n830), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n854), .B1(new_n857), .B2(new_n834), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n849), .B1(new_n841), .B2(new_n838), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(KEYINPUT53), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n441), .B1(new_n783), .B2(new_n781), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n863), .A2(new_n733), .A3(new_n732), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n633), .A3(new_n721), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n808), .B1(new_n857), .B2(new_n834), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n849), .A2(new_n814), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n816), .B2(new_n839), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n816), .A2(new_n839), .A3(new_n869), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n867), .A2(new_n868), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n852), .A2(new_n866), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n330), .A2(G952), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n749), .A2(new_n721), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n805), .A2(new_n441), .A3(new_n568), .A4(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n634), .A2(new_n642), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n862), .A2(new_n865), .A3(new_n873), .A4(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n690), .A2(new_n632), .A3(new_n721), .A4(new_n864), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT50), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n749), .A2(new_n863), .A3(new_n721), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n823), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n876), .A2(new_n634), .A3(new_n642), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n793), .A2(new_n797), .B1(new_n463), .B2(new_n801), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n864), .A2(new_n749), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT117), .Z(new_n890));
  OR2_X1    g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT51), .B1(new_n887), .B2(new_n891), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n884), .A2(new_n733), .A3(new_n754), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT48), .Z(new_n897));
  NOR4_X1   g711(.A1(new_n879), .A2(new_n894), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(G952), .A2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n807), .B1(new_n898), .B2(new_n899), .ZN(G75));
  AOI21_X1  g714(.A(new_n312), .B1(new_n852), .B2(new_n872), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(G210), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n304), .A2(new_n306), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n309), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n902), .B2(new_n903), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n330), .A2(G952), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(G51));
  XOR2_X1   g724(.A(new_n769), .B(KEYINPUT57), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AND4_X1   g726(.A1(new_n867), .A2(new_n868), .A3(new_n870), .A4(new_n871), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT53), .B1(new_n858), .B2(new_n859), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT54), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n912), .B1(new_n915), .B2(new_n873), .ZN(new_n916));
  INV_X1    g730(.A(new_n514), .ZN(new_n917));
  OAI21_X1  g731(.A(KEYINPUT119), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n768), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n901), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n852), .A2(new_n866), .A3(new_n872), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n866), .B1(new_n852), .B2(new_n872), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n911), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n924), .A3(new_n514), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n918), .A2(new_n920), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n909), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(G54));
  AND2_X1   g742(.A1(new_n901), .A2(KEYINPUT58), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n391), .B1(new_n929), .B2(G475), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n909), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(G475), .A3(new_n391), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n929), .A2(KEYINPUT120), .A3(G475), .A4(new_n391), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n931), .A2(new_n934), .A3(new_n935), .ZN(G60));
  OR2_X1    g750(.A1(new_n638), .A2(new_n639), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n921), .B2(new_n922), .ZN(new_n938));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n862), .B2(new_n873), .ZN(new_n941));
  OAI221_X1 g755(.A(new_n927), .B1(new_n938), .B2(new_n940), .C1(new_n937), .C2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT60), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n852), .B2(new_n872), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n565), .B(KEYINPUT122), .ZN(new_n948));
  OR3_X1    g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n946), .B2(new_n948), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(KEYINPUT61), .A3(new_n927), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n658), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT121), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT121), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n946), .A2(new_n954), .A3(new_n658), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n927), .B1(new_n946), .B2(new_n948), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n953), .B2(new_n955), .ZN(new_n958));
  OAI22_X1  g772(.A1(new_n951), .A2(new_n956), .B1(new_n958), .B2(KEYINPUT61), .ZN(G66));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n330), .B1(new_n442), .B2(G224), .ZN(new_n961));
  AOI22_X1  g775(.A1(new_n851), .A2(new_n330), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n960), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n904), .B1(G898), .B2(new_n330), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(G69));
  NAND2_X1  g779(.A1(new_n787), .A2(new_n824), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n787), .A2(KEYINPUT127), .A3(new_n824), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n776), .A2(new_n778), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(new_n733), .A3(new_n735), .A4(new_n754), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n799), .A2(new_n757), .A3(new_n759), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n970), .A2(new_n330), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n577), .A2(new_n578), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(new_n387), .ZN(new_n976));
  NAND2_X1  g790(.A1(G900), .A2(G953), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT125), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n749), .A2(new_n522), .A3(new_n622), .ZN(new_n981));
  INV_X1    g795(.A(new_n877), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n704), .B1(new_n982), .B2(new_n649), .ZN(new_n983));
  AOI22_X1  g797(.A1(new_n779), .A2(new_n786), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n712), .A2(KEYINPUT62), .A3(new_n824), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT62), .B1(new_n712), .B2(new_n824), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n984), .B(new_n799), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n980), .B1(new_n987), .B2(new_n330), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n976), .A2(new_n979), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n988), .A2(KEYINPUT126), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT126), .B1(new_n988), .B2(new_n989), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n978), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n330), .B1(G227), .B2(G900), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n993), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n978), .B(new_n995), .C1(new_n990), .C2(new_n991), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(G72));
  XOR2_X1   g811(.A(new_n697), .B(KEYINPUT63), .Z(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n987), .B2(new_n851), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n614), .A3(new_n585), .ZN(new_n1000));
  INV_X1    g814(.A(new_n596), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n615), .A2(new_n585), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n861), .B(new_n998), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1000), .A2(new_n1003), .A3(new_n927), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n970), .A2(new_n859), .A3(new_n972), .A4(new_n973), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n585), .B1(new_n1005), .B2(new_n998), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1004), .B1(new_n615), .B2(new_n1006), .ZN(G57));
endmodule


