//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n462), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  INV_X1    g046(.A(new_n464), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n460), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OAI21_X1  g054(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g056(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n482));
  OAI221_X1 g057(.A(G2104), .B1(G112), .B2(new_n460), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT68), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(new_n474), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n465), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT66), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n491), .B(new_n492), .ZN(G162));
  NOR2_X1   g068(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n494), .B1(new_n474), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n498));
  INV_X1    g073(.A(new_n494), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n498), .A2(G138), .A3(new_n499), .A4(new_n495), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n465), .A2(G126), .A3(G2105), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G2104), .C1(G114), .C2(new_n460), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n497), .A2(new_n500), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT71), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n509), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(G543), .B1(new_n509), .B2(KEYINPUT5), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n514), .A2(new_n522), .ZN(G166));
  INV_X1    g098(.A(new_n518), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n526), .B(new_n528), .C1(new_n529), .C2(new_n520), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n513), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n518), .A2(new_n534), .B1(new_n520), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  AOI22_X1  g112(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n513), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT72), .B(G81), .Z(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n518), .A2(new_n540), .B1(new_n520), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT73), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n511), .A2(new_n550), .A3(new_n515), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n550), .B1(new_n511), .B2(new_n515), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G91), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n513), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(G166), .ZN(G303));
  INV_X1    g137(.A(G49), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n520), .A2(KEYINPUT75), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT75), .B1(new_n520), .B2(new_n563), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n511), .A2(G74), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n564), .A2(new_n565), .B1(G651), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n553), .A2(G87), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n518), .A2(KEYINPUT74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n511), .A2(new_n550), .A3(new_n515), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n570), .A2(G86), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n570), .A2(KEYINPUT76), .A3(G86), .A4(new_n571), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n577), .A2(new_n513), .B1(new_n578), .B2(new_n520), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT77), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  AOI211_X1 g157(.A(new_n582), .B(new_n579), .C1(new_n574), .C2(new_n575), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n513), .ZN(new_n586));
  INV_X1    g161(.A(new_n520), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n524), .A2(G85), .B1(new_n587), .B2(G47), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G54), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n591), .A2(new_n513), .B1(new_n592), .B2(new_n520), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n570), .A2(new_n571), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n553), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n590), .B1(new_n599), .B2(G868), .ZN(G321));
  XNOR2_X1  g175(.A(G321), .B(KEYINPUT78), .ZN(G284));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  INV_X1    g177(.A(G299), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G297));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  INV_X1    g182(.A(new_n543), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n597), .A2(new_n598), .ZN(new_n611));
  INV_X1    g186(.A(new_n593), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n610), .B1(new_n614), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n465), .A2(new_n470), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT80), .B(KEYINPUT13), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT81), .B(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT82), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n488), .A2(G123), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  INV_X1    g201(.A(G111), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n626), .A2(KEYINPUT83), .B1(new_n627), .B2(G2105), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(KEYINPUT83), .B2(new_n626), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n498), .A2(G135), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n625), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  OAI211_X1 g207(.A(new_n624), .B(new_n632), .C1(new_n622), .C2(new_n621), .ZN(G156));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT15), .B(G2435), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2430), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n645), .A2(new_n648), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n635), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G14), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n645), .A2(new_n648), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n645), .A2(new_n648), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n634), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT86), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n657));
  NAND4_X1  g232(.A1(new_n653), .A2(new_n657), .A3(new_n634), .A4(new_n654), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n652), .B1(new_n656), .B2(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT87), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n660), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n662), .A2(new_n664), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  MUX2_X1   g246(.A(new_n660), .B(new_n668), .S(new_n671), .Z(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(new_n673), .Z(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n676), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(new_n679), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT20), .Z(new_n683));
  AOI211_X1 g258(.A(new_n681), .B(new_n683), .C1(new_n676), .C2(new_n680), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT89), .ZN(new_n685));
  XOR2_X1   g260(.A(G1981), .B(G1986), .Z(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n685), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(G6), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G305), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT32), .B(G1981), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n697), .ZN(new_n699));
  NOR2_X1   g274(.A1(G16), .A2(G23), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT93), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G288), .B2(new_n693), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT33), .B(G1976), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT92), .B(G16), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n698), .A2(new_n699), .A3(new_n704), .A4(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G25), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT90), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n498), .A2(G131), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n460), .A2(G107), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  INV_X1    g294(.A(G119), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n717), .B1(new_n718), .B2(new_n719), .C1(new_n720), .C2(new_n487), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n716), .B1(new_n725), .B2(G29), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n706), .A2(G24), .ZN(new_n730));
  INV_X1    g305(.A(G290), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n706), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G1986), .Z(new_n733));
  NAND4_X1  g308(.A1(new_n712), .A2(new_n713), .A3(new_n729), .A4(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n705), .A2(G20), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT23), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n603), .B2(new_n693), .ZN(new_n739));
  INV_X1    g314(.A(G1956), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G4), .A2(G16), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n599), .B2(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G1348), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n706), .A2(G19), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n543), .B2(new_n706), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1341), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n498), .A2(G140), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n460), .A2(G116), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G128), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n748), .B1(new_n749), .B2(new_n750), .C1(new_n751), .C2(new_n487), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G29), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n714), .A2(G26), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT28), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2067), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n747), .A2(new_n757), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n741), .A2(new_n744), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT26), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n488), .B2(G129), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n498), .A2(G141), .B1(G105), .B2(new_n470), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT96), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G29), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G29), .B2(G32), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT31), .B(G11), .Z(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT30), .B(G28), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n714), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G34), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n774), .A2(KEYINPUT24), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(KEYINPUT24), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n478), .B2(G29), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT95), .B(G2084), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n773), .B1(new_n714), .B2(new_n631), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n780), .B2(new_n782), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n769), .A2(new_n770), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n693), .A2(G5), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G171), .B2(new_n693), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(G1961), .ZN(new_n788));
  NOR2_X1   g363(.A1(G168), .A2(new_n693), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n693), .B2(G21), .ZN(new_n790));
  INV_X1    g365(.A(G1966), .ZN(new_n791));
  INV_X1    g366(.A(G2078), .ZN(new_n792));
  NAND2_X1  g367(.A1(G164), .A2(G29), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G27), .B2(G29), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n790), .A2(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n790), .A2(new_n791), .B1(G1961), .B2(new_n787), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n714), .A2(G33), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n465), .A2(G127), .ZN(new_n798));
  NAND2_X1  g373(.A1(G115), .A2(G2104), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(G2105), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT25), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n804), .A2(new_n805), .B1(new_n498), .B2(G139), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n797), .B1(new_n808), .B2(new_n714), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT94), .B(G2072), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n794), .A2(new_n792), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n796), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n785), .A2(new_n788), .A3(new_n795), .A4(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT97), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n759), .B1(G1348), .B2(new_n743), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(G29), .A2(G35), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G162), .B2(G29), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT29), .Z(new_n819));
  INV_X1    g394(.A(G2090), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n819), .A2(new_n820), .B1(new_n814), .B2(new_n815), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n820), .B2(new_n819), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n736), .A2(new_n816), .A3(new_n822), .ZN(G311));
  OR3_X1    g398(.A1(new_n736), .A2(new_n816), .A3(new_n822), .ZN(G150));
  AOI22_X1  g399(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  OR3_X1    g400(.A1(new_n825), .A2(KEYINPUT98), .A3(new_n513), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT98), .B1(new_n825), .B2(new_n513), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n524), .A2(G93), .B1(new_n587), .B2(G55), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n599), .A2(G559), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT38), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n829), .A2(new_n608), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n543), .A2(new_n826), .A3(new_n827), .A4(new_n828), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n833), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT99), .ZN(new_n840));
  INV_X1    g415(.A(G860), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n838), .B2(KEYINPUT39), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n831), .B1(new_n840), .B2(new_n842), .ZN(G145));
  AOI22_X1  g418(.A1(new_n488), .A2(G130), .B1(G142), .B2(new_n498), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n460), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT100), .B1(G106), .B2(G2105), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n844), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n725), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n619), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n765), .A2(new_n807), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n752), .B(new_n504), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n808), .A2(new_n764), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n854), .B2(new_n856), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n853), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(G162), .A2(G160), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(G162), .A2(G160), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n631), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(G162), .A2(G160), .ZN(new_n865));
  INV_X1    g440(.A(new_n631), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n861), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n860), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n853), .A2(new_n859), .A3(KEYINPUT101), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT101), .B1(new_n853), .B2(new_n859), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n853), .A2(new_n859), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n864), .A2(new_n875), .A3(new_n867), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT102), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n860), .B2(new_n868), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n879), .B(new_n880), .C1(new_n876), .C2(new_n874), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n878), .A2(KEYINPUT40), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT40), .B1(new_n878), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(G395));
  NAND2_X1  g459(.A1(new_n829), .A2(new_n609), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n836), .B(new_n614), .Z(new_n886));
  NAND3_X1  g461(.A1(new_n613), .A2(KEYINPUT103), .A3(new_n603), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n599), .B2(G299), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n599), .A2(G299), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT104), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(KEYINPUT41), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n887), .A2(new_n889), .A3(new_n896), .A4(new_n890), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n886), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT76), .B1(new_n553), .B2(G86), .ZN(new_n900));
  INV_X1    g475(.A(new_n575), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n580), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n582), .ZN(new_n903));
  XNOR2_X1  g478(.A(G166), .B(KEYINPUT105), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n579), .B1(new_n574), .B2(new_n575), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT77), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n908));
  XNOR2_X1  g483(.A(G166), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n581), .B2(new_n583), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n731), .A2(new_n568), .A3(new_n567), .ZN(new_n911));
  NAND2_X1  g486(.A1(G288), .A2(G290), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n907), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n907), .A2(new_n910), .A3(KEYINPUT106), .A4(new_n913), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n907), .A2(new_n910), .ZN(new_n920));
  INV_X1    g495(.A(new_n913), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI211_X1 g497(.A(KEYINPUT107), .B(new_n913), .C1(new_n907), .C2(new_n910), .ZN(new_n923));
  OAI22_X1  g498(.A1(new_n916), .A2(new_n918), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT42), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n899), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n885), .B1(new_n926), .B2(new_n609), .ZN(G295));
  OAI21_X1  g502(.A(new_n885), .B1(new_n926), .B2(new_n609), .ZN(G331));
  NAND2_X1  g503(.A1(new_n920), .A2(new_n921), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT107), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n920), .A2(new_n919), .A3(new_n921), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n914), .A2(new_n915), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n930), .A2(new_n931), .B1(new_n932), .B2(new_n917), .ZN(new_n933));
  NAND2_X1  g508(.A1(G286), .A2(G171), .ZN(new_n934));
  NAND2_X1  g509(.A1(G301), .A2(G168), .ZN(new_n935));
  AND4_X1   g510(.A1(new_n834), .A2(new_n934), .A3(new_n835), .A4(new_n935), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n935), .A2(new_n934), .B1(new_n834), .B2(new_n835), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n895), .A2(new_n897), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n891), .B1(new_n936), .B2(new_n937), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n933), .A2(new_n943), .A3(new_n941), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n939), .A2(new_n940), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT108), .B1(new_n924), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n942), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n949), .B(new_n942), .C1(new_n944), .C2(new_n946), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(KEYINPUT109), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n953), .A3(KEYINPUT43), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n952), .B1(new_n947), .B2(KEYINPUT43), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n950), .A2(KEYINPUT110), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n950), .A2(KEYINPUT110), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(new_n959), .ZN(G397));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n504), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G40), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n468), .A2(new_n476), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(G1996), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT46), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT125), .ZN(new_n968));
  INV_X1    g543(.A(G2067), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n752), .B(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT112), .ZN(new_n971));
  INV_X1    g546(.A(new_n764), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n965), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n966), .A2(KEYINPUT46), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n968), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n975), .B(KEYINPUT47), .Z(new_n976));
  INV_X1    g551(.A(G1996), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n971), .A2(new_n977), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n973), .A2(new_n978), .B1(new_n765), .B2(new_n966), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n725), .A2(new_n728), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT124), .Z(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(G2067), .B2(new_n752), .ZN(new_n983));
  INV_X1    g558(.A(new_n965), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n727), .B1(new_n723), .B2(new_n724), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n984), .B1(new_n980), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n979), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n965), .A2(G1986), .A3(G290), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT48), .Z(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n976), .A2(new_n985), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT126), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n992), .B(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(G303), .A2(G8), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT55), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n504), .A2(new_n998), .A3(new_n961), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n504), .B2(new_n961), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n469), .A2(G40), .A3(new_n477), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n820), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n504), .A2(new_n961), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n964), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(new_n962), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n709), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1004), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT113), .B1(new_n1009), .B2(new_n709), .ZN(new_n1013));
  OAI211_X1 g588(.A(G8), .B(new_n997), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT114), .B(G1981), .Z(new_n1016));
  NAND2_X1  g591(.A1(new_n905), .A2(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n524), .A2(G86), .ZN(new_n1018));
  OAI21_X1  g593(.A(G1981), .B1(new_n579), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT49), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(G8), .B1(new_n1005), .B2(new_n1002), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1017), .A2(new_n1019), .A3(KEYINPUT49), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G288), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1021), .B1(new_n1025), .B2(G1976), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1026), .B(new_n1027), .C1(G1976), .C2(new_n1025), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1024), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1024), .A2(new_n1031), .A3(new_n1025), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1017), .ZN(new_n1033));
  XOR2_X1   g608(.A(new_n1021), .B(KEYINPUT115), .Z(new_n1034));
  AOI22_X1  g609(.A1(new_n1015), .A2(new_n1030), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1010), .A2(new_n1004), .ZN(new_n1036));
  INV_X1    g611(.A(G8), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n996), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1030), .A2(new_n1014), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1005), .A2(KEYINPUT50), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1041), .A2(new_n964), .A3(new_n999), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n1043));
  OR3_X1    g618(.A1(new_n1042), .A2(new_n1043), .A3(G2084), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1042), .B2(G2084), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1044), .B(new_n1045), .C1(G1966), .C2(new_n1008), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1046), .A2(G8), .A3(G168), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT63), .B1(new_n1040), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(G8), .A3(G168), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT63), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n996), .ZN(new_n1053));
  AND4_X1   g628(.A1(new_n1014), .A2(new_n1051), .A3(new_n1053), .A4(new_n1030), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1035), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G168), .A2(new_n1037), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n1046), .B2(G8), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1047), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1046), .A2(new_n1057), .A3(G8), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1056), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT51), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT62), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n1009), .B2(G2078), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1008), .A2(KEYINPUT53), .A3(new_n792), .ZN(new_n1068));
  OR2_X1    g643(.A1(new_n1003), .A2(G1961), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1042), .A2(G2084), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1073), .A2(new_n1043), .B1(new_n1009), .B2(new_n791), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1037), .B1(new_n1074), .B2(new_n1044), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1049), .B1(new_n1075), .B2(new_n1059), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1056), .B1(new_n1075), .B2(new_n1057), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1076), .B(new_n1077), .C1(new_n1078), .C2(KEYINPUT51), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1065), .A2(new_n1072), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1003), .B2(G1956), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1042), .A2(KEYINPUT117), .A3(new_n740), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT56), .B(G2072), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1082), .A2(new_n1083), .B1(new_n1008), .B2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(G299), .B(KEYINPUT57), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT119), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n964), .A2(new_n961), .A3(new_n969), .A4(new_n504), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(KEYINPUT118), .ZN(new_n1090));
  INV_X1    g665(.A(G1348), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1042), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n613), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1008), .A2(new_n1084), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1042), .A2(KEYINPUT117), .A3(new_n740), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT117), .B1(new_n1042), .B2(new_n740), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n1086), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1088), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1087), .B(new_n1095), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1098), .A2(new_n1086), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1102), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT122), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n1108), .B(KEYINPUT61), .C1(new_n1104), .C2(new_n1102), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT120), .B(G1996), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1007), .A2(new_n962), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1005), .A2(new_n1002), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT58), .B(G1341), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n543), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n1117));
  NAND2_X1  g692(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n543), .B(new_n1118), .C1(new_n1112), .C2(new_n1115), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1090), .A2(new_n613), .A3(new_n1092), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT60), .B1(new_n1121), .B2(new_n1093), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n613), .A2(KEYINPUT60), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1090), .A2(new_n1123), .A3(new_n1092), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1085), .A2(KEYINPUT119), .A3(new_n1087), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1099), .B1(new_n1098), .B2(new_n1086), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1106), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1125), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1103), .B1(new_n1110), .B2(new_n1130), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1070), .A2(G171), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1132), .A2(new_n1071), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n1132), .B2(new_n1071), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n1134), .A2(new_n1135), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1080), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1055), .B1(new_n1137), .B2(new_n1040), .ZN(new_n1138));
  AND2_X1   g713(.A1(G290), .A2(G1986), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n989), .B1(new_n984), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT111), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n988), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n994), .B1(new_n1138), .B2(new_n1142), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n1145));
  OR2_X1    g719(.A1(G227), .A2(new_n458), .ZN(new_n1146));
  OAI21_X1  g720(.A(new_n1145), .B1(G401), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g721(.A1(G227), .A2(new_n458), .ZN(new_n1148));
  AND2_X1   g722(.A1(new_n656), .A2(new_n658), .ZN(new_n1149));
  OAI211_X1 g723(.A(KEYINPUT127), .B(new_n1148), .C1(new_n1149), .C2(new_n652), .ZN(new_n1150));
  NAND3_X1  g724(.A1(new_n1147), .A2(new_n1150), .A3(new_n691), .ZN(new_n1151));
  AOI21_X1  g725(.A(new_n1151), .B1(new_n878), .B2(new_n881), .ZN(new_n1152));
  AND3_X1   g726(.A1(new_n1152), .A2(new_n951), .A3(new_n954), .ZN(G308));
  NAND3_X1  g727(.A1(new_n1152), .A2(new_n954), .A3(new_n951), .ZN(G225));
endmodule


