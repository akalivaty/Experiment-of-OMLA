

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593;

  XNOR2_X1 U324 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n379) );
  XNOR2_X1 U325 ( .A(n464), .B(n463), .ZN(n533) );
  INV_X1 U326 ( .A(KEYINPUT73), .ZN(n306) );
  XOR2_X1 U327 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n368) );
  XOR2_X1 U328 ( .A(G85GAT), .B(G57GAT), .Z(n438) );
  XNOR2_X1 U329 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U330 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U331 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U332 ( .A(n380), .B(n379), .ZN(n387) );
  OR2_X1 U333 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U334 ( .A(n455), .B(n454), .ZN(n458) );
  NOR2_X1 U335 ( .A1(n476), .A2(n579), .ZN(n550) );
  XNOR2_X1 U336 ( .A(n462), .B(n461), .ZN(n463) );
  NOR2_X1 U337 ( .A1(n465), .A2(n525), .ZN(n571) );
  XNOR2_X1 U338 ( .A(n499), .B(KEYINPUT38), .ZN(n505) );
  XNOR2_X1 U339 ( .A(n466), .B(G190GAT), .ZN(n467) );
  XNOR2_X1 U340 ( .A(n468), .B(n467), .ZN(G1351GAT) );
  XOR2_X1 U341 ( .A(G92GAT), .B(G64GAT), .Z(n292) );
  XOR2_X1 U342 ( .A(G204GAT), .B(n292), .Z(n397) );
  XOR2_X1 U343 ( .A(KEYINPUT33), .B(G176GAT), .Z(n294) );
  XNOR2_X1 U344 ( .A(n438), .B(n368), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U346 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n296) );
  XNOR2_X1 U347 ( .A(KEYINPUT75), .B(KEYINPUT31), .ZN(n295) );
  XOR2_X1 U348 ( .A(n296), .B(n295), .Z(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n299) );
  NAND2_X1 U350 ( .A1(G230GAT), .A2(G233GAT), .ZN(n300) );
  NAND2_X1 U351 ( .A1(n299), .A2(n300), .ZN(n304) );
  INV_X1 U352 ( .A(n299), .ZN(n302) );
  INV_X1 U353 ( .A(n300), .ZN(n301) );
  NAND2_X1 U354 ( .A1(n302), .A2(n301), .ZN(n303) );
  NAND2_X1 U355 ( .A1(n304), .A2(n303), .ZN(n309) );
  XNOR2_X1 U356 ( .A(G148GAT), .B(G106GAT), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n305), .B(G78GAT), .ZN(n410) );
  XNOR2_X1 U358 ( .A(n410), .B(KEYINPUT76), .ZN(n307) );
  XOR2_X1 U359 ( .A(n397), .B(n310), .Z(n316) );
  INV_X1 U360 ( .A(G99GAT), .ZN(n311) );
  NAND2_X1 U361 ( .A1(G120GAT), .A2(n311), .ZN(n314) );
  INV_X1 U362 ( .A(G120GAT), .ZN(n312) );
  NAND2_X1 U363 ( .A1(n312), .A2(G99GAT), .ZN(n313) );
  NAND2_X1 U364 ( .A1(n314), .A2(n313), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n315), .B(G71GAT), .ZN(n451) );
  XNOR2_X1 U366 ( .A(n316), .B(n451), .ZN(n383) );
  XOR2_X1 U367 ( .A(KEYINPUT64), .B(KEYINPUT41), .Z(n317) );
  XNOR2_X1 U368 ( .A(n383), .B(n317), .ZN(n507) );
  XOR2_X1 U369 ( .A(G36GAT), .B(G8GAT), .Z(n403) );
  XOR2_X1 U370 ( .A(G197GAT), .B(n403), .Z(n319) );
  XOR2_X1 U371 ( .A(G1GAT), .B(KEYINPUT70), .Z(n367) );
  XNOR2_X1 U372 ( .A(G15GAT), .B(n367), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n325) );
  XOR2_X1 U374 ( .A(G141GAT), .B(G22GAT), .Z(n411) );
  XOR2_X1 U375 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n321) );
  XNOR2_X1 U376 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n340) );
  XOR2_X1 U378 ( .A(n411), .B(n340), .Z(n323) );
  NAND2_X1 U379 ( .A1(G229GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U381 ( .A(n325), .B(n324), .Z(n327) );
  XNOR2_X1 U382 ( .A(G50GAT), .B(G43GAT), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n335) );
  XOR2_X1 U384 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n329) );
  XNOR2_X1 U385 ( .A(G113GAT), .B(G169GAT), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U387 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n331) );
  XNOR2_X1 U388 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(n333), .B(n332), .Z(n334) );
  XOR2_X1 U391 ( .A(n335), .B(n334), .Z(n535) );
  INV_X1 U392 ( .A(n535), .ZN(n580) );
  NAND2_X1 U393 ( .A1(n507), .A2(n580), .ZN(n336) );
  XNOR2_X1 U394 ( .A(KEYINPUT46), .B(n336), .ZN(n378) );
  XOR2_X1 U395 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n338) );
  XNOR2_X1 U396 ( .A(G218GAT), .B(KEYINPUT78), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U398 ( .A(G134GAT), .B(G43GAT), .Z(n450) );
  XOR2_X1 U399 ( .A(n339), .B(n450), .Z(n345) );
  XOR2_X1 U400 ( .A(n340), .B(G85GAT), .Z(n342) );
  NAND2_X1 U401 ( .A1(G232GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U403 ( .A(G162GAT), .B(G50GAT), .Z(n416) );
  XNOR2_X1 U404 ( .A(n343), .B(n416), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n353) );
  XOR2_X1 U406 ( .A(G92GAT), .B(G190GAT), .Z(n347) );
  XNOR2_X1 U407 ( .A(KEYINPUT65), .B(KEYINPUT79), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U409 ( .A(G99GAT), .B(G106GAT), .Z(n349) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(KEYINPUT11), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U412 ( .A(n351), .B(n350), .Z(n352) );
  XOR2_X1 U413 ( .A(n353), .B(n352), .Z(n544) );
  INV_X1 U414 ( .A(n544), .ZN(n562) );
  XOR2_X1 U415 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n355) );
  XNOR2_X1 U416 ( .A(KEYINPUT14), .B(KEYINPUT80), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n376) );
  XOR2_X1 U418 ( .A(G64GAT), .B(G183GAT), .Z(n357) );
  XNOR2_X1 U419 ( .A(G57GAT), .B(G71GAT), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U421 ( .A(KEYINPUT83), .B(KEYINPUT12), .Z(n359) );
  XNOR2_X1 U422 ( .A(KEYINPUT85), .B(G8GAT), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U424 ( .A(n361), .B(n360), .Z(n366) );
  XOR2_X1 U425 ( .A(G127GAT), .B(G15GAT), .Z(n460) );
  XOR2_X1 U426 ( .A(KEYINPUT82), .B(KEYINPUT84), .Z(n363) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n460), .B(n364), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n372) );
  XOR2_X1 U431 ( .A(G22GAT), .B(G211GAT), .Z(n370) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U434 ( .A(n372), .B(n371), .Z(n374) );
  XNOR2_X1 U435 ( .A(G155GAT), .B(G78GAT), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U437 ( .A(n376), .B(n375), .Z(n541) );
  INV_X1 U438 ( .A(n541), .ZN(n587) );
  NOR2_X1 U439 ( .A1(n562), .A2(n587), .ZN(n377) );
  NAND2_X1 U440 ( .A1(n378), .A2(n377), .ZN(n380) );
  XOR2_X1 U441 ( .A(KEYINPUT36), .B(n544), .Z(n590) );
  NAND2_X1 U442 ( .A1(n587), .A2(n590), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n381), .B(KEYINPUT111), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n382), .B(KEYINPUT45), .ZN(n384) );
  INV_X1 U445 ( .A(n383), .ZN(n583) );
  NAND2_X1 U446 ( .A1(n384), .A2(n583), .ZN(n385) );
  NOR2_X1 U447 ( .A1(n580), .A2(n385), .ZN(n386) );
  NOR2_X1 U448 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n388), .B(KEYINPUT48), .ZN(n553) );
  XOR2_X1 U450 ( .A(G176GAT), .B(KEYINPUT17), .Z(n390) );
  XNOR2_X1 U451 ( .A(G183GAT), .B(KEYINPUT88), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U453 ( .A(KEYINPUT89), .B(KEYINPUT18), .Z(n392) );
  XNOR2_X1 U454 ( .A(G190GAT), .B(KEYINPUT90), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U456 ( .A(n394), .B(n393), .Z(n396) );
  XNOR2_X1 U457 ( .A(KEYINPUT19), .B(G169GAT), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n462) );
  XOR2_X1 U459 ( .A(n462), .B(n397), .Z(n407) );
  XOR2_X1 U460 ( .A(G197GAT), .B(KEYINPUT21), .Z(n399) );
  XNOR2_X1 U461 ( .A(G218GAT), .B(G211GAT), .ZN(n398) );
  XNOR2_X1 U462 ( .A(n399), .B(n398), .ZN(n422) );
  XOR2_X1 U463 ( .A(n422), .B(KEYINPUT100), .Z(n401) );
  NAND2_X1 U464 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U466 ( .A(n402), .B(KEYINPUT99), .Z(n405) );
  XNOR2_X1 U467 ( .A(n403), .B(KEYINPUT101), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U469 ( .A(n407), .B(n406), .Z(n488) );
  XNOR2_X1 U470 ( .A(KEYINPUT117), .B(n488), .ZN(n408) );
  NOR2_X1 U471 ( .A1(n553), .A2(n408), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n409), .B(KEYINPUT54), .ZN(n577) );
  XOR2_X1 U473 ( .A(KEYINPUT22), .B(n410), .Z(n415) );
  XNOR2_X1 U474 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n412) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U476 ( .A(G204GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n419) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U480 ( .A(n419), .B(n418), .Z(n424) );
  XOR2_X1 U481 ( .A(G155GAT), .B(KEYINPUT2), .Z(n421) );
  XNOR2_X1 U482 ( .A(KEYINPUT3), .B(KEYINPUT94), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n426), .B(n422), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n474) );
  XNOR2_X1 U486 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n425), .B(KEYINPUT86), .ZN(n456) );
  XNOR2_X1 U488 ( .A(n426), .B(n456), .ZN(n446) );
  XOR2_X1 U489 ( .A(KEYINPUT5), .B(G120GAT), .Z(n428) );
  XNOR2_X1 U490 ( .A(G141GAT), .B(G127GAT), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U492 ( .A(G1GAT), .B(KEYINPUT97), .Z(n430) );
  XNOR2_X1 U493 ( .A(KEYINPUT4), .B(KEYINPUT98), .ZN(n429) );
  XNOR2_X1 U494 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U495 ( .A(n432), .B(n431), .Z(n444) );
  XOR2_X1 U496 ( .A(KEYINPUT96), .B(KEYINPUT1), .Z(n434) );
  XNOR2_X1 U497 ( .A(KEYINPUT6), .B(KEYINPUT95), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n442) );
  XOR2_X1 U499 ( .A(G148GAT), .B(G134GAT), .Z(n436) );
  XNOR2_X1 U500 ( .A(G29GAT), .B(G162GAT), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U502 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U503 ( .A1(G225GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U506 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U507 ( .A(n446), .B(n445), .Z(n576) );
  INV_X1 U508 ( .A(n576), .ZN(n551) );
  NOR2_X1 U509 ( .A1(n474), .A2(n551), .ZN(n447) );
  AND2_X1 U510 ( .A1(n577), .A2(n447), .ZN(n449) );
  XNOR2_X1 U511 ( .A(KEYINPUT118), .B(KEYINPUT55), .ZN(n448) );
  XNOR2_X1 U512 ( .A(n449), .B(n448), .ZN(n465) );
  XNOR2_X1 U513 ( .A(n451), .B(n450), .ZN(n455) );
  NAND2_X1 U514 ( .A1(G227GAT), .A2(G233GAT), .ZN(n453) );
  INV_X1 U515 ( .A(KEYINPUT87), .ZN(n452) );
  XNOR2_X1 U516 ( .A(n456), .B(KEYINPUT20), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U518 ( .A(KEYINPUT91), .B(n459), .Z(n464) );
  XNOR2_X1 U519 ( .A(n460), .B(KEYINPUT92), .ZN(n461) );
  INV_X1 U520 ( .A(n533), .ZN(n525) );
  NAND2_X1 U521 ( .A1(n571), .A2(n562), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n466) );
  XNOR2_X1 U523 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n487) );
  NAND2_X1 U524 ( .A1(n583), .A2(n580), .ZN(n469) );
  XNOR2_X1 U525 ( .A(KEYINPUT77), .B(n469), .ZN(n498) );
  XOR2_X1 U526 ( .A(KEYINPUT27), .B(n488), .Z(n476) );
  XOR2_X1 U527 ( .A(n474), .B(KEYINPUT28), .Z(n529) );
  INV_X1 U528 ( .A(n529), .ZN(n492) );
  NOR2_X1 U529 ( .A1(n476), .A2(n492), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n551), .A2(n470), .ZN(n532) );
  XOR2_X1 U531 ( .A(KEYINPUT93), .B(n533), .Z(n471) );
  NOR2_X1 U532 ( .A1(n532), .A2(n471), .ZN(n482) );
  INV_X1 U533 ( .A(n488), .ZN(n523) );
  NOR2_X1 U534 ( .A1(n523), .A2(n525), .ZN(n472) );
  NOR2_X1 U535 ( .A1(n474), .A2(n472), .ZN(n473) );
  XOR2_X1 U536 ( .A(KEYINPUT25), .B(n473), .Z(n478) );
  NAND2_X1 U537 ( .A1(n474), .A2(n525), .ZN(n475) );
  XNOR2_X1 U538 ( .A(KEYINPUT26), .B(n475), .ZN(n579) );
  XNOR2_X1 U539 ( .A(n550), .B(KEYINPUT102), .ZN(n477) );
  NOR2_X1 U540 ( .A1(n478), .A2(n477), .ZN(n479) );
  NOR2_X1 U541 ( .A1(n551), .A2(n479), .ZN(n480) );
  XOR2_X1 U542 ( .A(KEYINPUT103), .B(n480), .Z(n481) );
  NOR2_X1 U543 ( .A1(n482), .A2(n481), .ZN(n496) );
  NOR2_X1 U544 ( .A1(n541), .A2(n562), .ZN(n483) );
  XOR2_X1 U545 ( .A(KEYINPUT16), .B(n483), .Z(n484) );
  NOR2_X1 U546 ( .A1(n496), .A2(n484), .ZN(n509) );
  NAND2_X1 U547 ( .A1(n498), .A2(n509), .ZN(n485) );
  XOR2_X1 U548 ( .A(KEYINPUT104), .B(n485), .Z(n493) );
  NAND2_X1 U549 ( .A1(n551), .A2(n493), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U551 ( .A1(n493), .A2(n488), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .Z(n491) );
  NAND2_X1 U554 ( .A1(n493), .A2(n533), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  NAND2_X1 U556 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n494), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U558 ( .A1(n541), .A2(n590), .ZN(n495) );
  XNOR2_X1 U559 ( .A(KEYINPUT37), .B(n497), .ZN(n519) );
  NAND2_X1 U560 ( .A1(n498), .A2(n519), .ZN(n499) );
  NOR2_X1 U561 ( .A1(n505), .A2(n576), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(n500), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(KEYINPUT39), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n505), .A2(n523), .ZN(n502) );
  XOR2_X1 U565 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U566 ( .A1(n505), .A2(n525), .ZN(n503) );
  XOR2_X1 U567 ( .A(KEYINPUT40), .B(n503), .Z(n504) );
  XNOR2_X1 U568 ( .A(n504), .B(G43GAT), .ZN(G1330GAT) );
  NOR2_X1 U569 ( .A1(n529), .A2(n505), .ZN(n506) );
  XOR2_X1 U570 ( .A(G50GAT), .B(n506), .Z(G1331GAT) );
  NAND2_X1 U571 ( .A1(n507), .A2(n535), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n508), .B(KEYINPUT105), .ZN(n520) );
  NAND2_X1 U573 ( .A1(n509), .A2(n520), .ZN(n516) );
  NOR2_X1 U574 ( .A1(n576), .A2(n516), .ZN(n510) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n510), .Z(n511) );
  XNOR2_X1 U576 ( .A(KEYINPUT42), .B(n511), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n523), .A2(n516), .ZN(n512) );
  XOR2_X1 U578 ( .A(KEYINPUT106), .B(n512), .Z(n513) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n513), .ZN(G1333GAT) );
  NOR2_X1 U580 ( .A1(n525), .A2(n516), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U583 ( .A1(n529), .A2(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n520), .ZN(n528) );
  NOR2_X1 U587 ( .A1(n576), .A2(n528), .ZN(n521) );
  XOR2_X1 U588 ( .A(KEYINPUT108), .B(n521), .Z(n522) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n528), .ZN(n524) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n528), .ZN(n527) );
  XNOR2_X1 U593 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(G1338GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(n530), .Z(n531) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n532), .A2(n553), .ZN(n534) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n545) );
  NOR2_X1 U600 ( .A1(n535), .A2(n545), .ZN(n536) );
  XOR2_X1 U601 ( .A(KEYINPUT112), .B(n536), .Z(n537) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  INV_X1 U603 ( .A(n507), .ZN(n538) );
  NOR2_X1 U604 ( .A1(n538), .A2(n545), .ZN(n540) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NOR2_X1 U607 ( .A1(n541), .A2(n545), .ZN(n542) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(n542), .Z(n543) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  NOR2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n547) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT114), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  XOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT115), .Z(n555) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n561), .A2(n580), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n555), .B(n554), .ZN(G1344GAT) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U622 ( .A1(n561), .A2(n507), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n587), .A2(n561), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT119), .Z(n565) );
  NAND2_X1 U630 ( .A1(n571), .A2(n580), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n567) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT120), .B(n568), .Z(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n507), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n587), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(KEYINPUT122), .ZN(n573) );
  XNOR2_X1 U640 ( .A(G183GAT), .B(n573), .ZN(G1350GAT) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(KEYINPUT60), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT59), .B(n575), .Z(n582) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n591) );
  NAND2_X1 U646 ( .A1(n591), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U649 ( .A1(n591), .A2(n383), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(G204GAT), .B(n586), .Z(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n591), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(KEYINPUT126), .ZN(n589) );
  XNOR2_X1 U654 ( .A(G211GAT), .B(n589), .ZN(G1354GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n592), .B(KEYINPUT62), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

