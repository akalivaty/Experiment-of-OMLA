

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U319 ( .A(n366), .B(n365), .ZN(n367) );
  AND2_X1 U320 ( .A1(G230GAT), .A2(G233GAT), .ZN(n287) );
  AND2_X1 U321 ( .A1(G232GAT), .A2(G233GAT), .ZN(n288) );
  XOR2_X1 U322 ( .A(n382), .B(n381), .Z(n289) );
  XNOR2_X1 U323 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n394) );
  XNOR2_X1 U324 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U325 ( .A(G50GAT), .B(G162GAT), .Z(n434) );
  XNOR2_X1 U326 ( .A(n376), .B(n288), .ZN(n360) );
  XNOR2_X1 U327 ( .A(n376), .B(n287), .ZN(n377) );
  XNOR2_X1 U328 ( .A(n361), .B(n360), .ZN(n363) );
  XNOR2_X1 U329 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U330 ( .A(n383), .B(n289), .ZN(n384) );
  XNOR2_X1 U331 ( .A(n368), .B(n367), .ZN(n371) );
  XNOR2_X1 U332 ( .A(n385), .B(n384), .ZN(n389) );
  XNOR2_X1 U333 ( .A(KEYINPUT97), .B(n458), .ZN(n563) );
  XNOR2_X1 U334 ( .A(n448), .B(G134GAT), .ZN(n449) );
  XNOR2_X1 U335 ( .A(n450), .B(n449), .ZN(G1343GAT) );
  XNOR2_X1 U336 ( .A(KEYINPUT27), .B(KEYINPUT98), .ZN(n307) );
  XOR2_X1 U337 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n291) );
  XNOR2_X1 U338 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n290) );
  XNOR2_X1 U339 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U340 ( .A(n292), .B(KEYINPUT84), .Z(n294) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(G183GAT), .ZN(n293) );
  XNOR2_X1 U342 ( .A(n294), .B(n293), .ZN(n311) );
  XNOR2_X1 U343 ( .A(G211GAT), .B(KEYINPUT87), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n295), .B(KEYINPUT21), .ZN(n296) );
  XOR2_X1 U345 ( .A(n296), .B(KEYINPUT86), .Z(n298) );
  XNOR2_X1 U346 ( .A(G197GAT), .B(G204GAT), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n441) );
  XNOR2_X1 U348 ( .A(G176GAT), .B(G64GAT), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n299), .B(KEYINPUT72), .ZN(n387) );
  XNOR2_X1 U350 ( .A(n441), .B(n387), .ZN(n305) );
  XOR2_X1 U351 ( .A(G92GAT), .B(G218GAT), .Z(n301) );
  XNOR2_X1 U352 ( .A(G36GAT), .B(G190GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n365) );
  XOR2_X1 U354 ( .A(n365), .B(G8GAT), .Z(n303) );
  NAND2_X1 U355 ( .A1(G226GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n311), .B(n306), .ZN(n540) );
  XNOR2_X1 U359 ( .A(n307), .B(n540), .ZN(n459) );
  XOR2_X1 U360 ( .A(G127GAT), .B(G71GAT), .Z(n309) );
  XNOR2_X1 U361 ( .A(G15GAT), .B(G120GAT), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n325) );
  XOR2_X1 U364 ( .A(G176GAT), .B(KEYINPUT80), .Z(n313) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(G190GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U367 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n315) );
  XNOR2_X1 U368 ( .A(KEYINPUT81), .B(KEYINPUT85), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U370 ( .A(n317), .B(n316), .Z(n323) );
  XNOR2_X1 U371 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n318), .B(KEYINPUT79), .ZN(n423) );
  XOR2_X1 U373 ( .A(G99GAT), .B(n423), .Z(n320) );
  NAND2_X1 U374 ( .A1(G227GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U376 ( .A(G134GAT), .B(n321), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n547) );
  XOR2_X1 U379 ( .A(KEYINPUT64), .B(KEYINPUT66), .Z(n327) );
  XNOR2_X1 U380 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n344) );
  XOR2_X1 U382 ( .A(G36GAT), .B(G50GAT), .Z(n329) );
  XNOR2_X1 U383 ( .A(G169GAT), .B(G29GAT), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U385 ( .A(G1GAT), .B(G141GAT), .Z(n331) );
  XNOR2_X1 U386 ( .A(G113GAT), .B(G197GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U388 ( .A(n333), .B(n332), .Z(n342) );
  XOR2_X1 U389 ( .A(G22GAT), .B(G15GAT), .Z(n335) );
  XNOR2_X1 U390 ( .A(KEYINPUT68), .B(G8GAT), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U392 ( .A(KEYINPUT67), .B(n336), .Z(n354) );
  XNOR2_X1 U393 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n337), .B(KEYINPUT7), .ZN(n369) );
  XOR2_X1 U395 ( .A(n369), .B(KEYINPUT65), .Z(n339) );
  NAND2_X1 U396 ( .A1(G229GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n354), .B(n340), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U400 ( .A(n344), .B(n343), .Z(n567) );
  INV_X1 U401 ( .A(n567), .ZN(n516) );
  XOR2_X1 U402 ( .A(KEYINPUT12), .B(G64GAT), .Z(n346) );
  XNOR2_X1 U403 ( .A(G155GAT), .B(G57GAT), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n358) );
  XNOR2_X1 U405 ( .A(G71GAT), .B(G78GAT), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n347), .B(KEYINPUT13), .ZN(n386) );
  XOR2_X1 U407 ( .A(G1GAT), .B(G127GAT), .Z(n407) );
  XOR2_X1 U408 ( .A(n386), .B(n407), .Z(n349) );
  XNOR2_X1 U409 ( .A(G183GAT), .B(G211GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U411 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n351) );
  NAND2_X1 U412 ( .A1(G231GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U414 ( .A(n353), .B(n352), .Z(n356) );
  XNOR2_X1 U415 ( .A(n354), .B(KEYINPUT77), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U417 ( .A(n358), .B(n357), .Z(n574) );
  XNOR2_X1 U418 ( .A(n434), .B(KEYINPUT9), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n359), .B(KEYINPUT11), .ZN(n361) );
  XOR2_X1 U420 ( .A(G99GAT), .B(G106GAT), .Z(n376) );
  INV_X1 U421 ( .A(KEYINPUT10), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n368) );
  XNOR2_X1 U423 ( .A(G29GAT), .B(G134GAT), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n364), .B(G85GAT), .ZN(n415) );
  XNOR2_X1 U425 ( .A(n415), .B(KEYINPUT75), .ZN(n366) );
  INV_X1 U426 ( .A(n369), .ZN(n370) );
  XOR2_X1 U427 ( .A(n371), .B(n370), .Z(n536) );
  INV_X1 U428 ( .A(KEYINPUT76), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n536), .B(n372), .ZN(n446) );
  XNOR2_X1 U430 ( .A(n446), .B(KEYINPUT36), .ZN(n476) );
  NOR2_X1 U431 ( .A1(n574), .A2(n476), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n373), .B(KEYINPUT45), .ZN(n390) );
  XOR2_X1 U433 ( .A(KEYINPUT70), .B(G92GAT), .Z(n375) );
  XNOR2_X1 U434 ( .A(G204GAT), .B(G85GAT), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n378) );
  XOR2_X1 U436 ( .A(n379), .B(KEYINPUT69), .Z(n385) );
  XOR2_X1 U437 ( .A(G120GAT), .B(G148GAT), .Z(n380) );
  XOR2_X1 U438 ( .A(G57GAT), .B(n380), .Z(n424) );
  XNOR2_X1 U439 ( .A(n424), .B(KEYINPUT71), .ZN(n383) );
  XOR2_X1 U440 ( .A(KEYINPUT31), .B(KEYINPUT73), .Z(n382) );
  XNOR2_X1 U441 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n389), .B(n388), .ZN(n571) );
  NAND2_X1 U444 ( .A1(n390), .A2(n571), .ZN(n392) );
  INV_X1 U445 ( .A(KEYINPUT111), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  NOR2_X1 U447 ( .A1(n516), .A2(n393), .ZN(n400) );
  XNOR2_X1 U448 ( .A(n571), .B(KEYINPUT41), .ZN(n518) );
  NAND2_X1 U449 ( .A1(n518), .A2(n516), .ZN(n395) );
  NAND2_X1 U450 ( .A1(n396), .A2(n574), .ZN(n397) );
  NOR2_X1 U451 ( .A1(n536), .A2(n397), .ZN(n398) );
  XOR2_X1 U452 ( .A(KEYINPUT47), .B(n398), .Z(n399) );
  NOR2_X1 U453 ( .A1(n400), .A2(n399), .ZN(n401) );
  XNOR2_X1 U454 ( .A(n401), .B(KEYINPUT48), .ZN(n541) );
  XOR2_X1 U455 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n403) );
  XNOR2_X1 U456 ( .A(KEYINPUT4), .B(KEYINPUT96), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n411) );
  XOR2_X1 U458 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n405) );
  XNOR2_X1 U459 ( .A(KEYINPUT95), .B(KEYINPUT93), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U461 ( .A(n406), .B(KEYINPUT91), .Z(n409) );
  XNOR2_X1 U462 ( .A(G162GAT), .B(n407), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U464 ( .A(n411), .B(n410), .Z(n421) );
  XOR2_X1 U465 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n413) );
  XNOR2_X1 U466 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(n414), .ZN(n442) );
  INV_X1 U469 ( .A(n442), .ZN(n419) );
  XOR2_X1 U470 ( .A(KEYINPUT1), .B(n415), .Z(n417) );
  NAND2_X1 U471 ( .A1(G225GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U474 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U475 ( .A(n423), .B(n422), .ZN(n425) );
  XNOR2_X1 U476 ( .A(n425), .B(n424), .ZN(n458) );
  NOR2_X1 U477 ( .A1(n541), .A2(n563), .ZN(n528) );
  NAND2_X1 U478 ( .A1(n547), .A2(n528), .ZN(n426) );
  NOR2_X1 U479 ( .A1(n459), .A2(n426), .ZN(n427) );
  XNOR2_X1 U480 ( .A(KEYINPUT112), .B(n427), .ZN(n444) );
  XOR2_X1 U481 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n429) );
  XNOR2_X1 U482 ( .A(G218GAT), .B(G106GAT), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U484 ( .A(G148GAT), .B(KEYINPUT22), .Z(n431) );
  XNOR2_X1 U485 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U487 ( .A(n433), .B(n432), .Z(n439) );
  XOR2_X1 U488 ( .A(n434), .B(G78GAT), .Z(n436) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U491 ( .A(G22GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n543) );
  XNOR2_X1 U495 ( .A(KEYINPUT28), .B(n543), .ZN(n512) );
  NAND2_X1 U496 ( .A1(n444), .A2(n512), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n445), .B(KEYINPUT113), .ZN(n521) );
  INV_X1 U498 ( .A(n446), .ZN(n447) );
  NAND2_X1 U499 ( .A1(n521), .A2(n447), .ZN(n450) );
  XOR2_X1 U500 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n448) );
  NOR2_X1 U501 ( .A1(n543), .A2(n547), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n451), .B(KEYINPUT26), .ZN(n565) );
  INV_X1 U503 ( .A(n565), .ZN(n452) );
  NOR2_X1 U504 ( .A1(n452), .A2(n459), .ZN(n527) );
  INV_X1 U505 ( .A(n547), .ZN(n508) );
  OR2_X1 U506 ( .A1(n540), .A2(n508), .ZN(n453) );
  NAND2_X1 U507 ( .A1(n453), .A2(n543), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n454), .B(KEYINPUT99), .ZN(n455) );
  XOR2_X1 U509 ( .A(KEYINPUT25), .B(n455), .Z(n456) );
  NOR2_X1 U510 ( .A1(n527), .A2(n456), .ZN(n457) );
  NOR2_X1 U511 ( .A1(n458), .A2(n457), .ZN(n463) );
  NOR2_X1 U512 ( .A1(n563), .A2(n459), .ZN(n460) );
  NAND2_X1 U513 ( .A1(n512), .A2(n460), .ZN(n461) );
  NOR2_X1 U514 ( .A1(n547), .A2(n461), .ZN(n462) );
  NOR2_X1 U515 ( .A1(n463), .A2(n462), .ZN(n477) );
  INV_X1 U516 ( .A(n574), .ZN(n522) );
  NAND2_X1 U517 ( .A1(n522), .A2(n446), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n464), .B(KEYINPUT16), .ZN(n465) );
  XNOR2_X1 U519 ( .A(n465), .B(KEYINPUT78), .ZN(n466) );
  NOR2_X1 U520 ( .A1(n477), .A2(n466), .ZN(n493) );
  NAND2_X1 U521 ( .A1(n516), .A2(n571), .ZN(n467) );
  XOR2_X1 U522 ( .A(KEYINPUT74), .B(n467), .Z(n481) );
  NAND2_X1 U523 ( .A1(n493), .A2(n481), .ZN(n474) );
  NOR2_X1 U524 ( .A1(n563), .A2(n474), .ZN(n469) );
  XNOR2_X1 U525 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U527 ( .A(G1GAT), .B(n470), .Z(G1324GAT) );
  NOR2_X1 U528 ( .A1(n540), .A2(n474), .ZN(n471) );
  XOR2_X1 U529 ( .A(G8GAT), .B(n471), .Z(G1325GAT) );
  NOR2_X1 U530 ( .A1(n508), .A2(n474), .ZN(n473) );
  XNOR2_X1 U531 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(G1326GAT) );
  NOR2_X1 U533 ( .A1(n512), .A2(n474), .ZN(n475) );
  XOR2_X1 U534 ( .A(G22GAT), .B(n475), .Z(G1327GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT38), .B(KEYINPUT103), .Z(n483) );
  NOR2_X1 U536 ( .A1(n476), .A2(n477), .ZN(n478) );
  NAND2_X1 U537 ( .A1(n574), .A2(n478), .ZN(n479) );
  XNOR2_X1 U538 ( .A(KEYINPUT37), .B(n479), .ZN(n480) );
  XNOR2_X1 U539 ( .A(KEYINPUT102), .B(n480), .ZN(n504) );
  NAND2_X1 U540 ( .A1(n481), .A2(n504), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(n490) );
  NOR2_X1 U542 ( .A1(n490), .A2(n563), .ZN(n486) );
  XOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT101), .Z(n484) );
  XNOR2_X1 U544 ( .A(KEYINPUT39), .B(n484), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  NOR2_X1 U546 ( .A1(n490), .A2(n540), .ZN(n487) );
  XOR2_X1 U547 ( .A(G36GAT), .B(n487), .Z(G1329GAT) );
  NOR2_X1 U548 ( .A1(n490), .A2(n508), .ZN(n488) );
  XOR2_X1 U549 ( .A(KEYINPUT40), .B(n488), .Z(n489) );
  XNOR2_X1 U550 ( .A(G43GAT), .B(n489), .ZN(G1330GAT) );
  NOR2_X1 U551 ( .A1(n512), .A2(n490), .ZN(n491) );
  XOR2_X1 U552 ( .A(G50GAT), .B(n491), .Z(G1331GAT) );
  INV_X1 U553 ( .A(n518), .ZN(n555) );
  NOR2_X1 U554 ( .A1(n516), .A2(n555), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n492), .B(KEYINPUT104), .ZN(n503) );
  NAND2_X1 U556 ( .A1(n493), .A2(n503), .ZN(n499) );
  NOR2_X1 U557 ( .A1(n563), .A2(n499), .ZN(n494) );
  XOR2_X1 U558 ( .A(G57GAT), .B(n494), .Z(n495) );
  XNOR2_X1 U559 ( .A(KEYINPUT42), .B(n495), .ZN(G1332GAT) );
  NOR2_X1 U560 ( .A1(n540), .A2(n499), .ZN(n496) );
  XOR2_X1 U561 ( .A(G64GAT), .B(n496), .Z(G1333GAT) );
  NOR2_X1 U562 ( .A1(n508), .A2(n499), .ZN(n498) );
  XNOR2_X1 U563 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n498), .B(n497), .ZN(G1334GAT) );
  NOR2_X1 U565 ( .A1(n512), .A2(n499), .ZN(n501) );
  XNOR2_X1 U566 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G78GAT), .B(n502), .ZN(G1335GAT) );
  NAND2_X1 U569 ( .A1(n504), .A2(n503), .ZN(n511) );
  NOR2_X1 U570 ( .A1(n563), .A2(n511), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n505), .B(KEYINPUT107), .ZN(n506) );
  XNOR2_X1 U572 ( .A(G85GAT), .B(n506), .ZN(G1336GAT) );
  NOR2_X1 U573 ( .A1(n540), .A2(n511), .ZN(n507) );
  XOR2_X1 U574 ( .A(G92GAT), .B(n507), .Z(G1337GAT) );
  NOR2_X1 U575 ( .A1(n508), .A2(n511), .ZN(n509) );
  XOR2_X1 U576 ( .A(KEYINPUT108), .B(n509), .Z(n510) );
  XNOR2_X1 U577 ( .A(G99GAT), .B(n510), .ZN(G1338GAT) );
  NOR2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n514) );
  XNOR2_X1 U579 ( .A(KEYINPUT109), .B(KEYINPUT44), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G106GAT), .B(n515), .ZN(G1339GAT) );
  NAND2_X1 U582 ( .A1(n516), .A2(n521), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U584 ( .A(G120GAT), .B(KEYINPUT49), .Z(n520) );
  NAND2_X1 U585 ( .A1(n521), .A2(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1341GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n526) );
  XOR2_X1 U588 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n524) );
  XNOR2_X1 U589 ( .A(G127GAT), .B(KEYINPUT114), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(G1342GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n537) );
  NOR2_X1 U593 ( .A1(n567), .A2(n537), .ZN(n529) );
  XOR2_X1 U594 ( .A(G141GAT), .B(n529), .Z(G1344GAT) );
  NOR2_X1 U595 ( .A1(n555), .A2(n537), .ZN(n534) );
  XOR2_X1 U596 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n531) );
  XNOR2_X1 U597 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(KEYINPUT52), .B(n532), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1345GAT) );
  NOR2_X1 U601 ( .A1(n574), .A2(n537), .ZN(n535) );
  XOR2_X1 U602 ( .A(G155GAT), .B(n535), .Z(G1346GAT) );
  INV_X1 U603 ( .A(n536), .ZN(n538) );
  NOR2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U605 ( .A(G162GAT), .B(n539), .Z(G1347GAT) );
  NOR2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(KEYINPUT54), .ZN(n564) );
  AND2_X1 U608 ( .A1(n563), .A2(n543), .ZN(n544) );
  NAND2_X1 U609 ( .A1(n564), .A2(n544), .ZN(n546) );
  XOR2_X1 U610 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n549), .B(KEYINPUT120), .ZN(n554) );
  NOR2_X1 U614 ( .A1(n554), .A2(n567), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(KEYINPUT121), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G169GAT), .B(n551), .ZN(G1348GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n553) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n557) );
  NOR2_X1 U620 ( .A1(n554), .A2(n555), .ZN(n556) );
  XOR2_X1 U621 ( .A(n557), .B(n556), .Z(G1349GAT) );
  NOR2_X1 U622 ( .A1(n574), .A2(n554), .ZN(n558) );
  XOR2_X1 U623 ( .A(G183GAT), .B(n558), .Z(G1350GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n560) );
  XNOR2_X1 U625 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n562) );
  NOR2_X1 U627 ( .A1(n446), .A2(n554), .ZN(n561) );
  XOR2_X1 U628 ( .A(n562), .B(n561), .Z(G1351GAT) );
  AND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n578) );
  NOR2_X1 U631 ( .A1(n567), .A2(n578), .ZN(n570) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n571), .A2(n578), .ZN(n573) );
  XNOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NOR2_X1 U638 ( .A1(n574), .A2(n578), .ZN(n576) );
  XNOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n476), .A2(n578), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

