//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT65), .Z(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT67), .B1(new_n461), .B2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n466), .A2(new_n467), .A3(G137), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(new_n464), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n470), .A2(G137), .A3(new_n468), .A4(new_n462), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n473), .B1(G2104), .B2(new_n468), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NOR3_X1   g050(.A1(new_n475), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n476));
  OR2_X1    g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(G101), .ZN(new_n479));
  OAI21_X1  g054(.A(G101), .B1(new_n474), .B2(new_n476), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT70), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n469), .A2(new_n472), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n464), .A2(new_n483), .A3(G125), .ZN(new_n484));
  NAND2_X1  g059(.A1(G113), .A2(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n468), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G160));
  NAND2_X1  g065(.A1(new_n466), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n466), .A2(new_n468), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G136), .ZN(new_n496));
  NOR2_X1   g071(.A1(G100), .A2(G2105), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT71), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n493), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G162));
  NAND4_X1  g076(.A1(new_n470), .A2(G138), .A3(new_n468), .A4(new_n462), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  AND4_X1   g080(.A1(new_n468), .A2(new_n505), .A3(new_n464), .A4(new_n483), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n470), .A2(G126), .A3(G2105), .A4(new_n462), .ZN(new_n509));
  OR2_X1    g084(.A1(G102), .A2(G2105), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n510), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n508), .A2(KEYINPUT72), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n506), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(new_n512), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(G164));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(new_n523), .B1(new_n520), .B2(G543), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n524), .A2(G62), .ZN(new_n532));
  NAND2_X1  g107(.A1(G75), .A2(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G166));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XOR2_X1   g114(.A(new_n539), .B(KEYINPUT7), .Z(new_n540));
  AND3_X1   g115(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n541));
  INV_X1    g116(.A(new_n528), .ZN(new_n542));
  AOI211_X1 g117(.A(new_n540), .B(new_n541), .C1(G51), .C2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n526), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G89), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(G168));
  AOI22_X1  g122(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n531), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n526), .A2(new_n550), .B1(new_n528), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(G171));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n526), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n531), .ZN(new_n557));
  AOI211_X1 g132(.A(new_n555), .B(new_n557), .C1(G43), .C2(new_n542), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND3_X1  g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT75), .Z(G176));
  XOR2_X1   g138(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n564));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(new_n524), .ZN(new_n569));
  XNOR2_X1  g144(.A(KEYINPUT78), .B(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT79), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n542), .A2(G53), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT9), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n544), .A2(G91), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT77), .Z(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  NAND2_X1  g155(.A1(G168), .A2(KEYINPUT80), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n546), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G286));
  INV_X1    g159(.A(G166), .ZN(G303));
  NAND2_X1  g160(.A1(new_n544), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n542), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n591));
  OR3_X1    g166(.A1(new_n590), .A2(new_n591), .A3(new_n531), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n590), .B2(new_n531), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n592), .A2(new_n593), .B1(G48), .B2(new_n542), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n524), .A2(G86), .A3(new_n525), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT82), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n531), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n526), .A2(new_n600), .B1(new_n528), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n544), .A2(G92), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n542), .A2(G54), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n524), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n531), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n605), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n605), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  XOR2_X1   g189(.A(G299), .B(KEYINPUT83), .Z(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT84), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g199(.A1(new_n464), .A2(new_n483), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n477), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n632), .B(new_n633), .C1(G111), .C2(new_n468), .ZN(new_n634));
  INV_X1    g209(.A(G135), .ZN(new_n635));
  INV_X1    g210(.A(G123), .ZN(new_n636));
  OAI221_X1 g211(.A(new_n634), .B1(new_n494), .B2(new_n635), .C1(new_n636), .C2(new_n491), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n629), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT15), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2435), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT87), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n650), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(new_n651), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n650), .A2(KEYINPUT87), .A3(new_n652), .ZN(new_n658));
  NAND4_X1  g233(.A1(new_n655), .A2(G14), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT88), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n663), .B(KEYINPUT17), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n664), .B1(new_n666), .B2(new_n662), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT90), .Z(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n662), .A3(new_n661), .ZN(new_n669));
  INV_X1    g244(.A(new_n662), .ZN(new_n670));
  INV_X1    g245(.A(new_n663), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n671), .A3(new_n661), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n668), .A2(new_n669), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT91), .Z(new_n676));
  XNOR2_X1  g251(.A(G2096), .B(G2100), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT92), .ZN(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n681), .A2(new_n682), .ZN(new_n688));
  AOI22_X1  g263(.A1(new_n686), .A2(new_n687), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  OR3_X1    g264(.A1(new_n683), .A2(new_n688), .A3(new_n685), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n689), .B(new_n690), .C1(new_n687), .C2(new_n686), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1986), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT93), .B(G1981), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  OAI21_X1  g274(.A(KEYINPUT99), .B1(G16), .B2(G21), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n546), .A2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(new_n700), .B(KEYINPUT99), .S(new_n702), .Z(new_n703));
  INV_X1    g278(.A(G1966), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT100), .Z(new_n706));
  NAND2_X1  g281(.A1(G299), .A2(G16), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n701), .A2(KEYINPUT23), .A3(G20), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT23), .ZN(new_n709));
  INV_X1    g284(.A(G20), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G16), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n707), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1956), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n701), .A2(G4), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n611), .B2(new_n701), .ZN(new_n715));
  INV_X1    g290(.A(G1348), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G27), .A2(G29), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G164), .B2(G29), .ZN(new_n719));
  INV_X1    g294(.A(G2078), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G35), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G162), .B2(new_n723), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G2090), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n701), .A2(G5), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G171), .B2(new_n701), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT101), .B(G1961), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  AND2_X1   g306(.A1(KEYINPUT24), .A2(G34), .ZN(new_n732));
  NOR2_X1   g307(.A1(KEYINPUT24), .A2(G34), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n732), .A2(new_n733), .A3(G29), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n489), .B2(G29), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT95), .Z(new_n736));
  OAI211_X1 g311(.A(new_n727), .B(new_n731), .C1(G2084), .C2(new_n736), .ZN(new_n737));
  NOR4_X1   g312(.A1(new_n706), .A2(new_n713), .A3(new_n722), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n723), .A2(G32), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n492), .A2(G129), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n495), .A2(G141), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n477), .A2(G105), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n740), .A2(new_n741), .A3(new_n742), .A4(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(new_n723), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT97), .Z(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n736), .A2(G2084), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  AOI22_X1  g329(.A1(new_n625), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  INV_X1    g330(.A(G139), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n754), .B1(new_n755), .B2(new_n468), .C1(new_n494), .C2(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G33), .B(new_n757), .S(G29), .Z(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(G2072), .Z(new_n759));
  NAND3_X1  g334(.A1(new_n751), .A2(new_n752), .A3(new_n759), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT98), .Z(new_n761));
  OAI22_X1  g336(.A1(new_n749), .A2(new_n750), .B1(G2090), .B2(new_n726), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n723), .A2(G26), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n492), .A2(G128), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n495), .A2(G140), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n468), .A2(G116), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n764), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n763), .B1(new_n768), .B2(G29), .ZN(new_n769));
  MUX2_X1   g344(.A(new_n763), .B(new_n769), .S(KEYINPUT28), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT30), .B(G28), .Z(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(G29), .B2(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n762), .B(new_n773), .C1(new_n704), .C2(new_n703), .ZN(new_n774));
  AND3_X1   g349(.A1(new_n738), .A2(new_n761), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n701), .A2(G23), .ZN(new_n776));
  INV_X1    g351(.A(G288), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n701), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT33), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1976), .ZN(new_n780));
  NOR2_X1   g355(.A1(G16), .A2(G22), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G166), .B2(G16), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G1971), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n701), .A2(G6), .ZN(new_n784));
  INV_X1    g359(.A(G305), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n701), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT32), .B(G1981), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT94), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n786), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n780), .A2(new_n783), .A3(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n701), .A2(G24), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n603), .B2(new_n701), .ZN(new_n793));
  INV_X1    g368(.A(G1986), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n723), .A2(G25), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n492), .A2(G119), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n495), .A2(G131), .ZN(new_n799));
  OR2_X1    g374(.A1(G95), .A2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(new_n723), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT35), .B(G1991), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n791), .A2(new_n795), .A3(new_n796), .A4(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT36), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT31), .B(G11), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n775), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n701), .A2(G19), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n558), .B2(new_n701), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1341), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n637), .A2(new_n723), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n811), .A2(new_n814), .A3(new_n815), .ZN(G311));
  INV_X1    g391(.A(G311), .ZN(G150));
  AOI22_X1  g392(.A1(new_n544), .A2(G93), .B1(new_n542), .B2(G55), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n524), .A2(G67), .ZN(new_n819));
  NAND2_X1  g394(.A1(G80), .A2(G543), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n818), .B1(new_n531), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  OR2_X1    g399(.A1(new_n558), .A2(new_n822), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n558), .A2(new_n822), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT39), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n611), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n824), .B1(new_n831), .B2(G860), .ZN(G145));
  XOR2_X1   g407(.A(new_n500), .B(KEYINPUT102), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n637), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n489), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n746), .B(new_n757), .Z(new_n836));
  NOR2_X1   g411(.A1(new_n516), .A2(new_n512), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n768), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n492), .A2(G130), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n495), .A2(G142), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n468), .A2(G118), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n627), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n802), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n839), .A2(KEYINPUT103), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n835), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n839), .B(new_n846), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n848), .B1(new_n850), .B2(KEYINPUT103), .ZN(new_n851));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n851), .B(new_n852), .C1(new_n850), .C2(new_n835), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g429(.A(G166), .B(G288), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G290), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n785), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n855), .A2(new_n603), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n855), .A2(new_n603), .ZN(new_n859));
  OAI21_X1  g434(.A(G305), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(KEYINPUT106), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT42), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT41), .ZN(new_n864));
  NAND2_X1  g439(.A1(G299), .A2(new_n611), .ZN(new_n865));
  INV_X1    g440(.A(new_n611), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n576), .A2(new_n866), .A3(new_n578), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT104), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(KEYINPUT104), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n864), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n865), .A2(new_n867), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n621), .B(new_n827), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n877), .B2(new_n873), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n863), .B(new_n879), .ZN(new_n880));
  MUX2_X1   g455(.A(new_n822), .B(new_n880), .S(G868), .Z(G295));
  MUX2_X1   g456(.A(new_n822), .B(new_n880), .S(G868), .Z(G331));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n546), .A2(G171), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G286), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n827), .B(new_n885), .C1(new_n886), .C2(G301), .ZN(new_n887));
  AOI21_X1  g462(.A(G301), .B1(new_n581), .B2(new_n583), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n826), .B(new_n825), .C1(new_n888), .C2(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n871), .B2(new_n875), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n872), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(G37), .B1(new_n894), .B2(new_n861), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n857), .A2(new_n860), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n891), .B2(new_n893), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT44), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n868), .A2(new_n870), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n887), .A2(new_n889), .A3(KEYINPUT41), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n892), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n873), .A2(new_n874), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n897), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n896), .B1(new_n895), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n883), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n906), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n908), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n899), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n896), .B1(new_n895), .B2(new_n898), .ZN(new_n912));
  INV_X1    g487(.A(new_n891), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n861), .A3(new_n892), .ZN(new_n914));
  AND4_X1   g489(.A1(new_n896), .A2(new_n914), .A3(new_n905), .A4(new_n852), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n911), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n910), .A2(new_n916), .ZN(G397));
  XOR2_X1   g492(.A(new_n768), .B(G2067), .Z(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G1384), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n516), .B2(new_n512), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n922));
  XOR2_X1   g497(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n924), .B(new_n920), .C1(new_n516), .C2(new_n512), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n469), .A2(new_n472), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n479), .A2(new_n481), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n488), .A2(new_n928), .A3(G40), .A4(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n919), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT112), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(G1996), .A3(new_n746), .ZN(new_n936));
  OR3_X1    g511(.A1(new_n932), .A2(KEYINPUT110), .A3(G1996), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT110), .B1(new_n932), .B2(G1996), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n939), .A2(KEYINPUT111), .A3(new_n747), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT111), .B1(new_n939), .B2(new_n747), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n935), .B(new_n936), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n802), .B(new_n806), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n942), .B1(new_n933), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n603), .B(new_n794), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n933), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT54), .ZN(new_n949));
  OAI211_X1 g524(.A(KEYINPUT45), .B(new_n920), .C1(new_n516), .C2(new_n512), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT53), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(G2078), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n950), .A2(new_n482), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G40), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n484), .A2(new_n485), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT121), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n956), .B2(G2105), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n926), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n926), .A2(new_n953), .A3(KEYINPUT122), .A4(new_n957), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n514), .A2(new_n920), .A3(new_n517), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n923), .ZN(new_n963));
  INV_X1    g538(.A(new_n950), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(new_n930), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(new_n965), .A3(new_n720), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n960), .A2(new_n961), .B1(new_n951), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n930), .B1(new_n962), .B2(KEYINPUT50), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n969), .B(new_n920), .C1(new_n516), .C2(new_n512), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT114), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1961), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT120), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT120), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n975), .B(G1961), .C1(new_n968), .C2(new_n971), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n967), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n949), .B1(new_n977), .B2(G171), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n972), .A2(new_n973), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n966), .A2(new_n951), .ZN(new_n980));
  INV_X1    g555(.A(new_n921), .ZN(new_n981));
  OAI221_X1 g556(.A(new_n931), .B1(KEYINPUT45), .B2(new_n981), .C1(new_n962), .C2(new_n923), .ZN(new_n982));
  INV_X1    g557(.A(new_n952), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n979), .B(new_n980), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n984), .A2(G171), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n978), .A2(KEYINPUT124), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT124), .B1(new_n978), .B2(new_n985), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n967), .B(G301), .C1(new_n974), .C2(new_n976), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(G171), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n949), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT123), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(KEYINPUT123), .A3(new_n949), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n997));
  INV_X1    g572(.A(G2084), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n968), .A2(new_n971), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n982), .A2(new_n704), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n968), .A2(new_n971), .A3(KEYINPUT116), .A4(new_n998), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n997), .B1(new_n1004), .B2(new_n546), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1001), .A2(G168), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n997), .B1(new_n1006), .B2(G8), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT119), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(KEYINPUT51), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT119), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1011), .B(new_n1012), .C1(new_n1007), .C2(new_n1005), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n536), .A2(G8), .A3(new_n537), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n963), .A2(new_n965), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT113), .B(G1971), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n921), .A2(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n931), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1024), .B2(G2090), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1017), .B1(new_n1025), .B2(G8), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  INV_X1    g602(.A(G1981), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n594), .A2(new_n1028), .A3(new_n596), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n595), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1028), .B1(new_n594), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1027), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n594), .A2(new_n1031), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT49), .B(new_n1029), .C1(new_n1034), .C2(new_n1028), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n931), .A2(new_n981), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n777), .A2(G1976), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(new_n1039), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1038), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1021), .B1(G2090), .B2(new_n972), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G8), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1017), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT115), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1046), .A2(new_n1017), .A3(new_n1050), .A4(G8), .ZN(new_n1051));
  AOI211_X1 g626(.A(new_n1026), .B(new_n1045), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n988), .A2(new_n996), .A3(new_n1014), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT125), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1036), .A2(G2067), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n716), .B2(new_n972), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(new_n866), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT118), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT57), .B1(new_n575), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(G299), .B(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1956), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1018), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT56), .B(G2072), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1024), .A2(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT61), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1067), .B(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT58), .B(G1341), .Z(new_n1071));
  NAND2_X1  g646(.A1(new_n1036), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1018), .B2(G1996), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n558), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1074), .B(KEYINPUT59), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1057), .A2(new_n1076), .A3(new_n611), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1070), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1057), .A2(new_n866), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1076), .B1(new_n1058), .B2(new_n1079), .ZN(new_n1080));
  OAI221_X1 g655(.A(new_n1068), .B1(new_n1062), .B2(new_n1066), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n978), .A2(new_n985), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n978), .A2(KEYINPUT124), .A3(new_n985), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1084), .A2(new_n1052), .A3(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1086), .A2(KEYINPUT125), .A3(new_n1014), .A4(new_n996), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1055), .A2(new_n1081), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1045), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1038), .A2(new_n1042), .A3(new_n777), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1029), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1090), .A2(new_n1091), .B1(new_n1037), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1004), .A2(G8), .A3(new_n886), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT63), .B1(new_n1052), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT63), .ZN(new_n1099));
  NOR4_X1   g674(.A1(new_n1090), .A2(new_n1045), .A3(new_n1095), .A4(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1014), .A2(KEYINPUT62), .ZN(new_n1101));
  INV_X1    g676(.A(new_n990), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1052), .B1(new_n1014), .B2(KEYINPUT62), .ZN(new_n1104));
  OAI221_X1 g679(.A(new_n1094), .B1(new_n1097), .B2(new_n1100), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n948), .B1(new_n1088), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n803), .A2(new_n806), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n942), .A2(new_n1107), .B1(G2067), .B2(new_n768), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1108), .A2(KEYINPUT126), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(KEYINPUT126), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n933), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n933), .B1(new_n919), .B2(new_n746), .ZN(new_n1112));
  INV_X1    g687(.A(new_n939), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1113), .A2(KEYINPUT46), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(KEYINPUT46), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT47), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n933), .A2(new_n794), .A3(new_n603), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT48), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n945), .A2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1111), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1106), .A2(new_n1121), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g697(.A(KEYINPUT127), .ZN(new_n1124));
  AND2_X1   g698(.A1(new_n659), .A2(new_n698), .ZN(new_n1125));
  OAI211_X1 g699(.A(new_n1125), .B(new_n678), .C1(new_n912), .C2(new_n915), .ZN(new_n1126));
  NAND2_X1  g700(.A1(new_n853), .A2(G319), .ZN(new_n1127));
  OAI21_X1  g701(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g702(.A1(new_n659), .A2(new_n698), .ZN(new_n1129));
  NAND3_X1  g703(.A1(new_n914), .A2(new_n898), .A3(new_n852), .ZN(new_n1130));
  NAND2_X1  g704(.A1(new_n1130), .A2(KEYINPUT43), .ZN(new_n1131));
  NAND3_X1  g705(.A1(new_n895), .A2(new_n896), .A3(new_n905), .ZN(new_n1132));
  AOI21_X1  g706(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g707(.A(new_n1127), .ZN(new_n1134));
  NAND4_X1  g708(.A1(new_n1133), .A2(new_n1134), .A3(KEYINPUT127), .A4(new_n678), .ZN(new_n1135));
  NAND2_X1  g709(.A1(new_n1128), .A2(new_n1135), .ZN(G308));
  NAND3_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n678), .ZN(G225));
endmodule


