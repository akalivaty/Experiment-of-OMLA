//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997;
  XOR2_X1   g000(.A(KEYINPUT93), .B(G29gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT94), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n202), .A2(KEYINPUT94), .A3(G36gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT92), .ZN(new_n208));
  OR3_X1    g007(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n207), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT92), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n205), .B(new_n206), .C1(new_n208), .C2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G43gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G50gat), .ZN(new_n215));
  INV_X1    g014(.A(G50gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G43gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT15), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n218), .B(KEYINPUT95), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(new_n206), .A3(new_n205), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT98), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n210), .B1(new_n209), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(new_n223), .B2(new_n209), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n217), .A2(KEYINPUT96), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT97), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n215), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n217), .A2(KEYINPUT96), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT97), .B1(new_n214), .B2(G50gat), .ZN(new_n230));
  NOR4_X1   g029(.A1(new_n226), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n225), .B1(new_n231), .B2(KEYINPUT15), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n220), .B1(new_n222), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT99), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G15gat), .B(G22gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(G1gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n238), .B2(G1gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  AOI211_X1 g039(.A(G8gat), .B(new_n237), .C1(new_n240), .C2(KEYINPUT101), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(KEYINPUT101), .B2(new_n240), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n236), .A2(G1gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT100), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n244), .A3(new_n239), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n245), .B(G8gat), .C1(new_n244), .C2(new_n239), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n220), .B(KEYINPUT99), .C1(new_n222), .C2(new_n232), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n235), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT17), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n251), .A3(new_n248), .ZN(new_n252));
  INV_X1    g051(.A(new_n247), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n233), .A2(new_n251), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G229gat), .A2(G233gat), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT102), .Z(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n250), .A2(new_n255), .A3(KEYINPUT18), .A4(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n257), .B(KEYINPUT13), .Z(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n247), .B1(new_n235), .B2(new_n248), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n249), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(G113gat), .B(G141gat), .Z(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT91), .B(G197gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT11), .B(G169gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT12), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n259), .A2(new_n263), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n250), .A2(new_n255), .A3(new_n258), .ZN(new_n271));
  XOR2_X1   g070(.A(KEYINPUT103), .B(KEYINPUT18), .Z(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT104), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(KEYINPUT104), .A3(new_n272), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n270), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n273), .A2(new_n263), .A3(new_n259), .ZN(new_n278));
  INV_X1    g077(.A(new_n269), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT83), .ZN(new_n283));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT75), .B(G211gat), .ZN(new_n285));
  INV_X1    g084(.A(G218gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n284), .B1(new_n287), .B2(KEYINPUT22), .ZN(new_n288));
  XNOR2_X1  g087(.A(G211gat), .B(G218gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(KEYINPUT76), .B(KEYINPUT29), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G183gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT27), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT27), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G183gat), .ZN(new_n296));
  INV_X1    g095(.A(G190gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(KEYINPUT28), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT27), .B(G183gat), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n299), .A2(KEYINPUT28), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n297), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OR3_X1    g107(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n308), .A2(new_n309), .B1(G183gat), .B2(G190gat), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n305), .A2(KEYINPUT68), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT68), .B1(new_n305), .B2(new_n310), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT24), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(G183gat), .A3(G190gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(G183gat), .B(G190gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(new_n315), .ZN(new_n318));
  INV_X1    g117(.A(G169gat), .ZN(new_n319));
  INV_X1    g118(.A(G176gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT23), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(G169gat), .B2(G176gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n323), .A3(new_n307), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n314), .B1(new_n318), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT65), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT65), .B(new_n314), .C1(new_n318), .C2(new_n324), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n315), .A2(G183gat), .A3(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n293), .A2(G190gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n297), .A2(G183gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n329), .B1(new_n332), .B2(KEYINPUT24), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n307), .A2(KEYINPUT66), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(new_n314), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n307), .A2(KEYINPUT66), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n321), .A2(new_n336), .A3(new_n323), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n327), .A2(new_n328), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n292), .B1(new_n313), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G226gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n305), .A2(new_n310), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n345));
  OAI22_X1  g144(.A1(new_n340), .A2(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n344), .A2(new_n345), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n290), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n339), .A2(new_n343), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n342), .A2(KEYINPUT29), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n313), .A2(new_n339), .A3(new_n342), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n288), .B(new_n289), .Z(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n313), .A2(new_n342), .A3(new_n339), .ZN(new_n357));
  INV_X1    g156(.A(new_n350), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n358), .B1(new_n339), .B2(new_n343), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n355), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT78), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n348), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT79), .ZN(new_n363));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n348), .A2(new_n368), .A3(new_n361), .A4(new_n356), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n363), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n348), .A2(new_n366), .A3(new_n361), .A4(new_n356), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT30), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n354), .B1(new_n353), .B2(new_n355), .ZN(new_n373));
  AOI211_X1 g172(.A(KEYINPUT78), .B(new_n290), .C1(new_n351), .C2(new_n352), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n366), .A4(new_n348), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n382));
  AND2_X1   g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(G141gat), .A2(G148gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G141gat), .ZN(new_n386));
  INV_X1    g185(.A(G148gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(KEYINPUT81), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391));
  OR3_X1    g190(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n385), .A2(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G155gat), .ZN(new_n394));
  INV_X1    g193(.A(G162gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n391), .ZN(new_n397));
  XOR2_X1   g196(.A(KEYINPUT80), .B(KEYINPUT2), .Z(new_n398));
  NOR2_X1   g197(.A1(new_n383), .A2(new_n384), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(new_n393), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n388), .A2(new_n389), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT80), .B(KEYINPUT2), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n391), .B(new_n396), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n385), .A2(new_n390), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n392), .A2(new_n391), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n402), .B(new_n405), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n401), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(G113gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n410), .A2(G120gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(G120gat), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(KEYINPUT71), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(KEYINPUT71), .B2(new_n412), .ZN(new_n414));
  INV_X1    g213(.A(G134gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G127gat), .ZN(new_n416));
  INV_X1    g215(.A(G127gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G134gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(KEYINPUT1), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT70), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT69), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G127gat), .B(G134gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT69), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT1), .ZN(new_n428));
  INV_X1    g227(.A(G120gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(G113gat), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n411), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n422), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n416), .A2(new_n418), .A3(KEYINPUT69), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT69), .B1(new_n416), .B2(new_n418), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n422), .B(new_n431), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n421), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n381), .B1(new_n409), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT70), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n435), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n393), .A2(new_n400), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n421), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n440), .A2(new_n435), .B1(new_n414), .B2(new_n420), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n446), .A2(KEYINPUT4), .A3(new_n442), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n438), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n443), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n446), .A2(new_n442), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n381), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(new_n451), .A3(KEYINPUT5), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453));
  XNOR2_X1  g252(.A(G1gat), .B(G29gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT0), .ZN(new_n455));
  XNOR2_X1  g254(.A(G57gat), .B(G85gat), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n455), .B(new_n456), .Z(new_n457));
  INV_X1    g256(.A(KEYINPUT5), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n438), .A2(new_n445), .A3(new_n458), .A4(new_n447), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n452), .A2(new_n453), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n452), .A2(new_n459), .ZN(new_n463));
  INV_X1    g262(.A(new_n457), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n457), .B1(new_n452), .B2(new_n459), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n457), .A3(new_n459), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(KEYINPUT82), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n466), .B1(new_n469), .B2(KEYINPUT6), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n283), .B1(new_n379), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n472));
  NAND2_X1  g271(.A1(G228gat), .A2(G233gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n355), .A2(new_n291), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n442), .B1(new_n474), .B2(new_n402), .ZN(new_n475));
  INV_X1    g274(.A(new_n408), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n290), .B1(new_n476), .B2(new_n292), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n473), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n442), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n290), .A2(KEYINPUT29), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(KEYINPUT3), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n482), .A2(G228gat), .A3(G233gat), .A4(new_n477), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n472), .B1(new_n484), .B2(G22gat), .ZN(new_n485));
  INV_X1    g284(.A(G22gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n479), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  XNOR2_X1  g286(.A(G78gat), .B(G106gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(new_n216), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT85), .ZN(new_n490));
  XOR2_X1   g289(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n484), .A2(new_n472), .A3(G22gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n290), .A2(new_n292), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n480), .B1(new_n496), .B2(KEYINPUT3), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n497), .A2(new_n477), .B1(G228gat), .B2(G233gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT29), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n355), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n442), .B1(new_n500), .B2(new_n402), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n477), .A2(G228gat), .A3(G233gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(KEYINPUT86), .B(G22gat), .C1(new_n498), .C2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n492), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(G22gat), .B1(new_n498), .B2(new_n503), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n487), .A3(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n494), .A2(new_n495), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n468), .A2(KEYINPUT82), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT6), .B1(new_n511), .B2(new_n465), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n467), .B1(new_n461), .B2(new_n460), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n514), .A2(KEYINPUT83), .A3(new_n370), .A4(new_n378), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n471), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n321), .A2(new_n323), .A3(new_n307), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT25), .B1(new_n333), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n338), .B1(new_n518), .B2(KEYINPUT65), .ZN(new_n519));
  INV_X1    g318(.A(new_n328), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n343), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n305), .A2(KEYINPUT68), .A3(new_n310), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n446), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n313), .A2(new_n339), .A3(new_n437), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G227gat), .A2(G233gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT64), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n532), .A2(KEYINPUT34), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(KEYINPUT34), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n526), .A2(new_n530), .A3(new_n527), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT32), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT33), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G15gat), .B(G43gat), .Z(new_n540));
  XNOR2_X1  g339(.A(G71gat), .B(G99gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n542), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n536), .B(KEYINPUT32), .C1(new_n538), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n535), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n533), .A2(new_n543), .A3(new_n534), .A4(new_n545), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(KEYINPUT74), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT74), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(KEYINPUT36), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT72), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n543), .A2(new_n554), .A3(new_n545), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n554), .B1(new_n543), .B2(new_n545), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n535), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT73), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT73), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n559), .B(new_n535), .C1(new_n555), .C2(new_n556), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n560), .A3(new_n548), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n553), .B1(new_n561), .B2(KEYINPUT36), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n355), .B1(new_n346), .B2(new_n347), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT37), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n564), .B1(new_n353), .B2(new_n290), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT38), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n348), .A2(new_n564), .A3(new_n361), .A4(new_n356), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n567), .A3(new_n367), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n568), .B(new_n371), .C1(new_n512), .C2(new_n513), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT89), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n470), .A2(KEYINPUT89), .A3(new_n568), .A4(new_n371), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n363), .A2(KEYINPUT37), .A3(new_n369), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n567), .A2(new_n367), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT38), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n437), .A2(new_n480), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(new_n443), .A3(new_n380), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT88), .Z(new_n580));
  AND2_X1   g379(.A1(new_n445), .A2(new_n447), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n409), .A2(new_n437), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n380), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n584), .A3(KEYINPUT39), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT39), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n464), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n585), .A2(new_n587), .A3(KEYINPUT40), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT40), .B1(new_n585), .B2(new_n587), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n588), .A2(new_n589), .A3(new_n467), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n510), .B1(new_n590), .B2(new_n379), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n577), .A2(new_n591), .A3(KEYINPUT90), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT90), .B1(new_n577), .B2(new_n591), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n516), .B(new_n562), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n509), .A2(new_n505), .A3(new_n504), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n507), .A2(KEYINPUT87), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n596), .A2(new_n495), .A3(new_n487), .A4(new_n492), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n600), .A2(new_n470), .A3(new_n379), .ZN(new_n601));
  INV_X1    g400(.A(new_n552), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n558), .A2(new_n598), .A3(new_n560), .A4(new_n548), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n471), .B2(new_n515), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n605), .B2(new_n599), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n282), .B1(new_n594), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G57gat), .B(G64gat), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G71gat), .B(G78gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT105), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(new_n417), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n247), .B1(new_n614), .B2(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n617), .B(G127gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n619), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(new_n394), .ZN(new_n626));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n620), .A2(new_n623), .A3(new_n628), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(KEYINPUT41), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n235), .A2(new_n248), .ZN(new_n638));
  NAND2_X1  g437(.A1(G85gat), .A2(G92gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT7), .ZN(new_n640));
  NAND2_X1  g439(.A1(G99gat), .A2(G106gat), .ZN(new_n641));
  INV_X1    g440(.A(G85gat), .ZN(new_n642));
  INV_X1    g441(.A(G92gat), .ZN(new_n643));
  AOI22_X1  g442(.A1(KEYINPUT8), .A2(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G99gat), .B(G106gat), .Z(new_n646));
  OR2_X1    g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n638), .A2(new_n649), .B1(KEYINPUT41), .B2(new_n633), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n651));
  INV_X1    g450(.A(new_n649), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n252), .A2(new_n254), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT107), .B(G190gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n286), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n651), .B1(new_n650), .B2(new_n653), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n656), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n650), .A2(new_n651), .A3(new_n653), .A4(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n637), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n665), .B(new_n636), .C1(new_n658), .C2(new_n657), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(G230gat), .A2(G233gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT10), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n648), .A2(KEYINPUT109), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n648), .A2(KEYINPUT109), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n671), .A2(new_n612), .A3(new_n647), .A4(new_n672), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n670), .B(new_n673), .C1(new_n614), .C2(new_n649), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n614), .A2(KEYINPUT10), .A3(new_n649), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n669), .B1(new_n676), .B2(KEYINPUT110), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n674), .A2(new_n678), .A3(new_n675), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n673), .B1(new_n614), .B2(new_n649), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n669), .ZN(new_n682));
  XNOR2_X1  g481(.A(G120gat), .B(G148gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(G176gat), .B(G204gat), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n683), .B(new_n684), .Z(new_n685));
  NAND3_X1  g484(.A1(new_n680), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n669), .B1(new_n674), .B2(new_n675), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n682), .ZN(new_n689));
  INV_X1    g488(.A(new_n685), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n632), .A2(new_n667), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n607), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n514), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(G1gat), .Z(G1324gat));
  INV_X1    g497(.A(KEYINPUT111), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n607), .A2(new_n379), .A3(new_n695), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT16), .B(G8gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n702), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n700), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(KEYINPUT42), .B2(new_n702), .ZN(G1325gat));
  XOR2_X1   g503(.A(new_n562), .B(KEYINPUT112), .Z(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G15gat), .B1(new_n696), .B2(new_n706), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n552), .A2(G15gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n696), .B2(new_n708), .ZN(G1326gat));
  NOR2_X1   g508(.A1(new_n696), .A2(new_n598), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT43), .B(G22gat), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n594), .A2(new_n606), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n664), .A2(new_n666), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n713), .ZN(new_n717));
  AND4_X1   g516(.A1(new_n598), .A2(new_n558), .A3(new_n560), .A4(new_n548), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n471), .A2(new_n515), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n599), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR4_X1   g519(.A1(new_n600), .A2(new_n552), .A3(new_n470), .A4(new_n379), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT113), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT113), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n603), .B(new_n723), .C1(new_n605), .C2(new_n599), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n717), .B1(new_n725), .B2(new_n594), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n716), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n632), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n693), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n282), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT114), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n593), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n577), .A2(new_n591), .A3(KEYINPUT90), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n562), .A2(new_n516), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n735), .A2(new_n736), .B1(new_n722), .B2(new_n724), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n667), .B1(new_n594), .B2(new_n606), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n737), .A2(new_n717), .B1(new_n738), .B2(new_n713), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(new_n740), .A3(new_n730), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n732), .A2(new_n470), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n202), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n738), .A2(new_n730), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n744), .A2(new_n514), .A3(new_n202), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT45), .Z(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(G1328gat));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n379), .A3(new_n741), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G36gat), .ZN(new_n749));
  INV_X1    g548(.A(new_n379), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n744), .A2(G36gat), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT46), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(G1329gat));
  NAND2_X1  g552(.A1(new_n739), .A2(new_n730), .ZN(new_n754));
  OAI21_X1  g553(.A(G43gat), .B1(new_n754), .B2(new_n562), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n552), .A2(G43gat), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n744), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n738), .A2(KEYINPUT115), .A3(new_n730), .A4(new_n757), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n761), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n732), .A2(new_n705), .A3(new_n741), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(G43gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n765), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g565(.A(G50gat), .B1(new_n754), .B2(new_n598), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n729), .A2(G50gat), .A3(new_n598), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n607), .A2(new_n715), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(KEYINPUT48), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n769), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n732), .A2(new_n510), .A3(new_n741), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(G50gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n773), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g573(.A1(new_n725), .A2(new_n594), .ZN(new_n775));
  NOR4_X1   g574(.A1(new_n728), .A2(new_n281), .A3(new_n715), .A4(new_n693), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n470), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g579(.A1(new_n777), .A2(new_n750), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  AND2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(G1333gat));
  NOR3_X1   g584(.A1(new_n777), .A2(G71gat), .A3(new_n552), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n778), .A2(new_n705), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(G71gat), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g588(.A1(new_n778), .A2(new_n510), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g590(.A1(new_n728), .A2(new_n282), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n667), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(new_n642), .A3(new_n470), .A4(new_n692), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n792), .A2(new_n693), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n739), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n470), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n797), .B1(new_n801), .B2(new_n642), .ZN(G1336gat));
  AOI21_X1  g601(.A(new_n643), .B1(new_n799), .B2(new_n379), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n750), .A2(new_n693), .A3(G92gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n796), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n804), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n794), .B(KEYINPUT51), .ZN(new_n809));
  INV_X1    g608(.A(new_n806), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT52), .B1(new_n811), .B2(new_n803), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n812), .ZN(G1337gat));
  OAI211_X1 g612(.A(new_n705), .B(new_n798), .C1(new_n716), .C2(new_n726), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n739), .A2(KEYINPUT116), .A3(new_n705), .A4(new_n798), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(G99gat), .A3(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n552), .A2(G99gat), .A3(new_n693), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n796), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT117), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1338gat));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n598), .A2(new_n693), .A3(G106gat), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n809), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n739), .A2(new_n510), .A3(new_n798), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G106gat), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT53), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT118), .B1(new_n796), .B2(new_n827), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n831), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(G1339gat));
  AND3_X1   g636(.A1(new_n270), .A2(new_n275), .A3(new_n276), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n250), .A2(new_n255), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n257), .ZN(new_n840));
  OR3_X1    g639(.A1(new_n249), .A2(new_n262), .A3(new_n261), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(new_n268), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n838), .A2(new_n693), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT54), .B1(new_n676), .B2(new_n668), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n846), .B1(new_n677), .B2(new_n679), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n685), .B1(new_n687), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n845), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n676), .A2(KEYINPUT110), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n852), .A2(new_n668), .A3(new_n679), .ZN(new_n853));
  OAI211_X1 g652(.A(KEYINPUT55), .B(new_n849), .C1(new_n853), .C2(new_n846), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n851), .A2(new_n854), .A3(new_n686), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n280), .B2(new_n277), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n667), .B1(new_n844), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT119), .B1(new_n838), .B2(new_n843), .ZN(new_n858));
  INV_X1    g657(.A(new_n843), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n277), .ZN(new_n861));
  INV_X1    g660(.A(new_n855), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n858), .A2(new_n715), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n728), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n695), .A2(new_n282), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n632), .B1(new_n857), .B2(new_n863), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n694), .A2(new_n281), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT120), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n510), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n379), .A2(new_n514), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n602), .A3(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(new_n410), .A3(new_n282), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n604), .B1(new_n868), .B2(new_n871), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n281), .A3(new_n873), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n410), .B2(new_n877), .ZN(G1340gat));
  NOR3_X1   g677(.A1(new_n874), .A2(new_n429), .A3(new_n693), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n876), .A2(new_n692), .A3(new_n873), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n429), .B2(new_n880), .ZN(G1341gat));
  OAI21_X1  g680(.A(G127gat), .B1(new_n874), .B2(new_n728), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n876), .A2(new_n873), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n632), .A2(new_n417), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT121), .ZN(G1342gat));
  NAND4_X1  g685(.A1(new_n876), .A2(new_n415), .A3(new_n715), .A4(new_n873), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n887), .A2(KEYINPUT56), .ZN(new_n888));
  OAI21_X1  g687(.A(G134gat), .B1(new_n874), .B2(new_n667), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(KEYINPUT56), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(G1343gat));
  NAND2_X1  g690(.A1(new_n562), .A2(new_n873), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n867), .B1(new_n865), .B2(new_n866), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT120), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n510), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n598), .A2(new_n896), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n869), .B2(new_n870), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n892), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n386), .B1(new_n900), .B2(new_n281), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n705), .A2(new_n514), .A3(new_n379), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n598), .B1(new_n868), .B2(new_n871), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(G141gat), .A3(new_n282), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT58), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n892), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n903), .A2(KEYINPUT57), .ZN(new_n908));
  INV_X1    g707(.A(new_n899), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G141gat), .B1(new_n910), .B2(new_n282), .ZN(new_n911));
  INV_X1    g710(.A(new_n905), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n906), .A2(new_n914), .ZN(G1344gat));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n632), .B1(new_n864), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n857), .A2(new_n863), .A3(KEYINPUT122), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n870), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n896), .B1(new_n919), .B2(new_n598), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n868), .A2(new_n871), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n898), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n692), .ZN(new_n924));
  OAI211_X1 g723(.A(KEYINPUT59), .B(G148gat), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT59), .B1(new_n904), .B2(new_n693), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n387), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n693), .A2(KEYINPUT59), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n925), .B(new_n927), .C1(new_n910), .C2(new_n928), .ZN(G1345gat));
  OAI21_X1  g728(.A(G155gat), .B1(new_n910), .B2(new_n728), .ZN(new_n930));
  INV_X1    g729(.A(new_n904), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n394), .A3(new_n632), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1346gat));
  NAND3_X1  g732(.A1(new_n931), .A2(new_n395), .A3(new_n715), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT123), .B1(new_n910), .B2(new_n667), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G162gat), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n910), .A2(KEYINPUT123), .A3(new_n667), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n750), .A2(new_n470), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n602), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n921), .A2(new_n598), .A3(new_n941), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n942), .A2(new_n319), .A3(new_n282), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n876), .A2(new_n939), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n281), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n943), .B1(new_n946), .B2(new_n319), .ZN(G1348gat));
  OAI21_X1  g746(.A(G176gat), .B1(new_n942), .B2(new_n693), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n692), .A2(new_n320), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n944), .B2(new_n949), .ZN(G1349gat));
  NAND3_X1  g749(.A1(new_n945), .A2(new_n302), .A3(new_n632), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT124), .B1(new_n942), .B2(new_n728), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G183gat), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n942), .A2(KEYINPUT124), .A3(new_n728), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT60), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n957), .B(new_n951), .C1(new_n953), .C2(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1350gat));
  NAND3_X1  g758(.A1(new_n872), .A2(new_n715), .A3(new_n941), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n960), .A2(new_n961), .A3(G190gat), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n960), .B2(G190gat), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n715), .A2(new_n297), .ZN(new_n964));
  OAI22_X1  g763(.A1(new_n962), .A2(new_n963), .B1(new_n944), .B2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI221_X1 g766(.A(KEYINPUT125), .B1(new_n944), .B2(new_n964), .C1(new_n962), .C2(new_n963), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1351gat));
  NAND3_X1  g768(.A1(new_n903), .A2(new_n706), .A3(new_n939), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n281), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n706), .A2(new_n939), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n973), .B1(new_n920), .B2(new_n922), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n281), .A2(G197gat), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1352gat));
  NOR3_X1   g775(.A1(new_n970), .A2(G204gat), .A3(new_n693), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT62), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n974), .A2(new_n692), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(G204gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1353gat));
  NAND3_X1  g780(.A1(new_n971), .A2(new_n285), .A3(new_n632), .ZN(new_n982));
  NAND2_X1  g781(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n983));
  INV_X1    g782(.A(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n984), .B1(new_n974), .B2(new_n632), .ZN(new_n985));
  NOR2_X1   g784(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n983), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g787(.A(new_n984), .B(new_n986), .C1(new_n974), .C2(new_n632), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(G1354gat));
  NOR3_X1   g789(.A1(new_n970), .A2(G218gat), .A3(new_n667), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n974), .A2(new_n715), .ZN(new_n994));
  OAI211_X1 g793(.A(new_n992), .B(new_n993), .C1(new_n994), .C2(new_n286), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n286), .B1(new_n974), .B2(new_n715), .ZN(new_n996));
  OAI21_X1  g795(.A(KEYINPUT127), .B1(new_n996), .B2(new_n991), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n995), .A2(new_n997), .ZN(G1355gat));
endmodule


