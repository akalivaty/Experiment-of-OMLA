

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776;

  INV_X1 U376 ( .A(n510), .ZN(n713) );
  XOR2_X1 U377 ( .A(G116), .B(G107), .Z(n535) );
  INV_X1 U378 ( .A(G953), .ZN(n764) );
  XOR2_X1 U379 ( .A(G119), .B(KEYINPUT3), .Z(n355) );
  NOR2_X2 U380 ( .A1(n648), .A2(n647), .ZN(n649) );
  AND2_X4 U381 ( .A1(n441), .A2(n363), .ZN(n739) );
  AND2_X2 U382 ( .A1(n425), .A2(n422), .ZN(n362) );
  INV_X4 U383 ( .A(G143), .ZN(n443) );
  NOR2_X1 U384 ( .A1(G953), .A2(n689), .ZN(n693) );
  XNOR2_X1 U385 ( .A(n719), .B(KEYINPUT81), .ZN(n620) );
  NOR2_X2 U386 ( .A1(n775), .A2(n776), .ZN(n500) );
  NAND2_X1 U387 ( .A1(n619), .A2(n627), .ZN(n719) );
  NAND2_X1 U388 ( .A1(n507), .A2(n504), .ZN(n619) );
  XNOR2_X1 U389 ( .A(n603), .B(KEYINPUT42), .ZN(n776) );
  INV_X1 U390 ( .A(n708), .ZN(n499) );
  AND2_X1 U391 ( .A1(n502), .A2(n501), .ZN(n507) );
  NOR2_X1 U392 ( .A1(n657), .A2(n709), .ZN(n624) );
  AND2_X1 U393 ( .A1(n430), .A2(n622), .ZN(n603) );
  XNOR2_X1 U394 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U395 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U396 ( .A1(n498), .A2(n620), .ZN(n427) );
  NOR2_X2 U397 ( .A1(n578), .A2(n420), .ZN(n419) );
  XNOR2_X1 U398 ( .A(n575), .B(n451), .ZN(n614) );
  XNOR2_X2 U399 ( .A(n562), .B(n561), .ZN(n396) );
  XNOR2_X1 U400 ( .A(n760), .B(G101), .ZN(n562) );
  NAND2_X1 U401 ( .A1(n358), .A2(n458), .ZN(n397) );
  XNOR2_X1 U402 ( .A(n470), .B(G125), .ZN(n538) );
  INV_X1 U403 ( .A(G146), .ZN(n470) );
  XNOR2_X1 U404 ( .A(n405), .B(G137), .ZN(n560) );
  INV_X1 U405 ( .A(G140), .ZN(n405) );
  XNOR2_X1 U406 ( .A(n616), .B(KEYINPUT103), .ZN(n509) );
  NAND2_X1 U407 ( .A1(n614), .A2(n615), .ZN(n616) );
  XNOR2_X1 U408 ( .A(n403), .B(n580), .ZN(n682) );
  XNOR2_X1 U409 ( .A(n400), .B(n399), .ZN(n599) );
  INV_X1 U410 ( .A(G469), .ZN(n399) );
  OR2_X1 U411 ( .A1(n732), .A2(G902), .ZN(n400) );
  XNOR2_X1 U412 ( .A(n432), .B(n431), .ZN(n521) );
  INV_X1 U413 ( .A(KEYINPUT8), .ZN(n431) );
  NAND2_X1 U414 ( .A1(n764), .A2(G234), .ZN(n432) );
  XNOR2_X1 U415 ( .A(n538), .B(n496), .ZN(n762) );
  XNOR2_X1 U416 ( .A(KEYINPUT10), .B(KEYINPUT65), .ZN(n496) );
  INV_X1 U417 ( .A(G478), .ZN(n446) );
  NOR2_X1 U418 ( .A1(G902), .A2(n640), .ZN(n546) );
  XNOR2_X1 U419 ( .A(n513), .B(n511), .ZN(n586) );
  XNOR2_X1 U420 ( .A(n554), .B(n512), .ZN(n511) );
  OR2_X1 U421 ( .A1(n735), .A2(G902), .ZN(n513) );
  INV_X1 U422 ( .A(G475), .ZN(n512) );
  INV_X1 U423 ( .A(KEYINPUT0), .ZN(n440) );
  NAND2_X1 U424 ( .A1(n623), .A2(n545), .ZN(n389) );
  NOR2_X1 U425 ( .A1(G902), .A2(n742), .ZN(n528) );
  NAND2_X1 U426 ( .A1(n406), .A2(n621), .ZN(n491) );
  XNOR2_X1 U427 ( .A(n585), .B(KEYINPUT92), .ZN(n406) );
  XNOR2_X1 U428 ( .A(G116), .B(G137), .ZN(n568) );
  XOR2_X1 U429 ( .A(KEYINPUT70), .B(KEYINPUT5), .Z(n569) );
  NOR2_X1 U430 ( .A1(G953), .A2(G237), .ZN(n570) );
  NAND2_X1 U431 ( .A1(n467), .A2(n468), .ZN(n464) );
  XOR2_X1 U432 ( .A(KEYINPUT75), .B(KEYINPUT85), .Z(n541) );
  XNOR2_X1 U433 ( .A(n471), .B(n538), .ZN(n494) );
  XNOR2_X1 U434 ( .A(n472), .B(KEYINPUT74), .ZN(n471) );
  XNOR2_X1 U435 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n472) );
  OR2_X1 U436 ( .A1(G902), .A2(G237), .ZN(n544) );
  BUF_X1 U437 ( .A(n618), .Z(n456) );
  NOR2_X1 U438 ( .A1(n663), .A2(n662), .ZN(n583) );
  NAND2_X1 U439 ( .A1(n392), .A2(n390), .ZN(n610) );
  AND2_X1 U440 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U441 ( .A1(n395), .A2(n638), .ZN(n393) );
  NAND2_X1 U442 ( .A1(n610), .A2(n654), .ZN(n618) );
  AND2_X1 U443 ( .A1(n723), .A2(n423), .ZN(n422) );
  XNOR2_X1 U444 ( .A(n536), .B(n495), .ZN(n751) );
  XNOR2_X1 U445 ( .A(n448), .B(n447), .ZN(n495) );
  INV_X1 U446 ( .A(n551), .ZN(n447) );
  NAND2_X1 U447 ( .A1(n464), .A2(n460), .ZN(n748) );
  AND2_X1 U448 ( .A1(n466), .A2(n465), .ZN(n460) );
  XNOR2_X1 U449 ( .A(n381), .B(n377), .ZN(n376) );
  XNOR2_X1 U450 ( .A(n517), .B(n516), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n379), .B(n378), .ZN(n377) );
  XOR2_X1 U452 ( .A(G140), .B(G131), .Z(n548) );
  XNOR2_X1 U453 ( .A(G143), .B(G113), .ZN(n547) );
  XNOR2_X1 U454 ( .A(n551), .B(n550), .ZN(n387) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n384) );
  INV_X1 U456 ( .A(KEYINPUT11), .ZN(n385) );
  NAND2_X1 U457 ( .A1(n570), .A2(G214), .ZN(n386) );
  NAND2_X1 U458 ( .A1(G214), .A2(n544), .ZN(n654) );
  XNOR2_X1 U459 ( .A(n609), .B(KEYINPUT39), .ZN(n632) );
  NOR2_X1 U460 ( .A1(n611), .A2(n651), .ZN(n609) );
  NOR2_X1 U461 ( .A1(n682), .A2(n439), .ZN(n402) );
  INV_X1 U462 ( .A(KEYINPUT6), .ZN(n451) );
  XNOR2_X1 U463 ( .A(n599), .B(KEYINPUT1), .ZN(n663) );
  XNOR2_X1 U464 ( .A(KEYINPUT68), .B(KEYINPUT22), .ZN(n559) );
  XNOR2_X1 U465 ( .A(n485), .B(n483), .ZN(n742) );
  XNOR2_X1 U466 ( .A(n524), .B(n514), .ZN(n485) );
  XNOR2_X1 U467 ( .A(n762), .B(n484), .ZN(n483) );
  XNOR2_X1 U468 ( .A(n411), .B(n567), .ZN(n401) );
  NOR2_X1 U469 ( .A1(G952), .A2(n764), .ZN(n744) );
  INV_X1 U470 ( .A(n665), .ZN(n429) );
  INV_X1 U471 ( .A(KEYINPUT45), .ZN(n469) );
  NAND2_X1 U472 ( .A1(n543), .A2(n525), .ZN(n391) );
  XNOR2_X1 U473 ( .A(n598), .B(KEYINPUT66), .ZN(n615) );
  AND2_X1 U474 ( .A1(n579), .A2(n360), .ZN(n598) );
  INV_X1 U475 ( .A(n722), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n380), .B(KEYINPUT98), .ZN(n379) );
  INV_X1 U477 ( .A(KEYINPUT96), .ZN(n380) );
  XNOR2_X1 U478 ( .A(G134), .B(KEYINPUT97), .ZN(n378) );
  XNOR2_X1 U479 ( .A(n396), .B(n478), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n572), .B(n573), .ZN(n478) );
  XNOR2_X1 U481 ( .A(n560), .B(n367), .ZN(n484) );
  NOR2_X1 U482 ( .A1(n748), .A2(n635), .ZN(n636) );
  NAND2_X1 U483 ( .A1(n461), .A2(n464), .ZN(n410) );
  XNOR2_X1 U484 ( .A(n560), .B(n404), .ZN(n757) );
  INV_X1 U485 ( .A(KEYINPUT88), .ZN(n404) );
  XNOR2_X1 U486 ( .A(G107), .B(G104), .ZN(n565) );
  XNOR2_X1 U487 ( .A(n409), .B(n407), .ZN(n563) );
  XNOR2_X1 U488 ( .A(KEYINPUT73), .B(KEYINPUT89), .ZN(n409) );
  NOR2_X1 U489 ( .A1(n408), .A2(G953), .ZN(n407) );
  INV_X1 U490 ( .A(G227), .ZN(n408) );
  XNOR2_X1 U491 ( .A(n562), .B(n493), .ZN(n492) );
  XNOR2_X1 U492 ( .A(n494), .B(n542), .ZN(n493) );
  XNOR2_X1 U493 ( .A(n382), .B(n602), .ZN(n681) );
  XNOR2_X1 U494 ( .A(n601), .B(n600), .ZN(n602) );
  NOR2_X1 U495 ( .A1(n651), .A2(n383), .ZN(n382) );
  XNOR2_X1 U496 ( .A(n374), .B(n373), .ZN(n617) );
  INV_X1 U497 ( .A(KEYINPUT99), .ZN(n373) );
  NAND2_X1 U498 ( .A1(n445), .A2(n586), .ZN(n374) );
  NOR2_X1 U499 ( .A1(n456), .A2(n370), .ZN(n506) );
  AND2_X1 U500 ( .A1(n608), .A2(n606), .ZN(n455) );
  XNOR2_X1 U501 ( .A(KEYINPUT30), .B(KEYINPUT105), .ZN(n604) );
  AND2_X1 U502 ( .A1(n480), .A2(n479), .ZN(n622) );
  INV_X1 U503 ( .A(n599), .ZN(n479) );
  XNOR2_X1 U504 ( .A(n482), .B(n481), .ZN(n480) );
  INV_X1 U505 ( .A(KEYINPUT28), .ZN(n481) );
  XNOR2_X1 U506 ( .A(n617), .B(n372), .ZN(n510) );
  INV_X1 U507 ( .A(KEYINPUT102), .ZN(n372) );
  NOR2_X1 U508 ( .A1(n662), .A2(n599), .ZN(n607) );
  XOR2_X1 U509 ( .A(n520), .B(n519), .Z(n640) );
  XNOR2_X1 U510 ( .A(n518), .B(n376), .ZN(n519) );
  XNOR2_X1 U511 ( .A(n387), .B(n384), .ZN(n552) );
  NAND2_X1 U512 ( .A1(n375), .A2(n631), .ZN(n723) );
  XNOR2_X1 U513 ( .A(n630), .B(KEYINPUT104), .ZN(n375) );
  XNOR2_X1 U514 ( .A(n450), .B(KEYINPUT40), .ZN(n775) );
  NOR2_X1 U515 ( .A1(n632), .A2(n617), .ZN(n450) );
  NAND2_X1 U516 ( .A1(n476), .A2(n582), .ZN(n475) );
  XNOR2_X1 U517 ( .A(n402), .B(KEYINPUT34), .ZN(n476) );
  INV_X1 U518 ( .A(KEYINPUT32), .ZN(n436) );
  XNOR2_X1 U519 ( .A(n413), .B(n412), .ZN(n715) );
  INV_X1 U520 ( .A(KEYINPUT31), .ZN(n412) );
  NAND2_X1 U521 ( .A1(n433), .A2(n434), .ZN(n415) );
  AND2_X1 U522 ( .A1(n418), .A2(n417), .ZN(n416) );
  NAND2_X1 U523 ( .A1(n663), .A2(n474), .ZN(n473) );
  NOR2_X1 U524 ( .A1(n614), .A2(n579), .ZN(n474) );
  XNOR2_X1 U525 ( .A(n740), .B(n452), .ZN(n743) );
  XNOR2_X1 U526 ( .A(n742), .B(n741), .ZN(n452) );
  XNOR2_X1 U527 ( .A(n730), .B(n449), .ZN(n733) );
  XNOR2_X1 U528 ( .A(n732), .B(n731), .ZN(n449) );
  XOR2_X1 U529 ( .A(G902), .B(KEYINPUT15), .Z(n638) );
  XNOR2_X1 U530 ( .A(KEYINPUT77), .B(n637), .ZN(n356) );
  OR2_X1 U531 ( .A1(n578), .A2(n473), .ZN(n489) );
  AND2_X1 U532 ( .A1(n489), .A2(KEYINPUT82), .ZN(n357) );
  AND2_X1 U533 ( .A1(n398), .A2(n459), .ZN(n358) );
  XOR2_X1 U534 ( .A(KEYINPUT91), .B(G472), .Z(n359) );
  AND2_X1 U535 ( .A1(n665), .A2(n606), .ZN(n360) );
  XOR2_X1 U536 ( .A(n527), .B(KEYINPUT25), .Z(n361) );
  AND2_X1 U537 ( .A1(n410), .A2(n638), .ZN(n363) );
  AND2_X1 U538 ( .A1(n425), .A2(n723), .ZN(n364) );
  NOR2_X1 U539 ( .A1(n663), .A2(n614), .ZN(n365) );
  AND2_X1 U540 ( .A1(n357), .A2(n491), .ZN(n366) );
  XOR2_X1 U541 ( .A(G128), .B(G119), .Z(n367) );
  INV_X1 U542 ( .A(n543), .ZN(n395) );
  AND2_X1 U543 ( .A1(n579), .A2(n437), .ZN(n368) );
  AND2_X1 U544 ( .A1(n364), .A2(n356), .ZN(n369) );
  NAND2_X1 U545 ( .A1(n416), .A2(n415), .ZN(n774) );
  XOR2_X1 U546 ( .A(KEYINPUT36), .B(KEYINPUT108), .Z(n370) );
  INV_X1 U547 ( .A(KEYINPUT100), .ZN(n437) );
  INV_X1 U548 ( .A(KEYINPUT82), .ZN(n490) );
  AND2_X1 U549 ( .A1(n490), .A2(KEYINPUT44), .ZN(n371) );
  INV_X1 U550 ( .A(n681), .ZN(n430) );
  NAND2_X1 U551 ( .A1(n650), .A2(n654), .ZN(n383) );
  XNOR2_X2 U552 ( .A(n388), .B(n559), .ZN(n578) );
  NAND2_X1 U553 ( .A1(n558), .A2(n557), .ZN(n388) );
  XNOR2_X2 U554 ( .A(n389), .B(n440), .ZN(n558) );
  OR2_X1 U555 ( .A1(n724), .A2(n391), .ZN(n390) );
  NAND2_X1 U556 ( .A1(n724), .A2(n395), .ZN(n394) );
  XNOR2_X1 U557 ( .A(n492), .B(n751), .ZN(n724) );
  NAND2_X1 U558 ( .A1(n773), .A2(n774), .ZN(n444) );
  XNOR2_X1 U559 ( .A(n419), .B(n436), .ZN(n773) );
  XNOR2_X1 U560 ( .A(n401), .B(n396), .ZN(n732) );
  NAND2_X1 U561 ( .A1(n397), .A2(n591), .ZN(n592) );
  NAND2_X1 U562 ( .A1(n772), .A2(n371), .ZN(n398) );
  NAND2_X1 U563 ( .A1(n583), .A2(n614), .ZN(n403) );
  OR2_X2 U564 ( .A1(n421), .A2(G902), .ZN(n477) );
  INV_X1 U565 ( .A(n410), .ZN(n648) );
  XNOR2_X1 U566 ( .A(n757), .B(n566), .ZN(n411) );
  INV_X1 U567 ( .A(n558), .ZN(n439) );
  NAND2_X1 U568 ( .A1(n414), .A2(n558), .ZN(n413) );
  INV_X1 U569 ( .A(n671), .ZN(n414) );
  NAND2_X1 U570 ( .A1(n578), .A2(KEYINPUT100), .ZN(n417) );
  OR2_X1 U571 ( .A1(n435), .A2(n437), .ZN(n418) );
  NAND2_X1 U572 ( .A1(n365), .A2(n579), .ZN(n420) );
  XNOR2_X1 U573 ( .A(n421), .B(n694), .ZN(n695) );
  XNOR2_X1 U574 ( .A(n424), .B(n497), .ZN(n425) );
  NAND2_X1 U575 ( .A1(n426), .A2(n427), .ZN(n424) );
  XNOR2_X1 U576 ( .A(n500), .B(KEYINPUT46), .ZN(n426) );
  NAND2_X1 U577 ( .A1(n428), .A2(n665), .ZN(n662) );
  INV_X1 U578 ( .A(n579), .ZN(n428) );
  AND2_X1 U579 ( .A1(n429), .A2(n579), .ZN(n666) );
  XNOR2_X2 U580 ( .A(n528), .B(n361), .ZN(n579) );
  AND2_X1 U581 ( .A1(n574), .A2(n368), .ZN(n433) );
  INV_X1 U582 ( .A(n578), .ZN(n434) );
  AND2_X1 U583 ( .A1(n574), .A2(n579), .ZN(n435) );
  AND2_X1 U584 ( .A1(n558), .A2(n438), .ZN(n584) );
  INV_X1 U585 ( .A(n668), .ZN(n438) );
  NOR2_X2 U586 ( .A1(n697), .A2(n744), .ZN(n453) );
  NOR2_X2 U587 ( .A1(n729), .A2(n744), .ZN(n454) );
  NAND2_X1 U588 ( .A1(n442), .A2(n644), .ZN(n441) );
  INV_X1 U589 ( .A(n636), .ZN(n442) );
  NAND2_X1 U590 ( .A1(n739), .A2(G478), .ZN(n639) );
  NAND2_X1 U591 ( .A1(n575), .A2(n654), .ZN(n605) );
  XNOR2_X2 U592 ( .A(n477), .B(n359), .ZN(n575) );
  XNOR2_X2 U593 ( .A(n539), .B(KEYINPUT4), .ZN(n760) );
  XNOR2_X2 U594 ( .A(n443), .B(G128), .ZN(n539) );
  XNOR2_X2 U595 ( .A(n444), .B(KEYINPUT83), .ZN(n590) );
  INV_X1 U596 ( .A(n586), .ZN(n587) );
  INV_X1 U597 ( .A(n588), .ZN(n445) );
  XNOR2_X2 U598 ( .A(n546), .B(n446), .ZN(n588) );
  XNOR2_X1 U599 ( .A(n553), .B(n552), .ZN(n735) );
  XNOR2_X1 U600 ( .A(n535), .B(n537), .ZN(n448) );
  NAND2_X1 U601 ( .A1(n592), .A2(n469), .ZN(n465) );
  NAND2_X1 U602 ( .A1(n366), .A2(n487), .ZN(n458) );
  XNOR2_X1 U603 ( .A(n453), .B(n698), .ZN(G57) );
  XNOR2_X1 U604 ( .A(n454), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U605 ( .A1(n607), .A2(n455), .ZN(n611) );
  NOR2_X2 U606 ( .A1(n590), .A2(n576), .ZN(n577) );
  NAND2_X1 U607 ( .A1(n465), .A2(n369), .ZN(n462) );
  XNOR2_X1 U608 ( .A(n457), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U609 ( .A1(n738), .A2(n744), .ZN(n457) );
  XNOR2_X2 U610 ( .A(n618), .B(KEYINPUT19), .ZN(n623) );
  NAND2_X1 U611 ( .A1(n486), .A2(n490), .ZN(n459) );
  NAND2_X1 U612 ( .A1(n593), .A2(n469), .ZN(n466) );
  NOR2_X1 U613 ( .A1(n463), .A2(n462), .ZN(n461) );
  INV_X1 U614 ( .A(n466), .ZN(n463) );
  INV_X1 U615 ( .A(n593), .ZN(n467) );
  NOR2_X1 U616 ( .A1(n592), .A2(n469), .ZN(n468) );
  XNOR2_X2 U617 ( .A(n475), .B(KEYINPUT35), .ZN(n772) );
  NAND2_X1 U618 ( .A1(n615), .A2(n668), .ZN(n482) );
  NAND2_X1 U619 ( .A1(n772), .A2(KEYINPUT44), .ZN(n487) );
  NAND2_X1 U620 ( .A1(n491), .A2(n489), .ZN(n486) );
  INV_X1 U621 ( .A(n489), .ZN(n488) );
  INV_X1 U622 ( .A(KEYINPUT48), .ZN(n497) );
  NAND2_X1 U623 ( .A1(n625), .A2(n499), .ZN(n498) );
  NAND2_X1 U624 ( .A1(n713), .A2(n370), .ZN(n501) );
  NAND2_X1 U625 ( .A1(n503), .A2(n370), .ZN(n502) );
  NAND2_X1 U626 ( .A1(n509), .A2(n508), .ZN(n503) );
  NAND2_X1 U627 ( .A1(n510), .A2(n509), .ZN(n626) );
  NAND2_X1 U628 ( .A1(n510), .A2(n505), .ZN(n504) );
  AND2_X1 U629 ( .A1(n509), .A2(n506), .ZN(n505) );
  INV_X1 U630 ( .A(n456), .ZN(n508) );
  XNOR2_X1 U631 ( .A(n610), .B(KEYINPUT38), .ZN(n651) );
  XOR2_X1 U632 ( .A(n523), .B(n522), .Z(n514) );
  AND2_X1 U633 ( .A1(G210), .A2(n570), .ZN(n515) );
  INV_X1 U634 ( .A(n651), .ZN(n655) );
  INV_X1 U635 ( .A(KEYINPUT71), .ZN(n634) );
  XNOR2_X1 U636 ( .A(n763), .B(n634), .ZN(n635) );
  XNOR2_X1 U637 ( .A(n571), .B(n515), .ZN(n572) );
  AND2_X1 U638 ( .A1(n650), .A2(n665), .ZN(n557) );
  INV_X1 U639 ( .A(KEYINPUT80), .ZN(n633) );
  XNOR2_X1 U640 ( .A(n758), .B(G146), .ZN(n561) );
  INV_X1 U641 ( .A(KEYINPUT59), .ZN(n734) );
  BUF_X1 U642 ( .A(n575), .Z(n668) );
  XNOR2_X1 U643 ( .A(n693), .B(n692), .ZN(G75) );
  NAND2_X1 U644 ( .A1(n521), .A2(G217), .ZN(n520) );
  XNOR2_X1 U645 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n516) );
  XNOR2_X1 U646 ( .A(G122), .B(KEYINPUT95), .ZN(n517) );
  XNOR2_X1 U647 ( .A(n539), .B(n535), .ZN(n518) );
  NAND2_X1 U648 ( .A1(G221), .A2(n521), .ZN(n524) );
  XOR2_X1 U649 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n523) );
  XNOR2_X1 U650 ( .A(G110), .B(KEYINPUT90), .ZN(n522) );
  INV_X1 U651 ( .A(n638), .ZN(n525) );
  NAND2_X1 U652 ( .A1(G234), .A2(n525), .ZN(n526) );
  XNOR2_X1 U653 ( .A(KEYINPUT20), .B(n526), .ZN(n555) );
  NAND2_X1 U654 ( .A1(n555), .A2(G217), .ZN(n527) );
  NAND2_X1 U655 ( .A1(G237), .A2(G234), .ZN(n529) );
  XNOR2_X1 U656 ( .A(n529), .B(KEYINPUT14), .ZN(n531) );
  NAND2_X1 U657 ( .A1(n531), .A2(G952), .ZN(n530) );
  XNOR2_X1 U658 ( .A(n530), .B(KEYINPUT87), .ZN(n679) );
  NAND2_X1 U659 ( .A1(n679), .A2(n764), .ZN(n597) );
  NAND2_X1 U660 ( .A1(G902), .A2(n531), .ZN(n594) );
  INV_X1 U661 ( .A(n594), .ZN(n532) );
  NOR2_X1 U662 ( .A1(G898), .A2(n764), .ZN(n753) );
  NAND2_X1 U663 ( .A1(n532), .A2(n753), .ZN(n533) );
  NAND2_X1 U664 ( .A1(n597), .A2(n533), .ZN(n545) );
  XNOR2_X1 U665 ( .A(KEYINPUT69), .B(KEYINPUT16), .ZN(n537) );
  XNOR2_X1 U666 ( .A(G113), .B(KEYINPUT67), .ZN(n534) );
  XNOR2_X1 U667 ( .A(n355), .B(n534), .ZN(n573) );
  XOR2_X1 U668 ( .A(KEYINPUT86), .B(G110), .Z(n564) );
  XNOR2_X1 U669 ( .A(n573), .B(n564), .ZN(n536) );
  XOR2_X1 U670 ( .A(G122), .B(G104), .Z(n551) );
  NAND2_X1 U671 ( .A1(G224), .A2(n764), .ZN(n540) );
  XNOR2_X1 U672 ( .A(n541), .B(n540), .ZN(n542) );
  NAND2_X1 U673 ( .A1(G210), .A2(n544), .ZN(n543) );
  XNOR2_X1 U674 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U675 ( .A(n762), .B(n549), .ZN(n553) );
  XOR2_X1 U676 ( .A(KEYINPUT93), .B(KEYINPUT12), .Z(n550) );
  XNOR2_X1 U677 ( .A(KEYINPUT94), .B(KEYINPUT13), .ZN(n554) );
  NOR2_X1 U678 ( .A1(n588), .A2(n586), .ZN(n650) );
  NAND2_X1 U679 ( .A1(n555), .A2(G221), .ZN(n556) );
  XOR2_X1 U680 ( .A(KEYINPUT21), .B(n556), .Z(n665) );
  XOR2_X1 U681 ( .A(G134), .B(G131), .Z(n758) );
  XOR2_X1 U682 ( .A(n563), .B(KEYINPUT72), .Z(n567) );
  XNOR2_X1 U683 ( .A(n565), .B(n564), .ZN(n566) );
  INV_X1 U684 ( .A(n663), .ZN(n627) );
  XNOR2_X1 U685 ( .A(n569), .B(n568), .ZN(n571) );
  NOR2_X1 U686 ( .A1(n627), .A2(n668), .ZN(n574) );
  INV_X1 U687 ( .A(KEYINPUT44), .ZN(n576) );
  XNOR2_X1 U688 ( .A(n577), .B(KEYINPUT64), .ZN(n593) );
  XOR2_X1 U689 ( .A(KEYINPUT84), .B(KEYINPUT33), .Z(n580) );
  NAND2_X1 U690 ( .A1(n586), .A2(n588), .ZN(n581) );
  XOR2_X1 U691 ( .A(n581), .B(KEYINPUT101), .Z(n613) );
  XOR2_X1 U692 ( .A(KEYINPUT76), .B(n613), .Z(n582) );
  NAND2_X1 U693 ( .A1(n668), .A2(n583), .ZN(n671) );
  NAND2_X1 U694 ( .A1(n607), .A2(n584), .ZN(n701) );
  NAND2_X1 U695 ( .A1(n715), .A2(n701), .ZN(n585) );
  NAND2_X1 U696 ( .A1(n588), .A2(n587), .ZN(n716) );
  NAND2_X1 U697 ( .A1(n617), .A2(n716), .ZN(n621) );
  NOR2_X1 U698 ( .A1(n772), .A2(KEYINPUT44), .ZN(n589) );
  NAND2_X1 U699 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U700 ( .A1(G900), .A2(n594), .ZN(n595) );
  NAND2_X1 U701 ( .A1(G953), .A2(n595), .ZN(n596) );
  NAND2_X1 U702 ( .A1(n597), .A2(n596), .ZN(n606) );
  XNOR2_X1 U703 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n601) );
  INV_X1 U704 ( .A(KEYINPUT106), .ZN(n600) );
  XNOR2_X1 U705 ( .A(n605), .B(n604), .ZN(n608) );
  INV_X1 U706 ( .A(n610), .ZN(n631) );
  OR2_X1 U707 ( .A1(n631), .A2(n611), .ZN(n612) );
  NOR2_X1 U708 ( .A1(n613), .A2(n612), .ZN(n708) );
  INV_X1 U709 ( .A(n621), .ZN(n657) );
  NAND2_X1 U710 ( .A1(n623), .A2(n622), .ZN(n709) );
  XNOR2_X1 U711 ( .A(n624), .B(KEYINPUT47), .ZN(n625) );
  NOR2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n654), .A2(n628), .ZN(n629) );
  XNOR2_X1 U714 ( .A(n629), .B(KEYINPUT43), .ZN(n630) );
  NOR2_X1 U715 ( .A1(n716), .A2(n632), .ZN(n722) );
  XNOR2_X2 U716 ( .A(n362), .B(n633), .ZN(n763) );
  INV_X1 U717 ( .A(KEYINPUT2), .ZN(n644) );
  OR2_X1 U718 ( .A1(n644), .A2(n722), .ZN(n637) );
  XNOR2_X1 U719 ( .A(n639), .B(n640), .ZN(n641) );
  NOR2_X2 U720 ( .A1(n641), .A2(n744), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n642), .B(KEYINPUT122), .ZN(G63) );
  NAND2_X1 U722 ( .A1(n644), .A2(n763), .ZN(n643) );
  XNOR2_X1 U723 ( .A(n643), .B(KEYINPUT78), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n644), .A2(n748), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U726 ( .A(KEYINPUT79), .B(n649), .ZN(n688) );
  INV_X1 U727 ( .A(n650), .ZN(n653) );
  NOR2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n652) );
  NOR2_X1 U729 ( .A1(n653), .A2(n652), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U733 ( .A(KEYINPUT117), .B(n660), .Z(n661) );
  NOR2_X1 U734 ( .A1(n682), .A2(n661), .ZN(n677) );
  NAND2_X1 U735 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U736 ( .A(n664), .B(KEYINPUT50), .ZN(n670) );
  XOR2_X1 U737 ( .A(KEYINPUT49), .B(n666), .Z(n667) );
  NOR2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n672) );
  NAND2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U741 ( .A(KEYINPUT51), .B(n673), .ZN(n674) );
  NOR2_X1 U742 ( .A1(n681), .A2(n674), .ZN(n675) );
  XNOR2_X1 U743 ( .A(n675), .B(KEYINPUT116), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U745 ( .A(KEYINPUT52), .B(n678), .Z(n680) );
  NAND2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n685) );
  NOR2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U748 ( .A(KEYINPUT118), .B(n683), .Z(n684) );
  NAND2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U750 ( .A(n686), .B(KEYINPUT119), .ZN(n687) );
  NAND2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U752 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n691) );
  INV_X1 U753 ( .A(KEYINPUT120), .ZN(n690) );
  XNOR2_X1 U754 ( .A(n691), .B(n690), .ZN(n692) );
  INV_X1 U755 ( .A(KEYINPUT63), .ZN(n698) );
  NAND2_X1 U756 ( .A1(n739), .A2(G472), .ZN(n696) );
  XOR2_X1 U757 ( .A(KEYINPUT62), .B(KEYINPUT109), .Z(n694) );
  XNOR2_X1 U758 ( .A(n696), .B(n695), .ZN(n697) );
  XOR2_X1 U759 ( .A(G101), .B(n488), .Z(G3) );
  NOR2_X1 U760 ( .A1(n713), .A2(n701), .ZN(n699) );
  XOR2_X1 U761 ( .A(KEYINPUT110), .B(n699), .Z(n700) );
  XNOR2_X1 U762 ( .A(G104), .B(n700), .ZN(G6) );
  NOR2_X1 U763 ( .A1(n701), .A2(n716), .ZN(n705) );
  XOR2_X1 U764 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n703) );
  XNOR2_X1 U765 ( .A(G107), .B(KEYINPUT111), .ZN(n702) );
  XNOR2_X1 U766 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U767 ( .A(n705), .B(n704), .ZN(G9) );
  NOR2_X1 U768 ( .A1(n716), .A2(n709), .ZN(n707) );
  XNOR2_X1 U769 ( .A(G128), .B(KEYINPUT29), .ZN(n706) );
  XNOR2_X1 U770 ( .A(n707), .B(n706), .ZN(G30) );
  XOR2_X1 U771 ( .A(G143), .B(n708), .Z(G45) );
  NOR2_X1 U772 ( .A1(n713), .A2(n709), .ZN(n711) );
  XNOR2_X1 U773 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n710) );
  XNOR2_X1 U774 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U775 ( .A(G146), .B(n712), .ZN(G48) );
  NOR2_X1 U776 ( .A1(n713), .A2(n715), .ZN(n714) );
  XOR2_X1 U777 ( .A(G113), .B(n714), .Z(G15) );
  NOR2_X1 U778 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U779 ( .A(KEYINPUT114), .B(n717), .Z(n718) );
  XNOR2_X1 U780 ( .A(G116), .B(n718), .ZN(G18) );
  XNOR2_X1 U781 ( .A(KEYINPUT115), .B(KEYINPUT37), .ZN(n720) );
  XNOR2_X1 U782 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U783 ( .A(G125), .B(n721), .ZN(G27) );
  XOR2_X1 U784 ( .A(G134), .B(n722), .Z(G36) );
  XNOR2_X1 U785 ( .A(G140), .B(n723), .ZN(G42) );
  NAND2_X1 U786 ( .A1(n739), .A2(G210), .ZN(n728) );
  BUF_X1 U787 ( .A(n724), .Z(n726) );
  XOR2_X1 U788 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n725) );
  XNOR2_X1 U789 ( .A(n728), .B(n727), .ZN(n729) );
  XOR2_X1 U790 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n731) );
  NAND2_X1 U791 ( .A1(n739), .A2(G469), .ZN(n730) );
  NOR2_X1 U792 ( .A1(n744), .A2(n733), .ZN(G54) );
  NAND2_X1 U793 ( .A1(n739), .A2(G475), .ZN(n737) );
  XNOR2_X1 U794 ( .A(n737), .B(n736), .ZN(n738) );
  XOR2_X1 U795 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n741) );
  NAND2_X1 U796 ( .A1(n739), .A2(G217), .ZN(n740) );
  NOR2_X1 U797 ( .A1(n744), .A2(n743), .ZN(G66) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n745) );
  XNOR2_X1 U799 ( .A(KEYINPUT61), .B(n745), .ZN(n746) );
  NAND2_X1 U800 ( .A1(n746), .A2(G898), .ZN(n747) );
  XNOR2_X1 U801 ( .A(n747), .B(KEYINPUT125), .ZN(n750) );
  NOR2_X1 U802 ( .A1(n748), .A2(G953), .ZN(n749) );
  NOR2_X1 U803 ( .A1(n750), .A2(n749), .ZN(n756) );
  XOR2_X1 U804 ( .A(n751), .B(G101), .Z(n752) );
  NOR2_X1 U805 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U806 ( .A(KEYINPUT126), .B(n754), .Z(n755) );
  XNOR2_X1 U807 ( .A(n756), .B(n755), .ZN(G69) );
  XOR2_X1 U808 ( .A(n758), .B(n757), .Z(n759) );
  XNOR2_X1 U809 ( .A(n760), .B(n759), .ZN(n761) );
  XOR2_X1 U810 ( .A(n762), .B(n761), .Z(n766) );
  XOR2_X1 U811 ( .A(n763), .B(n766), .Z(n765) );
  NAND2_X1 U812 ( .A1(n765), .A2(n764), .ZN(n770) );
  XOR2_X1 U813 ( .A(G227), .B(n766), .Z(n767) );
  NAND2_X1 U814 ( .A1(n767), .A2(G900), .ZN(n768) );
  NAND2_X1 U815 ( .A1(n768), .A2(G953), .ZN(n769) );
  NAND2_X1 U816 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U817 ( .A(KEYINPUT127), .B(n771), .Z(G72) );
  XOR2_X1 U818 ( .A(n772), .B(G122), .Z(G24) );
  XNOR2_X1 U819 ( .A(G119), .B(n773), .ZN(G21) );
  XNOR2_X1 U820 ( .A(G110), .B(n774), .ZN(G12) );
  XOR2_X1 U821 ( .A(n775), .B(G131), .Z(G33) );
  XOR2_X1 U822 ( .A(n776), .B(G137), .Z(G39) );
endmodule

