

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U323 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U324 ( .A(KEYINPUT54), .B(KEYINPUT116), .ZN(n409) );
  XNOR2_X1 U325 ( .A(n455), .B(n454), .ZN(n563) );
  XNOR2_X1 U326 ( .A(n427), .B(KEYINPUT55), .ZN(n445) );
  XNOR2_X1 U327 ( .A(n429), .B(n428), .ZN(n430) );
  INV_X1 U328 ( .A(KEYINPUT32), .ZN(n369) );
  XNOR2_X1 U329 ( .A(n431), .B(n430), .ZN(n435) );
  XNOR2_X1 U330 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U331 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n454) );
  XNOR2_X1 U332 ( .A(n408), .B(KEYINPUT48), .ZN(n539) );
  XNOR2_X1 U333 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U334 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U335 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U336 ( .A(n446), .B(G190GAT), .ZN(n447) );
  XNOR2_X1 U337 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U338 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n477), .B(n476), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT11), .B(G218GAT), .Z(n292) );
  XNOR2_X1 U341 ( .A(G134GAT), .B(G106GAT), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U343 ( .A(KEYINPUT77), .B(KEYINPUT10), .Z(n294) );
  XNOR2_X1 U344 ( .A(KEYINPUT66), .B(KEYINPUT9), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U346 ( .A(n296), .B(n295), .Z(n305) );
  XOR2_X1 U347 ( .A(KEYINPUT70), .B(KEYINPUT7), .Z(n298) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G29GAT), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U350 ( .A(KEYINPUT8), .B(n299), .Z(n355) );
  XNOR2_X1 U351 ( .A(G36GAT), .B(G190GAT), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n300), .B(KEYINPUT79), .ZN(n329) );
  XNOR2_X1 U353 ( .A(G50GAT), .B(G162GAT), .ZN(n425) );
  XNOR2_X1 U354 ( .A(n329), .B(n425), .ZN(n302) );
  NAND2_X1 U355 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n355), .B(n303), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U359 ( .A(n306), .B(KEYINPUT78), .Z(n310) );
  XOR2_X1 U360 ( .A(KEYINPUT74), .B(G92GAT), .Z(n308) );
  XNOR2_X1 U361 ( .A(G99GAT), .B(G85GAT), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n361) );
  XNOR2_X1 U363 ( .A(n361), .B(KEYINPUT65), .ZN(n309) );
  XOR2_X1 U364 ( .A(n310), .B(n309), .Z(n478) );
  XNOR2_X1 U365 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n311), .B(KEYINPUT2), .ZN(n419) );
  XOR2_X1 U367 ( .A(G134GAT), .B(KEYINPUT0), .Z(n428) );
  XOR2_X1 U368 ( .A(n419), .B(n428), .Z(n313) );
  NAND2_X1 U369 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n328) );
  XOR2_X1 U371 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n315) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(KEYINPUT1), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U374 ( .A(G57GAT), .B(KEYINPUT4), .Z(n317) );
  XNOR2_X1 U375 ( .A(KEYINPUT89), .B(KEYINPUT6), .ZN(n316) );
  XNOR2_X1 U376 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n326) );
  XOR2_X1 U378 ( .A(G85GAT), .B(G148GAT), .Z(n321) );
  XNOR2_X1 U379 ( .A(G120GAT), .B(G162GAT), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U381 ( .A(n322), .B(G127GAT), .Z(n324) );
  XOR2_X1 U382 ( .A(G113GAT), .B(G1GAT), .Z(n348) );
  XNOR2_X1 U383 ( .A(G29GAT), .B(n348), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U386 ( .A(n328), .B(n327), .Z(n512) );
  INV_X1 U387 ( .A(n512), .ZN(n469) );
  XOR2_X1 U388 ( .A(G8GAT), .B(G183GAT), .Z(n383) );
  XOR2_X1 U389 ( .A(KEYINPUT91), .B(n329), .Z(n333) );
  XOR2_X1 U390 ( .A(G64GAT), .B(KEYINPUT75), .Z(n331) );
  XNOR2_X1 U391 ( .A(G176GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n366) );
  XNOR2_X1 U393 ( .A(n366), .B(G92GAT), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U395 ( .A(n383), .B(n334), .Z(n336) );
  NAND2_X1 U396 ( .A1(G226GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n336), .B(n335), .ZN(n342) );
  XOR2_X1 U398 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n338) );
  XNOR2_X1 U399 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n338), .B(n337), .ZN(n431) );
  XOR2_X1 U401 ( .A(G211GAT), .B(KEYINPUT21), .Z(n340) );
  XNOR2_X1 U402 ( .A(G197GAT), .B(G218GAT), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n340), .B(n339), .ZN(n412) );
  XOR2_X1 U404 ( .A(n431), .B(n412), .Z(n341) );
  XOR2_X1 U405 ( .A(n342), .B(n341), .Z(n514) );
  INV_X1 U406 ( .A(n514), .ZN(n494) );
  XOR2_X1 U407 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n344) );
  XNOR2_X1 U408 ( .A(KEYINPUT71), .B(KEYINPUT29), .ZN(n343) );
  XNOR2_X1 U409 ( .A(n344), .B(n343), .ZN(n359) );
  XOR2_X1 U410 ( .A(G8GAT), .B(G197GAT), .Z(n346) );
  XNOR2_X1 U411 ( .A(G50GAT), .B(G36GAT), .ZN(n345) );
  XNOR2_X1 U412 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U413 ( .A(n347), .B(G15GAT), .Z(n350) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(n348), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U416 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n352) );
  NAND2_X1 U417 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U419 ( .A(n354), .B(n353), .Z(n357) );
  XOR2_X1 U420 ( .A(G141GAT), .B(G22GAT), .Z(n424) );
  XNOR2_X1 U421 ( .A(n355), .B(n424), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U423 ( .A(n359), .B(n358), .Z(n542) );
  INV_X1 U424 ( .A(n542), .ZN(n565) );
  XNOR2_X1 U425 ( .A(G106GAT), .B(G78GAT), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n360), .B(G148GAT), .ZN(n420) );
  XNOR2_X1 U427 ( .A(n420), .B(n361), .ZN(n374) );
  XOR2_X1 U428 ( .A(KEYINPUT76), .B(KEYINPUT33), .Z(n363) );
  NAND2_X1 U429 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U430 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U431 ( .A(n364), .B(KEYINPUT31), .Z(n368) );
  XNOR2_X1 U432 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n365), .B(KEYINPUT72), .ZN(n386) );
  XNOR2_X1 U434 ( .A(n366), .B(n386), .ZN(n367) );
  XNOR2_X1 U435 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U436 ( .A(G120GAT), .B(G71GAT), .Z(n439) );
  XNOR2_X1 U437 ( .A(n439), .B(KEYINPUT73), .ZN(n370) );
  XOR2_X1 U438 ( .A(n374), .B(n373), .Z(n571) );
  INV_X1 U439 ( .A(n571), .ZN(n449) );
  XNOR2_X1 U440 ( .A(KEYINPUT36), .B(n478), .ZN(n582) );
  XOR2_X1 U441 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n376) );
  XNOR2_X1 U442 ( .A(KEYINPUT14), .B(KEYINPUT85), .ZN(n375) );
  XNOR2_X1 U443 ( .A(n376), .B(n375), .ZN(n396) );
  XOR2_X1 U444 ( .A(KEYINPUT80), .B(KEYINPUT84), .Z(n378) );
  XNOR2_X1 U445 ( .A(KEYINPUT71), .B(KEYINPUT12), .ZN(n377) );
  XNOR2_X1 U446 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U447 ( .A(KEYINPUT82), .B(G64GAT), .Z(n380) );
  XNOR2_X1 U448 ( .A(G22GAT), .B(G1GAT), .ZN(n379) );
  XNOR2_X1 U449 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n382), .B(n381), .ZN(n394) );
  XOR2_X1 U451 ( .A(n383), .B(G155GAT), .Z(n385) );
  XOR2_X1 U452 ( .A(G15GAT), .B(G127GAT), .Z(n429) );
  XNOR2_X1 U453 ( .A(n429), .B(G78GAT), .ZN(n384) );
  XNOR2_X1 U454 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U455 ( .A(n386), .B(KEYINPUT15), .Z(n388) );
  NAND2_X1 U456 ( .A1(G231GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U458 ( .A(n390), .B(n389), .Z(n392) );
  XNOR2_X1 U459 ( .A(G71GAT), .B(G211GAT), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U462 ( .A(n396), .B(n395), .Z(n548) );
  INV_X1 U463 ( .A(n548), .ZN(n576) );
  NOR2_X1 U464 ( .A1(n582), .A2(n576), .ZN(n397) );
  XOR2_X1 U465 ( .A(KEYINPUT45), .B(n397), .Z(n398) );
  NOR2_X1 U466 ( .A1(n449), .A2(n398), .ZN(n399) );
  NAND2_X1 U467 ( .A1(n565), .A2(n399), .ZN(n407) );
  INV_X1 U468 ( .A(n478), .ZN(n551) );
  XOR2_X1 U469 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n400) );
  XOR2_X1 U470 ( .A(n571), .B(n400), .Z(n544) );
  NAND2_X1 U471 ( .A1(n542), .A2(n544), .ZN(n401) );
  XNOR2_X1 U472 ( .A(n401), .B(KEYINPUT46), .ZN(n402) );
  NAND2_X1 U473 ( .A1(n402), .A2(n576), .ZN(n403) );
  NOR2_X1 U474 ( .A1(n551), .A2(n403), .ZN(n405) );
  XNOR2_X1 U475 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n404) );
  XNOR2_X1 U476 ( .A(n405), .B(n404), .ZN(n406) );
  NAND2_X1 U477 ( .A1(n407), .A2(n406), .ZN(n408) );
  NAND2_X1 U478 ( .A1(n494), .A2(n539), .ZN(n410) );
  NOR2_X1 U479 ( .A1(n469), .A2(n411), .ZN(n564) );
  XOR2_X1 U480 ( .A(n412), .B(G204GAT), .Z(n414) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U482 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U483 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n416) );
  XNOR2_X1 U484 ( .A(KEYINPUT22), .B(KEYINPUT88), .ZN(n415) );
  XNOR2_X1 U485 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U486 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U487 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U488 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n460) );
  NAND2_X1 U491 ( .A1(n564), .A2(n460), .ZN(n427) );
  XOR2_X1 U492 ( .A(G176GAT), .B(G183GAT), .Z(n433) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U495 ( .A(n435), .B(n434), .Z(n442) );
  XOR2_X1 U496 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n437) );
  XNOR2_X1 U497 ( .A(G190GAT), .B(KEYINPUT87), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U499 ( .A(G113GAT), .B(n438), .ZN(n440) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(G99GAT), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n524) );
  INV_X1 U502 ( .A(n524), .ZN(n473) );
  NAND2_X1 U503 ( .A1(n445), .A2(n473), .ZN(n561) );
  NOR2_X1 U504 ( .A1(n478), .A2(n561), .ZN(n448) );
  XNOR2_X1 U505 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n446) );
  XOR2_X1 U506 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n468) );
  NOR2_X1 U507 ( .A1(n449), .A2(n565), .ZN(n482) );
  NAND2_X1 U508 ( .A1(n473), .A2(n494), .ZN(n450) );
  XOR2_X1 U509 ( .A(KEYINPUT93), .B(n450), .Z(n451) );
  NAND2_X1 U510 ( .A1(n460), .A2(n451), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n452), .B(KEYINPUT94), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n453), .B(KEYINPUT25), .ZN(n457) );
  XNOR2_X1 U513 ( .A(KEYINPUT27), .B(n514), .ZN(n459) );
  NOR2_X1 U514 ( .A1(n473), .A2(n460), .ZN(n455) );
  INV_X1 U515 ( .A(n563), .ZN(n541) );
  NOR2_X1 U516 ( .A1(n459), .A2(n541), .ZN(n456) );
  NOR2_X1 U517 ( .A1(n457), .A2(n456), .ZN(n458) );
  NOR2_X1 U518 ( .A1(n458), .A2(n469), .ZN(n462) );
  NOR2_X1 U519 ( .A1(n512), .A2(n459), .ZN(n538) );
  XOR2_X1 U520 ( .A(KEYINPUT28), .B(n460), .Z(n498) );
  INV_X1 U521 ( .A(n498), .ZN(n519) );
  NAND2_X1 U522 ( .A1(n538), .A2(n519), .ZN(n523) );
  NOR2_X1 U523 ( .A1(n473), .A2(n523), .ZN(n461) );
  NOR2_X1 U524 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U525 ( .A(KEYINPUT95), .B(n463), .ZN(n481) );
  NAND2_X1 U526 ( .A1(n576), .A2(n481), .ZN(n464) );
  NOR2_X1 U527 ( .A1(n582), .A2(n464), .ZN(n466) );
  XNOR2_X1 U528 ( .A(KEYINPUT37), .B(KEYINPUT101), .ZN(n465) );
  XNOR2_X1 U529 ( .A(n466), .B(n465), .ZN(n511) );
  NAND2_X1 U530 ( .A1(n482), .A2(n511), .ZN(n467) );
  XNOR2_X1 U531 ( .A(n468), .B(n467), .ZN(n497) );
  NAND2_X1 U532 ( .A1(n497), .A2(n469), .ZN(n472) );
  XOR2_X1 U533 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n470) );
  XNOR2_X1 U534 ( .A(n470), .B(G29GAT), .ZN(n471) );
  XNOR2_X1 U535 ( .A(n472), .B(n471), .ZN(G1328GAT) );
  NAND2_X1 U536 ( .A1(n497), .A2(n473), .ZN(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n475) );
  XNOR2_X1 U538 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n474) );
  NAND2_X1 U539 ( .A1(n548), .A2(n478), .ZN(n479) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(n479), .Z(n480) );
  AND2_X1 U541 ( .A1(n481), .A2(n480), .ZN(n500) );
  NAND2_X1 U542 ( .A1(n482), .A2(n500), .ZN(n491) );
  NOR2_X1 U543 ( .A1(n512), .A2(n491), .ZN(n484) );
  XNOR2_X1 U544 ( .A(KEYINPUT34), .B(KEYINPUT96), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U546 ( .A(G1GAT), .B(n485), .Z(G1324GAT) );
  NOR2_X1 U547 ( .A1(n514), .A2(n491), .ZN(n487) );
  XNOR2_X1 U548 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U550 ( .A1(n524), .A2(n491), .ZN(n489) );
  XNOR2_X1 U551 ( .A(KEYINPUT35), .B(KEYINPUT98), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U553 ( .A(G15GAT), .B(n490), .ZN(G1326GAT) );
  NOR2_X1 U554 ( .A1(n519), .A2(n491), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(G1327GAT) );
  XOR2_X1 U557 ( .A(G36GAT), .B(KEYINPUT103), .Z(n496) );
  NAND2_X1 U558 ( .A1(n497), .A2(n494), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1329GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U562 ( .A(n544), .ZN(n558) );
  NOR2_X1 U563 ( .A1(n542), .A2(n558), .ZN(n510) );
  NAND2_X1 U564 ( .A1(n510), .A2(n500), .ZN(n506) );
  NOR2_X1 U565 ( .A1(n512), .A2(n506), .ZN(n502) );
  XNOR2_X1 U566 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n503), .Z(G1332GAT) );
  NOR2_X1 U569 ( .A1(n514), .A2(n506), .ZN(n504) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n524), .A2(n506), .ZN(n505) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n519), .A2(n506), .ZN(n508) );
  XNOR2_X1 U574 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U576 ( .A(G78GAT), .B(n509), .Z(G1335GAT) );
  NAND2_X1 U577 ( .A1(n511), .A2(n510), .ZN(n518) );
  NOR2_X1 U578 ( .A1(n512), .A2(n518), .ZN(n513) );
  XOR2_X1 U579 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U580 ( .A1(n514), .A2(n518), .ZN(n515) );
  XOR2_X1 U581 ( .A(KEYINPUT108), .B(n515), .Z(n516) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(n516), .ZN(G1337GAT) );
  NOR2_X1 U583 ( .A1(n524), .A2(n518), .ZN(n517) );
  XOR2_X1 U584 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  NOR2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n521) );
  XNOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U590 ( .A1(n525), .A2(n539), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n526), .B(KEYINPUT111), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n534), .A2(n542), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(KEYINPUT112), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n530) );
  NAND2_X1 U596 ( .A1(n534), .A2(n544), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n532) );
  NAND2_X1 U599 ( .A1(n534), .A2(n548), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n536) );
  NAND2_X1 U603 ( .A1(n534), .A2(n551), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(n537), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n552), .A2(n542), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  NAND2_X1 U611 ( .A1(n552), .A2(n544), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(n547), .ZN(G1345GAT) );
  XOR2_X1 U614 ( .A(G155GAT), .B(KEYINPUT115), .Z(n550) );
  NAND2_X1 U615 ( .A1(n552), .A2(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U619 ( .A1(n565), .A2(n561), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(KEYINPUT117), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT118), .B(KEYINPUT57), .Z(n557) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n560) );
  NOR2_X1 U625 ( .A1(n558), .A2(n561), .ZN(n559) );
  XOR2_X1 U626 ( .A(n560), .B(n559), .Z(G1349GAT) );
  NOR2_X1 U627 ( .A1(n576), .A2(n561), .ZN(n562) );
  XOR2_X1 U628 ( .A(G183GAT), .B(n562), .Z(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n581) );
  NOR2_X1 U630 ( .A1(n565), .A2(n581), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT121), .Z(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT120), .B(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n581), .A2(n571), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT123), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n581), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT124), .B(n577), .Z(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n580) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(n584), .B(n583), .Z(G1355GAT) );
endmodule

