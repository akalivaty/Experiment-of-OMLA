//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(KEYINPUT22), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G148gat), .ZN(new_n212));
  INV_X1    g011(.A(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G141gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(KEYINPUT82), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT82), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT2), .B1(new_n212), .B2(new_n214), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(new_n219), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n211), .A2(G148gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(KEYINPUT83), .B2(new_n212), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n212), .A2(KEYINPUT83), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n219), .B1(new_n218), .B2(KEYINPUT2), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n210), .B1(new_n234), .B2(KEYINPUT29), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT85), .B1(G228gat), .B2(G233gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(new_n210), .B2(KEYINPUT29), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n236), .B1(new_n238), .B2(new_n233), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT31), .B(G22gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(KEYINPUT85), .A2(G228gat), .A3(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(G50gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n235), .A2(new_n239), .A3(new_n241), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n247), .B1(new_n243), .B2(new_n248), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n203), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n243), .A2(new_n248), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n246), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n202), .A3(new_n249), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT77), .ZN(new_n257));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n261));
  INV_X1    g060(.A(G169gat), .ZN(new_n262));
  INV_X1    g061(.A(G176gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT23), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n260), .A2(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(G169gat), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n263), .A2(KEYINPUT64), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n263), .A2(KEYINPUT64), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT24), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n273), .B(new_n274), .C1(G183gat), .C2(G190gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n266), .A2(new_n270), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT25), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n279), .B1(new_n273), .B2(KEYINPUT66), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n271), .A2(new_n281), .A3(new_n272), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n274), .A2(KEYINPUT67), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n274), .A2(KEYINPUT67), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n280), .A2(new_n282), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  AND3_X1   g084(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  OAI22_X1  g087(.A1(new_n286), .A2(new_n287), .B1(KEYINPUT23), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT25), .B1(new_n264), .B2(new_n265), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n278), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n271), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT69), .ZN(new_n295));
  AOI22_X1  g094(.A1(KEYINPUT26), .A2(new_n295), .B1(new_n260), .B2(new_n261), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT26), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n288), .A2(KEYINPUT69), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n294), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G190gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(KEYINPUT68), .B2(KEYINPUT28), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n306));
  OAI22_X1  g105(.A1(new_n302), .A2(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT27), .B(G183gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n305), .A2(new_n306), .ZN(new_n309));
  AOI21_X1  g108(.A(G190gat), .B1(new_n305), .B2(new_n306), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n299), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n299), .B2(new_n312), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n293), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OR2_X1    g115(.A1(G127gat), .A2(G134gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(G127gat), .A2(G134gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(G113gat), .B2(G120gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT71), .B(G113gat), .ZN(new_n323));
  INV_X1    g122(.A(G120gat), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n319), .B(new_n322), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G113gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(new_n324), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n317), .B(new_n318), .C1(new_n327), .C2(new_n321), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT72), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n325), .A2(new_n331), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n332), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n331), .B1(new_n325), .B2(new_n328), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n337), .B(new_n293), .C1(new_n315), .C2(new_n314), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G227gat), .ZN(new_n340));
  INV_X1    g139(.A(G233gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT34), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT73), .B1(new_n339), .B2(new_n342), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n347));
  INV_X1    g146(.A(new_n342), .ZN(new_n348));
  AOI211_X1 g147(.A(new_n347), .B(new_n348), .C1(new_n334), .C2(new_n338), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT32), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT33), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(new_n346), .B2(new_n349), .ZN(new_n352));
  XOR2_X1   g151(.A(G15gat), .B(G43gat), .Z(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT76), .ZN(new_n354));
  XOR2_X1   g153(.A(G71gat), .B(G99gat), .Z(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n350), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  OAI221_X1 g159(.A(KEYINPUT32), .B1(new_n351), .B2(new_n358), .C1(new_n346), .C2(new_n349), .ZN(new_n361));
  AOI211_X1 g160(.A(new_n257), .B(new_n345), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n345), .A3(new_n361), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n257), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n256), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367));
  INV_X1    g166(.A(G85gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT0), .B(G57gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n329), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n221), .A2(new_n225), .B1(new_n230), .B2(new_n231), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(new_n237), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n333), .B2(new_n233), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n373), .A2(KEYINPUT4), .A3(new_n372), .ZN(new_n379));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(KEYINPUT5), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n376), .A2(new_n378), .A3(new_n379), .A4(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n373), .A2(new_n330), .A3(KEYINPUT4), .A4(new_n332), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n380), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n329), .B1(new_n233), .B2(KEYINPUT3), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n373), .A2(new_n237), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT4), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n372), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n233), .A2(new_n329), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n389), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n391), .B1(new_n393), .B2(new_n381), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n371), .B(new_n383), .C1(new_n390), .C2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n399));
  INV_X1    g198(.A(new_n371), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n383), .B1(new_n390), .B2(new_n395), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n398), .A2(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n396), .A2(KEYINPUT84), .A3(new_n397), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n400), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT81), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n278), .A2(new_n292), .B1(new_n299), .B2(new_n312), .ZN(new_n411));
  NAND2_X1  g210(.A1(G226gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n277), .A2(new_n276), .B1(new_n285), .B2(new_n291), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n309), .B1(new_n308), .B2(new_n310), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n295), .A2(KEYINPUT26), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n260), .A2(new_n261), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(new_n298), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n271), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT70), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n299), .A2(new_n312), .A3(new_n313), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n415), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n413), .A2(KEYINPUT29), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n210), .B(new_n414), .C1(new_n425), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT78), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n316), .A2(new_n426), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT78), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n430), .A2(new_n431), .A3(new_n210), .A4(new_n414), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n412), .B1(new_n411), .B2(KEYINPUT29), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT79), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n316), .A2(new_n413), .ZN(new_n436));
  INV_X1    g235(.A(new_n210), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n438), .B(new_n412), .C1(new_n411), .C2(KEYINPUT29), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n435), .A2(new_n436), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n433), .A2(KEYINPUT80), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT80), .B1(new_n433), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n410), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n433), .A2(new_n440), .A3(new_n409), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n433), .A2(KEYINPUT30), .A3(new_n440), .A4(new_n409), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n406), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT35), .B1(new_n366), .B2(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n252), .A2(new_n255), .ZN(new_n452));
  INV_X1    g251(.A(new_n383), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n377), .B1(new_n374), .B2(new_n375), .ZN(new_n454));
  INV_X1    g253(.A(new_n389), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n380), .B(new_n384), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n456), .B2(new_n394), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n371), .B(KEYINPUT87), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n396), .B(new_n397), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n459), .A2(new_n405), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n452), .A2(new_n460), .A3(KEYINPUT35), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n360), .A2(new_n361), .ZN(new_n462));
  INV_X1    g261(.A(new_n345), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n363), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n461), .B(new_n449), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT36), .B1(new_n362), .B2(new_n365), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT36), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n464), .A2(new_n470), .A3(new_n363), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT40), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT39), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n381), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n458), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT39), .B1(new_n393), .B2(new_n381), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n381), .B2(new_n475), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n474), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n458), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n401), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n475), .A2(new_n381), .ZN(new_n484));
  INV_X1    g283(.A(new_n479), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n486), .A2(KEYINPUT40), .A3(new_n458), .A4(new_n477), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n481), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n410), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n316), .A2(new_n426), .B1(new_n413), .B2(new_n411), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n431), .B1(new_n490), .B2(new_n210), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n428), .A2(KEYINPUT78), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n440), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT80), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n433), .A2(KEYINPUT80), .A3(new_n440), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n489), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n446), .A2(new_n447), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n488), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n256), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n433), .A2(new_n501), .A3(new_n440), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT38), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n410), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n490), .B2(new_n437), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n435), .A2(new_n436), .A3(new_n210), .A4(new_n439), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n459), .A2(new_n508), .A3(new_n405), .A4(new_n444), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT37), .B1(new_n441), .B2(new_n442), .ZN(new_n510));
  INV_X1    g309(.A(new_n409), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n509), .B1(new_n514), .B2(KEYINPUT38), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n473), .B1(new_n500), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n256), .B(KEYINPUT86), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n450), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n452), .B1(new_n448), .B2(new_n488), .ZN(new_n519));
  AND4_X1   g318(.A1(new_n405), .A2(new_n459), .A3(new_n508), .A4(new_n444), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n495), .A2(new_n496), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n512), .B1(new_n521), .B2(KEYINPUT37), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n522), .B2(new_n503), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(new_n523), .A3(KEYINPUT88), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n472), .A2(new_n516), .A3(new_n518), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n468), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT16), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(G1gat), .B1(new_n527), .B2(KEYINPUT91), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G8gat), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(G57gat), .A2(G64gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(G57gat), .A2(G64gat), .ZN(new_n539));
  AND2_X1   g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n538), .B(new_n539), .C1(new_n540), .C2(KEYINPUT9), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(KEYINPUT94), .B2(new_n540), .ZN(new_n542));
  NOR2_X1   g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n542), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT95), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT21), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n545), .A2(KEYINPUT21), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n537), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550));
  INV_X1    g349(.A(G183gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(new_n205), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n548), .A2(new_n537), .ZN(new_n554));
  OR3_X1    g353(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n549), .B2(new_n554), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G127gat), .B(G155gat), .Z(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n558), .B(new_n559), .Z(new_n560));
  OR2_X1    g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n555), .A2(new_n560), .A3(new_n556), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G134gat), .B(G162gat), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT14), .ZN(new_n568));
  INV_X1    g367(.A(G29gat), .ZN(new_n569));
  INV_X1    g368(.A(G36gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n571), .A2(new_n572), .B1(G29gat), .B2(G36gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(G43gat), .B(G50gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT90), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(new_n573), .A3(new_n575), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  INV_X1    g381(.A(G92gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(KEYINPUT8), .A2(new_n582), .B1(new_n368), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT7), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(new_n368), .B2(new_n583), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G99gat), .B(G106gat), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n588), .B(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT17), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n567), .B1(new_n581), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n580), .ZN(new_n594));
  NOR3_X1   g393(.A1(new_n594), .A2(KEYINPUT17), .A3(new_n591), .ZN(new_n595));
  XOR2_X1   g394(.A(G190gat), .B(G218gat), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OR3_X1    g396(.A1(new_n593), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n593), .B2(new_n595), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n566), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n598), .A2(new_n566), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n599), .A2(KEYINPUT96), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT97), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n601), .A2(new_n602), .A3(new_n606), .A4(new_n603), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n600), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n563), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT98), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT98), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n563), .A2(new_n611), .A3(new_n608), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n526), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT17), .ZN(new_n617));
  INV_X1    g416(.A(new_n537), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n617), .B1(new_n618), .B2(KEYINPUT92), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n581), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n581), .A2(KEYINPUT17), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n618), .B1(new_n621), .B2(KEYINPUT92), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n616), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  OR3_X1    g422(.A1(new_n623), .A2(KEYINPUT93), .A3(KEYINPUT18), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n537), .B(new_n594), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n615), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT18), .B1(new_n623), .B2(KEYINPUT93), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(G113gat), .B(G141gat), .Z(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT89), .B(G197gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT11), .B(G169gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT12), .Z(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n636), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n624), .A2(new_n638), .A3(new_n628), .A4(new_n629), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(G230gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n341), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n546), .A2(KEYINPUT10), .A3(new_n591), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n545), .B1(new_n645), .B2(new_n590), .ZN(new_n646));
  INV_X1    g445(.A(new_n591), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n545), .B(new_n591), .C1(new_n645), .C2(new_n590), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n643), .B1(new_n644), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n643), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n648), .B2(new_n649), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT100), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n655), .A2(KEYINPUT100), .A3(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n641), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n614), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n406), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT101), .B(G1gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1324gat));
  INV_X1    g467(.A(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n448), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT42), .B1(new_n671), .B2(new_n534), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  MUX2_X1   g473(.A(KEYINPUT42), .B(new_n672), .S(new_n674), .Z(G1325gat));
  INV_X1    g474(.A(new_n472), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n669), .A2(new_n676), .A3(G15gat), .ZN(new_n677));
  INV_X1    g476(.A(G15gat), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n465), .A2(new_n466), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n665), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n681), .B2(new_n680), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n669), .A2(new_n517), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT103), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  NOR3_X1   g486(.A1(new_n500), .A2(new_n515), .A3(new_n473), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT88), .B1(new_n519), .B2(new_n523), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n469), .A2(new_n471), .B1(new_n450), .B2(new_n517), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n690), .A2(new_n691), .B1(new_n451), .B2(new_n467), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(new_n608), .A3(new_n563), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n664), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G29gat), .A3(new_n406), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n563), .B(KEYINPUT104), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n664), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT105), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n692), .B2(new_n608), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n608), .A2(KEYINPUT106), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n705));
  AOI211_X1 g504(.A(new_n705), .B(new_n600), .C1(new_n605), .C2(new_n607), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n526), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n701), .B1(new_n702), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n703), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n468), .B2(new_n525), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(KEYINPUT107), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n700), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n406), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n569), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n696), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1328gat));
  OAI21_X1  g518(.A(G36gat), .B1(new_n713), .B2(new_n449), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n693), .A2(new_n570), .A3(new_n664), .A4(new_n448), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n721), .A2(new_n722), .A3(KEYINPUT46), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(KEYINPUT46), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n721), .B2(KEYINPUT46), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n720), .A2(new_n723), .A3(new_n724), .A4(new_n725), .ZN(G1329gat));
  NOR3_X1   g525(.A1(new_n694), .A2(G43gat), .A3(new_n679), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n714), .A2(new_n676), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(G43gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g529(.A(G50gat), .B1(new_n713), .B2(new_n256), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n517), .A2(new_n245), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n694), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(KEYINPUT48), .A3(new_n734), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n517), .B(new_n700), .C1(new_n709), .C2(new_n712), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G50gat), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n736), .A2(KEYINPUT110), .A3(G50gat), .ZN(new_n740));
  AOI211_X1 g539(.A(KEYINPUT111), .B(KEYINPUT48), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742));
  INV_X1    g541(.A(new_n517), .ZN(new_n743));
  INV_X1    g542(.A(new_n608), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n703), .B1(new_n526), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT107), .B1(new_n745), .B2(new_n711), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n708), .A2(new_n701), .ZN(new_n747));
  AOI211_X1 g546(.A(new_n743), .B(new_n699), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n738), .B1(new_n748), .B2(new_n245), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n740), .A3(new_n734), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n742), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n735), .B1(new_n741), .B2(new_n752), .ZN(G1331gat));
  INV_X1    g552(.A(new_n663), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n640), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n614), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n715), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g558(.A1(new_n756), .A2(new_n449), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  AND2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n760), .B2(new_n761), .ZN(G1333gat));
  OAI21_X1  g563(.A(G71gat), .B1(new_n756), .B2(new_n472), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n679), .A2(G71gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n756), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g567(.A1(new_n757), .A2(new_n517), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g569(.A1(new_n693), .A2(new_n641), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT51), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n693), .A2(new_n773), .A3(new_n641), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n663), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n715), .ZN(new_n777));
  INV_X1    g576(.A(new_n563), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n755), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n746), .B2(new_n747), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n406), .A2(new_n368), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(G1336gat));
  NAND2_X1  g581(.A1(new_n448), .A2(new_n583), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n775), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n583), .B1(new_n780), .B2(new_n448), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n785), .B2(KEYINPUT112), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n786), .B(new_n788), .Z(G1337gat));
  OR2_X1    g588(.A1(new_n775), .A2(new_n679), .ZN(new_n790));
  INV_X1    g589(.A(G99gat), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n472), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n790), .A2(new_n791), .B1(new_n780), .B2(new_n792), .ZN(G1338gat));
  INV_X1    g592(.A(G106gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n776), .A2(new_n794), .A3(new_n452), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n517), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G106gat), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n794), .B1(new_n780), .B2(new_n452), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n795), .A2(new_n799), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n798), .A2(new_n799), .B1(new_n800), .B2(new_n801), .ZN(G1339gat));
  INV_X1    g601(.A(new_n697), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n644), .A2(new_n651), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n653), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n805), .A2(new_n806), .A3(new_n652), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n660), .B1(new_n652), .B2(new_n806), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(KEYINPUT55), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  INV_X1    g610(.A(new_n809), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n655), .A2(new_n659), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n810), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n637), .B2(new_n639), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817));
  OR3_X1    g616(.A1(new_n625), .A2(new_n817), .A3(new_n627), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n620), .A2(new_n616), .A3(new_n622), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n625), .B2(new_n627), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n635), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(KEYINPUT114), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(KEYINPUT114), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n823), .A2(new_n639), .A3(new_n663), .A4(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT115), .B1(new_n816), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n828), .B(new_n825), .C1(new_n641), .C2(new_n815), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n704), .A2(new_n706), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n823), .A2(new_n639), .A3(new_n824), .ZN(new_n832));
  INV_X1    g631(.A(new_n815), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n803), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n640), .A2(new_n663), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n610), .A2(new_n612), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n366), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n406), .A2(new_n448), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n323), .A3(new_n640), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n840), .A2(new_n679), .A3(new_n517), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n842), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(KEYINPUT116), .A3(new_n842), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n851), .A2(new_n640), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n845), .B1(new_n852), .B2(new_n326), .ZN(G1340gat));
  NAND3_X1  g652(.A1(new_n844), .A2(new_n324), .A3(new_n663), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n851), .A2(new_n663), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n324), .ZN(G1341gat));
  NAND2_X1  g655(.A1(new_n844), .A2(new_n563), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(KEYINPUT117), .ZN(new_n858));
  AOI21_X1  g657(.A(G127gat), .B1(new_n857), .B2(KEYINPUT117), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n803), .A2(G127gat), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n858), .A2(new_n859), .B1(new_n851), .B2(new_n860), .ZN(G1342gat));
  NAND2_X1  g660(.A1(new_n744), .A2(new_n449), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(G134gat), .A3(new_n406), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n841), .A2(new_n863), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT118), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(KEYINPUT118), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n849), .A2(new_n744), .A3(new_n850), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G134gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n865), .A2(KEYINPUT56), .A3(new_n866), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(G1343gat));
  NAND2_X1  g672(.A1(new_n472), .A2(new_n842), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n815), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n810), .A2(KEYINPUT119), .A3(new_n813), .A4(new_n814), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n640), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n744), .B1(new_n878), .B2(new_n825), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n778), .B1(new_n879), .B2(new_n835), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT120), .ZN(new_n881));
  INV_X1    g680(.A(new_n839), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n883), .B(new_n778), .C1(new_n879), .C2(new_n835), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n743), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n452), .B1(new_n837), .B2(new_n839), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n888), .A2(new_n889), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n887), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n839), .B1(new_n880), .B2(KEYINPUT120), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n884), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT121), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n874), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n211), .B1(new_n896), .B2(new_n640), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n676), .A2(new_n256), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n406), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI221_X1 g700(.A(new_n901), .B1(new_n900), .B2(new_n899), .C1(new_n837), .C2(new_n839), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n448), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n211), .A3(new_n640), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT58), .B1(new_n897), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n874), .ZN(new_n907));
  INV_X1    g706(.A(new_n890), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n908), .A2(KEYINPUT57), .B1(new_n894), .B2(KEYINPUT121), .ZN(new_n909));
  INV_X1    g708(.A(new_n895), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G141gat), .B1(new_n911), .B2(new_n641), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n904), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n906), .A2(new_n914), .ZN(G1344gat));
  NAND3_X1  g714(.A1(new_n903), .A2(new_n213), .A3(new_n663), .ZN(new_n916));
  AOI211_X1 g715(.A(KEYINPUT59), .B(new_n213), .C1(new_n896), .C2(new_n663), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n839), .A2(KEYINPUT123), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n839), .A2(KEYINPUT123), .ZN(new_n920));
  INV_X1    g719(.A(new_n834), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n879), .B1(new_n744), .B2(new_n921), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n919), .B(new_n920), .C1(new_n563), .C2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n886), .A3(new_n517), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n890), .A2(KEYINPUT57), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n663), .A3(new_n907), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n918), .B1(new_n927), .B2(G148gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n916), .B1(new_n917), .B2(new_n928), .ZN(G1345gat));
  AOI21_X1  g728(.A(G155gat), .B1(new_n903), .B2(new_n563), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n803), .A2(G155gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n896), .B2(new_n931), .ZN(G1346gat));
  OAI21_X1  g731(.A(G162gat), .B1(new_n911), .B2(new_n830), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n862), .A2(G162gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n902), .B2(new_n934), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n715), .A2(new_n449), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n841), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n262), .A3(new_n640), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n846), .A2(new_n936), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n640), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT124), .B1(new_n942), .B2(G169gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n939), .B1(new_n944), .B2(new_n945), .ZN(G1348gat));
  AOI21_X1  g745(.A(G176gat), .B1(new_n938), .B2(new_n663), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n754), .A2(new_n268), .A3(new_n269), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n941), .B2(new_n948), .ZN(G1349gat));
  NAND3_X1  g748(.A1(new_n938), .A2(new_n563), .A3(new_n308), .ZN(new_n950));
  OAI21_X1  g749(.A(G183gat), .B1(new_n940), .B2(new_n697), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n938), .A2(new_n303), .A3(new_n707), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n941), .A2(new_n744), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n956), .A3(G190gat), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n956), .B1(new_n955), .B2(G190gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  AND2_X1   g759(.A1(new_n472), .A2(new_n936), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n908), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT125), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n641), .A2(G197gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(new_n965), .ZN(new_n967));
  OAI21_X1  g766(.A(KEYINPUT125), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(G197gat), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n924), .A2(new_n925), .A3(new_n961), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n971), .B1(new_n972), .B2(new_n640), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT126), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n972), .A2(new_n640), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n969), .B(new_n975), .C1(new_n976), .C2(new_n971), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n974), .A2(new_n977), .ZN(G1352gat));
  NOR3_X1   g777(.A1(new_n962), .A2(G204gat), .A3(new_n754), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT62), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n926), .A2(new_n663), .A3(new_n961), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(G204gat), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1353gat));
  NAND3_X1  g782(.A1(new_n963), .A2(new_n205), .A3(new_n563), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n972), .A2(KEYINPUT127), .A3(new_n563), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n924), .A2(new_n925), .A3(new_n563), .A4(new_n961), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n205), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n985), .A2(new_n988), .A3(KEYINPUT63), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n985), .B2(new_n988), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n984), .B1(new_n989), .B2(new_n990), .ZN(G1354gat));
  AOI21_X1  g790(.A(G218gat), .B1(new_n963), .B2(new_n707), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n608), .A2(new_n206), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n992), .B1(new_n972), .B2(new_n993), .ZN(G1355gat));
endmodule


