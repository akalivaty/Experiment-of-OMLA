//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT0), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(KEYINPUT0), .B2(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n198), .A2(KEYINPUT66), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n199), .B1(new_n191), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G131), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n207), .A2(new_n209), .A3(new_n213), .A4(new_n210), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n204), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n218));
  INV_X1    g032(.A(G113), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n220), .A2(new_n221), .B1(KEYINPUT2), .B2(G113), .ZN(new_n222));
  INV_X1    g036(.A(G116), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(G119), .ZN(new_n224));
  INV_X1    g038(.A(G119), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT69), .B1(new_n225), .B2(G116), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n223), .A3(G119), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n222), .A2(new_n229), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n189), .B(G146), .C1(new_n193), .C2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n193), .A2(new_n187), .A3(G143), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT67), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n233), .A2(new_n237), .A3(new_n234), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n188), .A3(new_n190), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n206), .A2(G137), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n208), .A2(G134), .ZN(new_n243));
  OAI21_X1  g057(.A(G131), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n214), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n216), .A2(new_n232), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n222), .B(new_n229), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n200), .B1(new_n198), .B2(KEYINPUT66), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n191), .A2(new_n202), .A3(new_n199), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n255), .A2(new_n197), .B1(new_n212), .B2(new_n214), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n235), .A2(KEYINPUT67), .B1(new_n198), .B2(new_n239), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n245), .B1(new_n257), .B2(new_n238), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n252), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n249), .B1(new_n259), .B2(new_n248), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n251), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT71), .B(G237), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(G210), .A3(new_n263), .ZN(new_n264));
  XOR2_X1   g078(.A(KEYINPUT26), .B(G101), .Z(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n248), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT70), .B1(new_n256), .B2(new_n258), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT64), .B1(new_n216), .B2(new_n247), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT30), .B(new_n273), .C1(new_n274), .C2(KEYINPUT70), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n256), .A2(new_n258), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n276), .B(new_n277), .C1(new_n278), .C2(KEYINPUT64), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n272), .B1(new_n280), .B2(new_n252), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT31), .B1(new_n281), .B2(new_n269), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n232), .B1(new_n275), .B2(new_n279), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  NOR4_X1   g098(.A1(new_n283), .A2(new_n284), .A3(new_n272), .A4(new_n268), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n271), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n287));
  NOR2_X1   g101(.A1(G472), .A2(G902), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n288), .B(KEYINPUT73), .Z(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n286), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n287), .B1(new_n286), .B2(new_n290), .ZN(new_n292));
  INV_X1    g106(.A(G472), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n259), .A2(new_n248), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT28), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT74), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n294), .A2(new_n297), .A3(KEYINPUT28), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n268), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n296), .A2(new_n250), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n268), .B1(new_n283), .B2(new_n272), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT29), .B1(new_n261), .B2(new_n269), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n293), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(KEYINPUT75), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT75), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n309), .B(new_n293), .C1(new_n303), .C2(new_n306), .ZN(new_n310));
  OAI22_X1  g124(.A1(new_n291), .A2(new_n292), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n193), .A2(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT76), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(new_n225), .B2(G128), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n313), .B(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G110), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT24), .B(G110), .Z(new_n318));
  XNOR2_X1  g132(.A(G119), .B(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G125), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT16), .ZN(new_n325));
  OR3_X1    g139(.A1(new_n323), .A2(KEYINPUT16), .A3(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT77), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n323), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(KEYINPUT77), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(G146), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n325), .B2(new_n326), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n334), .A2(new_n187), .A3(new_n330), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n317), .B(new_n320), .C1(new_n332), .C2(new_n335), .ZN(new_n336));
  OAI22_X1  g150(.A1(new_n316), .A2(G110), .B1(new_n319), .B2(new_n318), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n328), .A2(G146), .A3(new_n331), .ZN(new_n338));
  XNOR2_X1  g152(.A(G125), .B(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n187), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G137), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n343), .B(new_n344), .Z(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n336), .A2(new_n341), .A3(new_n345), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n302), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT25), .A4(new_n302), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G217), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(G234), .B2(new_n302), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT78), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n353), .A2(new_n358), .A3(new_n355), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n347), .A2(new_n348), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n355), .A2(G902), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT79), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n357), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT9), .B(G234), .ZN(new_n365));
  OAI21_X1  g179(.A(G221), .B1(new_n365), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G469), .ZN(new_n368));
  XNOR2_X1  g182(.A(G110), .B(G140), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n263), .A2(G227), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n240), .A2(KEYINPUT81), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n233), .A2(new_n234), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n198), .A2(new_n374), .A3(new_n239), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(new_n377), .B2(G107), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  INV_X1    g193(.A(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G104), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(G107), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n378), .A2(new_n381), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n377), .A2(G107), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n380), .A2(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(G101), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n376), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n378), .A2(new_n381), .A3(new_n383), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G101), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n395), .A3(G101), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n204), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n241), .A2(KEYINPUT10), .A3(new_n388), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n391), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n215), .ZN(new_n400));
  INV_X1    g214(.A(new_n215), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n391), .A2(new_n397), .A3(new_n401), .A4(new_n398), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n371), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n389), .B1(new_n241), .B2(new_n388), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n405), .A2(KEYINPUT12), .A3(new_n215), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT12), .B1(new_n405), .B2(new_n215), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n402), .A2(new_n371), .ZN(new_n409));
  OAI22_X1  g223(.A1(new_n403), .A2(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI211_X1 g224(.A(KEYINPUT83), .B(new_n371), .C1(new_n400), .C2(new_n402), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n368), .B(new_n302), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n368), .A2(new_n302), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n402), .B1(new_n406), .B2(new_n407), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n371), .B(KEYINPUT80), .Z(new_n415));
  INV_X1    g229(.A(new_n409), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n414), .A2(new_n415), .B1(new_n416), .B2(new_n400), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n413), .B1(new_n417), .B2(G469), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n367), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n189), .A2(G128), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n193), .A2(G143), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(new_n206), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n223), .A2(KEYINPUT14), .A3(G122), .ZN(new_n424));
  XNOR2_X1  g238(.A(G116), .B(G122), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(G107), .B(new_n424), .C1(new_n426), .C2(KEYINPUT14), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n423), .B(new_n427), .C1(G107), .C2(new_n426), .ZN(new_n428));
  INV_X1    g242(.A(new_n420), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n429), .A2(KEYINPUT13), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n421), .B1(new_n429), .B2(KEYINPUT13), .ZN(new_n431));
  OAI21_X1  g245(.A(G134), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n422), .A2(new_n206), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n425), .B(new_n380), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n365), .A2(new_n354), .A3(G953), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n428), .A2(new_n435), .A3(new_n437), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n302), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n441), .B2(new_n302), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(G475), .A2(G902), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n332), .A2(new_n335), .ZN(new_n450));
  AND2_X1   g264(.A1(KEYINPUT71), .A2(G237), .ZN(new_n451));
  NOR2_X1   g265(.A1(KEYINPUT71), .A2(G237), .ZN(new_n452));
  OAI211_X1 g266(.A(G214), .B(new_n263), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT86), .B(G143), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OR2_X1    g269(.A1(KEYINPUT86), .A2(G143), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n262), .A2(G214), .A3(new_n263), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G131), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT17), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(new_n457), .A3(new_n213), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n213), .B1(new_n455), .B2(new_n457), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT17), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n450), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G113), .B(G122), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(new_n377), .ZN(new_n467));
  NAND2_X1  g281(.A1(KEYINPUT18), .A2(G131), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n455), .A2(new_n457), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n339), .B(new_n187), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n471));
  INV_X1    g285(.A(new_n468), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n458), .B2(new_n472), .ZN(new_n473));
  AOI211_X1 g287(.A(KEYINPUT87), .B(new_n468), .C1(new_n455), .C2(new_n457), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n469), .B(new_n470), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n465), .A2(new_n467), .A3(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n339), .B(KEYINPUT19), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n187), .ZN(new_n478));
  INV_X1    g292(.A(new_n461), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n478), .B(new_n338), .C1(new_n479), .C2(new_n463), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n467), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n449), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT20), .ZN(new_n483));
  INV_X1    g297(.A(new_n467), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n469), .A2(new_n470), .ZN(new_n485));
  INV_X1    g299(.A(new_n473), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n458), .A2(new_n471), .A3(new_n472), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n480), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n484), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n465), .A2(new_n467), .A3(new_n475), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n449), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n467), .B1(new_n465), .B2(new_n475), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n302), .B1(new_n476), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n483), .A2(new_n494), .B1(G475), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n419), .A2(new_n448), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G214), .B1(G237), .B2(G902), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n204), .A2(G125), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n241), .A2(new_n323), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n263), .A2(G224), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT84), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n226), .A2(new_n228), .ZN(new_n510));
  INV_X1    g324(.A(new_n224), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(KEYINPUT5), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT5), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n219), .B1(new_n224), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n222), .A2(new_n229), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n388), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n396), .B1(new_n230), .B2(new_n231), .ZN(new_n518));
  INV_X1    g332(.A(new_n394), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(G110), .B(G122), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n517), .B(new_n521), .C1(new_n518), .C2(new_n519), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n509), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n508), .B1(new_n520), .B2(new_n522), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n505), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n521), .B(KEYINPUT8), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n515), .A2(new_n388), .A3(new_n516), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n388), .B1(new_n515), .B2(new_n516), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n323), .B1(new_n255), .B2(new_n197), .ZN(new_n532));
  AOI21_X1  g346(.A(G125), .B1(new_n257), .B2(new_n238), .ZN(new_n533));
  OAI211_X1 g347(.A(KEYINPUT7), .B(new_n504), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n504), .A2(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n501), .A2(new_n502), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT85), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n531), .A2(new_n534), .A3(KEYINPUT85), .A4(new_n536), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n524), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n527), .A2(new_n541), .A3(new_n302), .ZN(new_n542));
  OAI21_X1  g356(.A(G210), .B1(G237), .B2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n527), .A2(new_n541), .A3(new_n302), .A4(new_n543), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n500), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(G234), .A2(G237), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(G952), .A3(new_n263), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(G902), .A3(G953), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT21), .B(G898), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n547), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n498), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n311), .A2(new_n364), .A3(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(G101), .ZN(G3));
  NAND2_X1  g373(.A1(new_n280), .A2(new_n252), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n248), .A3(new_n269), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n284), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n281), .A2(KEYINPUT31), .A3(new_n269), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n270), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(new_n289), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n293), .B1(new_n286), .B2(new_n302), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n357), .A2(new_n359), .A3(new_n363), .ZN(new_n568));
  INV_X1    g382(.A(new_n419), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n496), .A2(G475), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n493), .B1(new_n492), .B2(new_n449), .ZN(new_n573));
  INV_X1    g387(.A(new_n449), .ZN(new_n574));
  AOI211_X1 g388(.A(KEYINPUT20), .B(new_n574), .C1(new_n490), .C2(new_n491), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n572), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(KEYINPUT88), .A2(KEYINPUT33), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n441), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(KEYINPUT88), .A2(KEYINPUT33), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n439), .B(new_n440), .C1(new_n580), .C2(new_n577), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n579), .A2(G478), .A3(new_n581), .A4(new_n302), .ZN(new_n582));
  INV_X1    g396(.A(new_n441), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n442), .B1(new_n583), .B2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n576), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n556), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n571), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT34), .B(G104), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G6));
  INV_X1    g404(.A(KEYINPUT89), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n483), .A2(new_n494), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n446), .A2(new_n447), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n572), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n591), .B1(new_n594), .B2(new_n554), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n497), .A2(KEYINPUT89), .A3(new_n555), .A4(new_n593), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n595), .A2(new_n547), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n571), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT35), .B(G107), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G9));
  OR2_X1    g414(.A1(new_n346), .A2(KEYINPUT36), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n342), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n342), .A2(new_n601), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n362), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT90), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n357), .A3(new_n359), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n557), .A2(new_n567), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT37), .B(G110), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G12));
  INV_X1    g424(.A(KEYINPUT92), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n545), .A2(new_n546), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n499), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n549), .B(KEYINPUT91), .Z(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(G900), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(new_n552), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n497), .A2(new_n593), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n611), .B1(new_n613), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n594), .A2(new_n617), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(KEYINPUT92), .A3(new_n547), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n358), .B1(new_n353), .B2(new_n355), .ZN(new_n624));
  INV_X1    g438(.A(new_n355), .ZN(new_n625));
  AOI211_X1 g439(.A(KEYINPUT78), .B(new_n625), .C1(new_n351), .C2(new_n352), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n624), .A2(new_n626), .A3(new_n605), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n569), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n623), .A2(new_n311), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G128), .ZN(G30));
  XNOR2_X1  g444(.A(new_n612), .B(KEYINPUT38), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n497), .A2(new_n448), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(new_n499), .A3(new_n627), .A4(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n561), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n294), .A2(new_n268), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n635), .B(KEYINPUT93), .Z(new_n636));
  OAI21_X1  g450(.A(new_n302), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G472), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n638), .B1(new_n291), .B2(new_n292), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT94), .ZN(new_n641));
  OR3_X1    g455(.A1(new_n633), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n641), .B1(new_n633), .B2(new_n640), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n617), .B(KEYINPUT39), .Z(new_n644));
  NAND2_X1  g458(.A1(new_n419), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT95), .B(KEYINPUT40), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G143), .ZN(G45));
  NAND3_X1  g463(.A1(new_n576), .A2(new_n585), .A3(new_n618), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT96), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n576), .A2(new_n652), .A3(new_n585), .A4(new_n618), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n613), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n311), .A3(new_n628), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT97), .B(G146), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G48));
  OAI21_X1  g472(.A(new_n302), .B1(new_n410), .B2(new_n411), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(G469), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n366), .A3(new_n412), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n660), .A2(KEYINPUT98), .A3(new_n366), .A4(new_n412), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n311), .A2(new_n665), .A3(new_n364), .A4(new_n587), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT41), .B(G113), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G15));
  NAND4_X1  g482(.A1(new_n311), .A2(new_n665), .A3(new_n597), .A4(new_n364), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G116), .ZN(G18));
  AND3_X1   g484(.A1(new_n663), .A2(new_n547), .A3(new_n664), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n576), .A2(new_n593), .A3(new_n554), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n671), .A2(new_n311), .A3(new_n607), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G119), .ZN(G21));
  NAND2_X1  g488(.A1(new_n562), .A2(new_n563), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n298), .A2(new_n250), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n260), .A2(new_n297), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n268), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n289), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n566), .A2(new_n679), .A3(new_n568), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n547), .A2(new_n632), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n554), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n665), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G122), .ZN(G24));
  AND2_X1   g498(.A1(new_n651), .A2(new_n653), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n566), .A2(new_n679), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n686), .A3(new_n607), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n663), .A2(new_n547), .A3(new_n664), .ZN(new_n688));
  OAI21_X1  g502(.A(KEYINPUT99), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n566), .A2(new_n627), .A3(new_n679), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n671), .A2(new_n690), .A3(new_n691), .A4(new_n685), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT100), .B(G125), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G27));
  OAI21_X1  g509(.A(KEYINPUT32), .B1(new_n564), .B2(new_n289), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n286), .A2(new_n287), .A3(new_n290), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n301), .A2(new_n302), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n304), .B2(new_n305), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n309), .B1(new_n699), .B2(new_n293), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n307), .A2(KEYINPUT75), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n696), .A2(new_n697), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT102), .B1(new_n702), .B2(new_n568), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n311), .A2(new_n704), .A3(new_n364), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n412), .A2(new_n418), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n367), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n545), .A2(new_n499), .A3(new_n546), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n412), .A2(new_n418), .A3(KEYINPUT101), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n711), .A2(new_n654), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n703), .A2(new_n705), .A3(new_n713), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n311), .A2(new_n364), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n712), .B1(new_n716), .B2(new_n654), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G131), .ZN(G33));
  NAND4_X1  g533(.A1(new_n311), .A2(new_n364), .A3(new_n715), .A4(new_n621), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G134), .ZN(G36));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n576), .B(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n585), .A2(KEYINPUT43), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n497), .A2(new_n585), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  OAI22_X1  g541(.A1(new_n724), .A2(new_n725), .B1(KEYINPUT43), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n567), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n607), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT44), .A4(new_n607), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n417), .A2(KEYINPUT45), .ZN(new_n734));
  OAI21_X1  g548(.A(G469), .B1(new_n417), .B2(KEYINPUT45), .ZN(new_n735));
  OAI22_X1  g549(.A1(new_n734), .A2(new_n735), .B1(new_n368), .B2(new_n302), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT46), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n412), .A3(new_n739), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(new_n366), .A3(new_n644), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n732), .A2(new_n709), .A3(new_n733), .A4(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT104), .B(G137), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G39));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n366), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(KEYINPUT105), .B2(KEYINPUT47), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n545), .A2(new_n499), .A3(new_n546), .ZN(new_n747));
  NOR4_X1   g561(.A1(new_n311), .A2(new_n364), .A3(new_n654), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n740), .A2(new_n366), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n746), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(KEYINPUT106), .B(G140), .Z(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G42));
  NAND2_X1  g567(.A1(new_n660), .A2(new_n412), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n631), .B1(KEYINPUT49), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n585), .A2(new_n499), .A3(new_n366), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n724), .A2(new_n568), .A3(new_n756), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n754), .A2(KEYINPUT49), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n755), .A2(new_n640), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n754), .A2(new_n366), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n746), .B2(new_n750), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n728), .A2(new_n615), .A3(new_n680), .A4(new_n709), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT51), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n728), .A2(new_n615), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n663), .A2(new_n664), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n765), .A2(new_n766), .A3(new_n747), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n690), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n568), .A2(new_n549), .A3(new_n747), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n640), .A2(new_n665), .A3(new_n769), .ZN(new_n770));
  OR3_X1    g584(.A1(new_n770), .A2(new_n576), .A3(new_n585), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n768), .A2(new_n771), .A3(KEYINPUT112), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT112), .B1(new_n768), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(G472), .B1(new_n564), .B2(G902), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n675), .A2(new_n678), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n775), .B(new_n364), .C1(new_n289), .C2(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n765), .A2(new_n766), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n631), .A2(new_n499), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT50), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(KEYINPUT50), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n764), .B1(new_n774), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n782), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n785), .B(KEYINPUT113), .C1(new_n772), .C2(new_n773), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n763), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n767), .A2(new_n703), .A3(new_n705), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT48), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n778), .A2(new_n547), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT114), .Z(new_n791));
  OAI211_X1 g605(.A(G952), .B(new_n263), .C1(new_n770), .C2(new_n586), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n768), .B(new_n771), .C1(new_n761), .C2(new_n762), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n783), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n789), .B(new_n793), .C1(new_n795), .C2(KEYINPUT51), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n681), .A2(new_n607), .A3(new_n617), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n708), .A2(new_n710), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n639), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n629), .A2(new_n656), .A3(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n801), .A2(new_n693), .A3(KEYINPUT52), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(new_n801), .B2(new_n693), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n556), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT108), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n586), .B(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n567), .A2(new_n805), .A3(new_n570), .A4(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n558), .A2(KEYINPUT109), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT109), .B1(new_n558), .B2(new_n808), .ZN(new_n810));
  INV_X1    g624(.A(new_n594), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n567), .A2(new_n805), .A3(new_n570), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n608), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n809), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n576), .A2(new_n593), .A3(new_n617), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT110), .B1(new_n709), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n592), .A2(new_n448), .A3(new_n572), .A4(new_n618), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT110), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n747), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n311), .A3(new_n628), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n690), .A2(new_n685), .A3(new_n715), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n720), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n717), .B2(new_n714), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n669), .A2(new_n673), .A3(new_n666), .A4(new_n683), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT107), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n777), .A2(new_n766), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n607), .A2(new_n672), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n696), .A2(new_n697), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n700), .A2(new_n701), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n827), .A2(new_n682), .B1(new_n831), .B2(new_n671), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT107), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n666), .A4(new_n669), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n814), .A2(new_n824), .A3(new_n826), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n797), .B1(new_n804), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n810), .A2(new_n813), .ZN(new_n837));
  INV_X1    g651(.A(new_n809), .ZN(new_n838));
  INV_X1    g652(.A(new_n823), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n718), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n623), .A2(new_n311), .A3(new_n628), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n689), .B2(new_n692), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n656), .A2(new_n800), .A3(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n629), .A2(new_n656), .A3(new_n800), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n692), .B2(new_n689), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n846), .B2(KEYINPUT52), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n825), .A2(new_n797), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n840), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n814), .A2(new_n849), .A3(new_n824), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n801), .A2(new_n693), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n852), .A2(new_n853), .B1(new_n842), .B2(new_n843), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT111), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n836), .A2(new_n850), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT53), .B1(new_n804), .B2(new_n835), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n826), .A2(new_n834), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n840), .A2(new_n847), .A3(new_n859), .A4(new_n797), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(KEYINPUT54), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n787), .A2(new_n796), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(G952), .A2(G953), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n759), .B1(new_n863), .B2(new_n864), .ZN(G75));
  NOR2_X1   g679(.A1(new_n263), .A2(G952), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n836), .A2(new_n855), .A3(new_n850), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n868), .A2(G210), .A3(G902), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT56), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n525), .A2(new_n526), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(new_n505), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT55), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n867), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n874), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT115), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n871), .A2(new_n878), .A3(new_n874), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n875), .B1(new_n877), .B2(new_n879), .ZN(G51));
  NAND2_X1  g694(.A1(new_n868), .A2(KEYINPUT54), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n881), .A2(new_n857), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n413), .B(KEYINPUT57), .Z(new_n883));
  OAI22_X1  g697(.A1(new_n882), .A2(new_n883), .B1(new_n411), .B2(new_n410), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n734), .A2(new_n735), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n868), .A2(G902), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n886), .B(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n866), .B1(new_n884), .B2(new_n888), .ZN(G54));
  AND2_X1   g703(.A1(KEYINPUT58), .A2(G475), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n868), .A2(G902), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n892));
  INV_X1    g706(.A(new_n492), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n892), .B1(new_n891), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n867), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n868), .A2(G902), .A3(new_n492), .A4(new_n890), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT117), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(G60));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT59), .Z(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n857), .B2(new_n861), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n579), .A2(new_n581), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n881), .A2(new_n857), .ZN(new_n906));
  INV_X1    g720(.A(new_n904), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n902), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n905), .A2(new_n867), .A3(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n903), .A2(new_n900), .A3(new_n904), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(G63));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT120), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT60), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n868), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(new_n360), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n602), .A2(new_n603), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n868), .A2(new_n919), .A3(new_n915), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n920), .A2(new_n867), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n917), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n867), .B(new_n920), .C1(new_n916), .C2(new_n360), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n923), .A3(new_n922), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(G66));
  AOI21_X1  g743(.A(G953), .B1(new_n859), .B2(new_n814), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT122), .ZN(new_n931));
  INV_X1    g745(.A(G224), .ZN(new_n932));
  OAI21_X1  g746(.A(G953), .B1(new_n553), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(G898), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n872), .B1(new_n935), .B2(G953), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n934), .B(new_n936), .Z(G69));
  INV_X1    g751(.A(G227), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n938), .B2(new_n616), .ZN(new_n939));
  INV_X1    g753(.A(new_n681), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n741), .A2(new_n703), .A3(new_n940), .A4(new_n705), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n742), .A2(new_n751), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n842), .A2(new_n656), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT125), .B1(new_n718), .B2(new_n720), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n718), .A2(KEYINPUT125), .A3(new_n720), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n944), .B(new_n263), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n280), .B(new_n477), .Z(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(G900), .B2(G953), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n939), .B1(new_n951), .B2(KEYINPUT124), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n807), .A2(new_n811), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n953), .A2(new_n645), .A3(new_n747), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n364), .A3(new_n311), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n742), .A2(new_n751), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n648), .A2(new_n656), .A3(new_n842), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(KEYINPUT62), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n648), .A2(new_n959), .A3(new_n656), .A4(new_n842), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n958), .A2(KEYINPUT123), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT123), .B1(new_n958), .B2(new_n960), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n263), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n948), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n952), .A2(new_n964), .A3(new_n950), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n952), .B1(new_n964), .B2(new_n950), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(G72));
  NAND2_X1  g781(.A1(new_n859), .A2(new_n814), .ZN(new_n968));
  OR3_X1    g782(.A1(new_n961), .A2(new_n962), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT63), .Z(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT126), .ZN(new_n972));
  AOI211_X1 g786(.A(new_n268), .B(new_n281), .C1(new_n969), .C2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n972), .B1(new_n974), .B2(new_n968), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(new_n268), .A3(new_n281), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n634), .A2(KEYINPUT127), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(new_n304), .Z(new_n978));
  NAND4_X1  g792(.A1(new_n858), .A2(new_n860), .A3(new_n971), .A4(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n976), .A2(new_n867), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n973), .A2(new_n980), .ZN(G57));
endmodule


