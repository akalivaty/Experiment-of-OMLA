//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT0), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT0), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n189), .A2(new_n191), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT0), .A4(G128), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n200), .A2(KEYINPUT64), .A3(KEYINPUT0), .A4(G128), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n196), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  OR3_X1    g017(.A1(new_n202), .A2(KEYINPUT88), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n200), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n207));
  OAI21_X1  g021(.A(G128), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(G143), .B2(new_n188), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT68), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n205), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n200), .A2(new_n209), .A3(G128), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n203), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT88), .B1(new_n202), .B2(new_n203), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G224), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G953), .ZN(new_n218));
  XOR2_X1   g032(.A(new_n216), .B(new_n218), .Z(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT82), .B(G107), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n220), .A2(new_n222), .B1(new_n221), .B2(G107), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT3), .B1(new_n221), .B2(G107), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT81), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n226), .B(KEYINPUT3), .C1(new_n221), .C2(G107), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G101), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n223), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G107), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G104), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(new_n220), .B2(G104), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G101), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G116), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(G113), .B1(new_n238), .B2(KEYINPUT5), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT5), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n243), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n236), .A2(new_n247), .ZN(new_n248));
  XOR2_X1   g062(.A(G110), .B(G122), .Z(new_n249));
  INV_X1    g063(.A(new_n227), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n226), .B1(new_n232), .B2(KEYINPUT3), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT82), .A2(G107), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT82), .A2(G107), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n222), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n221), .A2(G107), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT83), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n223), .A2(new_n228), .A3(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n258), .A2(KEYINPUT84), .A3(G101), .A4(new_n260), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n258), .A2(G101), .A3(new_n260), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n230), .A2(KEYINPUT84), .ZN(new_n263));
  OAI211_X1 g077(.A(KEYINPUT4), .B(new_n261), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n241), .B(new_n242), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  AOI211_X1 g082(.A(new_n248), .B(new_n249), .C1(new_n264), .C2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n248), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n261), .A2(KEYINPUT4), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n256), .B(new_n255), .C1(new_n250), .C2(new_n251), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n229), .B1(new_n272), .B2(KEYINPUT83), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n273), .A2(new_n260), .B1(KEYINPUT84), .B2(new_n230), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n267), .A3(new_n260), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n265), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n270), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n249), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT87), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n269), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n278), .A2(KEYINPUT6), .A3(new_n281), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n219), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G210), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n214), .B1(new_n203), .B2(new_n202), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT7), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n218), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n235), .A2(new_n247), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n249), .B(KEYINPUT8), .Z(new_n296));
  NAND2_X1  g110(.A1(new_n244), .A2(KEYINPUT89), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n297), .A2(new_n246), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n244), .A2(KEYINPUT89), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n243), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n295), .B(new_n296), .C1(new_n235), .C2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n294), .B(new_n301), .C1(new_n216), .C2(new_n293), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n289), .B1(new_n269), .B2(new_n302), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n286), .A2(new_n288), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n248), .B1(new_n264), .B2(new_n268), .ZN(new_n305));
  INV_X1    g119(.A(new_n281), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n283), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n279), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n285), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n219), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n303), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n287), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n187), .B1(new_n304), .B2(new_n313), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT9), .B(G234), .Z(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G221), .B1(new_n316), .B2(G902), .ZN(new_n317));
  XNOR2_X1  g131(.A(G110), .B(G140), .ZN(new_n318));
  INV_X1    g132(.A(G953), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n319), .A2(G227), .ZN(new_n320));
  XOR2_X1   g134(.A(new_n318), .B(new_n320), .Z(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT85), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n276), .A2(new_n202), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n275), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G134), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT65), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT65), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G134), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G137), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT11), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(KEYINPUT11), .A3(G134), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT11), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G137), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n327), .A2(new_n329), .B1(KEYINPUT11), .B2(new_n331), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n337), .ZN(new_n341));
  OAI21_X1  g155(.A(G131), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n342), .A3(KEYINPUT69), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n276), .A2(new_n202), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n264), .A2(new_n348), .A3(KEYINPUT85), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n212), .A2(new_n213), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n236), .A2(KEYINPUT10), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n210), .A2(new_n192), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n213), .B1(new_n352), .B2(new_n200), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n230), .A2(new_n234), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n325), .A2(new_n347), .A3(new_n349), .A4(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n202), .B(new_n276), .C1(new_n271), .C2(new_n274), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n357), .B1(new_n361), .B2(new_n323), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n347), .B1(new_n362), .B2(new_n349), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n322), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n354), .B1(new_n236), .B2(new_n350), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT12), .A3(new_n343), .ZN(new_n366));
  INV_X1    g180(.A(new_n347), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n366), .B1(new_n368), .B2(KEYINPUT12), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n359), .A2(new_n321), .A3(new_n369), .ZN(new_n370));
  AOI211_X1 g184(.A(G469), .B(G902), .C1(new_n364), .C2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n325), .A2(new_n349), .A3(new_n358), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n367), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n359), .A3(new_n321), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n359), .A2(new_n369), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n322), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n376), .A3(G469), .ZN(new_n377));
  NAND2_X1  g191(.A1(G469), .A2(G902), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n317), .B1(new_n371), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT86), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(new_n317), .C1(new_n371), .C2(new_n379), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n314), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n345), .A2(new_n202), .A3(new_n346), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n334), .B1(G134), .B2(G137), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT65), .B(G134), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(new_n387), .B2(G137), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n350), .A2(new_n339), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n265), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n266), .A3(new_n389), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT28), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT28), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(G237), .A2(G953), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G210), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(new_n229), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(G902), .B1(new_n397), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT67), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n340), .A2(new_n341), .A3(G131), .ZN(new_n407));
  INV_X1    g221(.A(new_n386), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n330), .B2(new_n331), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n406), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n339), .A2(KEYINPUT67), .A3(new_n388), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n350), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT66), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n343), .A2(new_n413), .A3(new_n202), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n343), .B2(new_n202), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n265), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n392), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n418), .A2(KEYINPUT28), .B1(KEYINPUT72), .B2(new_n396), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT72), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n420), .B(new_n395), .C1(new_n417), .C2(new_n392), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n402), .B(KEYINPUT71), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n403), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT70), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n385), .A2(new_n426), .A3(KEYINPUT30), .A4(new_n389), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT70), .B1(new_n416), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n390), .A2(new_n428), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n265), .B(new_n427), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n392), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n402), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n405), .B1(new_n425), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G472), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n431), .A2(new_n392), .A3(new_n434), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT31), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n424), .B1(new_n419), .B2(new_n421), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT31), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n431), .A2(new_n441), .A3(new_n392), .A4(new_n434), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(G472), .A2(G902), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n443), .A2(KEYINPUT32), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT32), .B1(new_n443), .B2(new_n444), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT73), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n443), .A2(KEYINPUT32), .A3(new_n444), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT73), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n437), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n237), .A2(G128), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT23), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT75), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n237), .A2(G128), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT23), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n456), .A2(KEYINPUT76), .ZN(new_n457));
  OAI22_X1  g271(.A1(new_n456), .A2(KEYINPUT76), .B1(new_n237), .B2(G128), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n455), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(new_n452), .ZN(new_n461));
  XOR2_X1   g275(.A(KEYINPUT24), .B(G110), .Z(new_n462));
  OAI22_X1  g276(.A1(new_n459), .A2(G110), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G140), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n203), .A2(G140), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT16), .ZN(new_n467));
  OR3_X1    g281(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(G146), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n465), .A2(new_n466), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT78), .A3(new_n188), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT78), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n465), .A2(new_n466), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n472), .B1(new_n473), .B2(G146), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n463), .A2(new_n469), .A3(new_n475), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n459), .A2(G110), .B1(new_n461), .B2(new_n462), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT77), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n469), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(G146), .B1(new_n467), .B2(new_n468), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n478), .B(G146), .C1(new_n467), .C2(new_n468), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n319), .A2(G221), .A3(G234), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT79), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT22), .B(G137), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n476), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n488), .B1(new_n476), .B2(new_n484), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G217), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(G234), .B2(new_n289), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(G902), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n491), .ZN(new_n498));
  AOI21_X1  g312(.A(G902), .B1(new_n498), .B2(new_n489), .ZN(new_n499));
  OR2_X1    g313(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n500), .ZN(new_n502));
  NAND2_X1  g316(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n494), .B(KEYINPUT74), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n497), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT99), .ZN(new_n507));
  INV_X1    g321(.A(G478), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G122), .ZN(new_n511));
  OR3_X1    g325(.A1(new_n511), .A2(KEYINPUT14), .A3(G116), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT14), .B1(new_n511), .B2(G116), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n512), .B(new_n513), .C1(new_n239), .C2(G122), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G107), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT97), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(G116), .B(G122), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n220), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n190), .A2(G128), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n192), .A2(G143), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(new_n387), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n514), .A2(KEYINPUT97), .A3(G107), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n517), .A2(new_n519), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n522), .A2(new_n387), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n518), .A2(new_n220), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n527), .B2(new_n519), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT96), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT13), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT95), .B1(new_n520), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n520), .A2(new_n530), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n521), .A3(new_n532), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n520), .A2(KEYINPUT95), .A3(new_n530), .ZN(new_n534));
  OAI21_X1  g348(.A(G134), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n528), .A2(new_n529), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n529), .B1(new_n528), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n525), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n316), .A2(new_n493), .A3(G953), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n525), .B(new_n539), .C1(new_n536), .C2(new_n537), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n510), .B1(new_n543), .B2(new_n289), .ZN(new_n544));
  AOI211_X1 g358(.A(G902), .B(new_n509), .C1(new_n541), .C2(new_n542), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n398), .A2(G214), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n190), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n398), .A2(G143), .A3(G214), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(KEYINPUT18), .A2(G131), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT90), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n188), .B1(new_n465), .B2(new_n466), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n475), .B2(new_n555), .ZN(new_n556));
  AOI211_X1 g370(.A(KEYINPUT90), .B(new_n554), .C1(new_n471), .C2(new_n474), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n334), .B1(new_n548), .B2(new_n549), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT17), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n548), .A2(new_n334), .A3(new_n549), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(KEYINPUT17), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n563), .B(new_n564), .C1(new_n481), .C2(new_n482), .ZN(new_n565));
  XNOR2_X1  g379(.A(G113), .B(G122), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(new_n221), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n558), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n558), .B2(new_n565), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n289), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT94), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT94), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n573), .B(new_n289), .C1(new_n569), .C2(new_n570), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(G475), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT20), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT93), .ZN(new_n577));
  INV_X1    g391(.A(new_n551), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n550), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n475), .A2(new_n555), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT90), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n475), .A2(new_n553), .A3(new_n555), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n562), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n469), .B1(new_n584), .B2(new_n559), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n473), .B2(KEYINPUT92), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT19), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n586), .B(KEYINPUT19), .C1(new_n473), .C2(KEYINPUT92), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n470), .A2(KEYINPUT91), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n585), .B1(new_n593), .B2(new_n188), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n577), .B1(new_n583), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n567), .ZN(new_n596));
  OAI221_X1 g410(.A(new_n469), .B1(new_n559), .B2(new_n584), .C1(new_n592), .C2(G146), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n558), .A3(KEYINPUT93), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n568), .ZN(new_n600));
  NOR2_X1   g414(.A1(G475), .A2(G902), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n576), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n601), .ZN(new_n603));
  AOI211_X1 g417(.A(KEYINPUT20), .B(new_n603), .C1(new_n599), .C2(new_n568), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n546), .B(new_n575), .C1(new_n602), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(G234), .A2(G237), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n606), .A2(G952), .A3(new_n319), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(G902), .A3(G953), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n608), .B(KEYINPUT98), .Z(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT21), .B(G898), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n507), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n597), .A2(new_n558), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n567), .B1(new_n613), .B2(new_n577), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n569), .B1(new_n614), .B2(new_n598), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT20), .B1(new_n615), .B2(new_n603), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n600), .A2(new_n576), .A3(new_n601), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n574), .A2(G475), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n616), .A2(new_n617), .B1(new_n618), .B2(new_n572), .ZN(new_n619));
  INV_X1    g433(.A(new_n611), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(KEYINPUT99), .A3(new_n620), .A4(new_n546), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n612), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n384), .A2(new_n451), .A3(new_n506), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  NAND2_X1  g439(.A1(new_n443), .A2(new_n289), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(G472), .ZN(new_n628));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n443), .B(new_n289), .C1(KEYINPUT100), .C2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n506), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n381), .B2(new_n383), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n543), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n541), .A2(KEYINPUT33), .A3(new_n542), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(G478), .B1(new_n636), .B2(G902), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n543), .A2(new_n508), .A3(new_n289), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n638), .B1(new_n637), .B2(new_n639), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n619), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n620), .B(new_n187), .C1(new_n304), .C2(new_n313), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n632), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT34), .B(G104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  INV_X1    g463(.A(new_n546), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n619), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n632), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NAND2_X1  g469(.A1(new_n628), .A2(new_n630), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n504), .A2(new_n505), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n476), .A2(new_n484), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n488), .A2(KEYINPUT36), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n495), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n384), .A2(new_n623), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n607), .B1(new_n609), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n651), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n384), .A2(new_n451), .A3(new_n662), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  NAND2_X1  g486(.A1(new_n443), .A2(new_n444), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT32), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n449), .A3(new_n448), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n445), .A2(KEYINPUT73), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n438), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n424), .B2(new_n393), .ZN(new_n680));
  OAI21_X1  g494(.A(G472), .B1(new_n680), .B2(G902), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n304), .A2(new_n313), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT38), .Z(new_n684));
  INV_X1    g498(.A(new_n187), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n619), .A2(new_n546), .A3(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n682), .A2(new_n684), .A3(new_n663), .A4(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n381), .A2(new_n383), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n669), .B(KEYINPUT39), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT40), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n687), .A2(new_n688), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n689), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT103), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n689), .A2(new_n695), .A3(new_n699), .A4(new_n696), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n190), .ZN(G45));
  INV_X1    g516(.A(new_n669), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n643), .B(new_n703), .C1(new_n640), .C2(new_n641), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n384), .A2(new_n451), .A3(new_n662), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  AOI21_X1  g521(.A(new_n321), .B1(new_n373), .B2(new_n359), .ZN(new_n708));
  INV_X1    g522(.A(new_n370), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n289), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n364), .A2(new_n370), .ZN(new_n712));
  INV_X1    g526(.A(G469), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n289), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n711), .A2(new_n317), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n711), .A2(new_n714), .A3(KEYINPUT104), .A4(new_n317), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n451), .A2(new_n506), .A3(new_n646), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT105), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n720), .B(new_n722), .ZN(G15));
  NAND4_X1  g537(.A1(new_n451), .A2(new_n506), .A3(new_n652), .A4(new_n719), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NOR3_X1   g539(.A1(new_n622), .A2(new_n715), .A3(new_n314), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n451), .A2(new_n662), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  OAI21_X1  g542(.A(new_n288), .B1(new_n286), .B2(new_n303), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n311), .A2(new_n287), .A3(new_n312), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n685), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n619), .A2(new_n546), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n620), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n717), .B2(new_n718), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n439), .B(new_n442), .C1(new_n423), .C2(new_n397), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n444), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n626), .B2(G472), .ZN(new_n738));
  AOI211_X1 g552(.A(KEYINPUT106), .B(new_n629), .C1(new_n443), .C2(new_n289), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n506), .B(new_n736), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  OAI211_X1 g557(.A(new_n662), .B(new_n736), .C1(new_n738), .C2(new_n739), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n704), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n715), .A2(new_n314), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  NOR2_X1   g562(.A1(new_n445), .A2(new_n446), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n437), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n506), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n729), .A2(new_n187), .A3(new_n730), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n317), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n359), .A2(new_n321), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n756), .A2(new_n373), .B1(new_n375), .B2(new_n322), .ZN(new_n757));
  OAI21_X1  g571(.A(G469), .B1(new_n757), .B2(G902), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n755), .B1(new_n758), .B2(new_n714), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n729), .A2(new_n730), .A3(KEYINPUT107), .A4(new_n187), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n705), .A2(new_n754), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT42), .B1(new_n751), .B2(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n754), .A2(new_n759), .A3(new_n760), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n704), .A2(KEYINPUT42), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n451), .A2(new_n763), .A3(new_n506), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n334), .ZN(G33));
  NAND4_X1  g581(.A1(new_n451), .A2(new_n763), .A3(new_n506), .A4(new_n670), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  OR2_X1    g583(.A1(new_n757), .A2(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n757), .A2(KEYINPUT45), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(G469), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n378), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n714), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT46), .B1(new_n772), .B2(new_n378), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n317), .B(new_n692), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT108), .ZN(new_n777));
  INV_X1    g591(.A(new_n775), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n714), .A3(new_n773), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n780), .A3(new_n317), .A4(new_n692), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n754), .A2(new_n760), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n619), .B1(new_n640), .B2(new_n641), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n784), .A2(new_n785), .A3(KEYINPUT43), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n656), .A3(new_n662), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n783), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n792), .A2(KEYINPUT110), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n792), .A2(KEYINPUT110), .B1(new_n791), .B2(new_n790), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n782), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  NAND2_X1  g610(.A1(new_n779), .A2(new_n317), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT47), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n779), .A2(new_n799), .A3(new_n317), .ZN(new_n800));
  INV_X1    g614(.A(new_n783), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n801), .A2(new_n451), .A3(new_n506), .A4(new_n704), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n798), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  INV_X1    g618(.A(G952), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n319), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT117), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n684), .A2(new_n187), .A3(new_n715), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n788), .A2(new_n607), .A3(new_n789), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n740), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n812));
  OR3_X1    g626(.A1(new_n808), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n812), .B1(new_n808), .B2(new_n811), .ZN(new_n814));
  INV_X1    g628(.A(new_n744), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n809), .A2(new_n801), .A3(new_n715), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n813), .A2(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n715), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n783), .A2(new_n607), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n678), .A2(new_n506), .A3(new_n681), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n642), .A2(new_n643), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n711), .A2(new_n714), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n798), .A2(new_n800), .B1(new_n755), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n810), .A2(new_n783), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n817), .B(new_n825), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n644), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n822), .A2(new_n832), .A3(new_n823), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n805), .B(G953), .C1(new_n810), .C2(new_n746), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n816), .A2(new_n506), .A3(new_n750), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT48), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n834), .B1(new_n833), .B2(new_n835), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n839), .A2(KEYINPUT116), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT116), .B1(new_n839), .B2(new_n840), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n829), .A2(new_n830), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n831), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n671), .A2(new_n747), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n731), .A2(new_n732), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n847), .A2(new_n380), .A3(new_n669), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n682), .A2(new_n663), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n845), .A2(new_n846), .A3(new_n706), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(new_n645), .B2(new_n651), .ZN(new_n852));
  INV_X1    g666(.A(new_n651), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n731), .A2(KEYINPUT111), .A3(new_n620), .A4(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n632), .B1(new_n855), .B2(new_n646), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n624), .A3(new_n665), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n720), .A2(new_n724), .A3(new_n742), .A4(new_n727), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n671), .A2(new_n706), .A3(new_n747), .A4(new_n849), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT52), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n762), .A2(new_n765), .A3(new_n768), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n745), .A2(new_n763), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n605), .A2(new_n669), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n754), .A2(new_n760), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n451), .A2(new_n690), .A3(new_n865), .A4(new_n662), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n850), .A2(new_n859), .A3(new_n861), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT53), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n860), .B(new_n846), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n754), .A2(new_n760), .A3(new_n864), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n381), .B2(new_n383), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n663), .B1(new_n678), .B2(new_n437), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n873), .A2(new_n874), .B1(new_n745), .B2(new_n763), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n762), .A3(new_n765), .A4(new_n768), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n876), .A2(new_n857), .A3(new_n858), .ZN(new_n877));
  XNOR2_X1  g691(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n871), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n870), .A2(new_n880), .A3(KEYINPUT54), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n869), .A2(new_n879), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n768), .A2(KEYINPUT53), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n857), .A2(new_n766), .A3(new_n867), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n858), .A2(KEYINPUT113), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n874), .A2(new_n726), .B1(new_n741), .B2(new_n734), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT113), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n720), .A4(new_n724), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n884), .A2(new_n850), .A3(new_n861), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n882), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n807), .B1(new_n844), .B2(new_n893), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n826), .B(KEYINPUT49), .Z(new_n895));
  NAND4_X1  g709(.A1(new_n642), .A2(new_n619), .A3(new_n187), .A4(new_n317), .ZN(new_n896));
  OR3_X1    g710(.A1(new_n895), .A2(new_n684), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n894), .B1(new_n820), .B2(new_n897), .ZN(G75));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n289), .B1(new_n882), .B2(new_n890), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n900), .B2(G210), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n309), .B(new_n219), .ZN(new_n902));
  XNOR2_X1  g716(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n902), .B(new_n903), .Z(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n899), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(G210), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n907), .B(new_n289), .C1(new_n882), .C2(new_n890), .ZN(new_n908));
  OAI211_X1 g722(.A(KEYINPUT119), .B(new_n904), .C1(new_n908), .C2(KEYINPUT56), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n319), .A2(G952), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n904), .A2(KEYINPUT56), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n900), .A2(G210), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n908), .A2(KEYINPUT120), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n910), .A2(new_n917), .ZN(G51));
  XOR2_X1   g732(.A(new_n378), .B(KEYINPUT57), .Z(new_n919));
  INV_X1    g733(.A(new_n892), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n891), .B1(new_n882), .B2(new_n890), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n712), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n882), .A2(new_n890), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(G902), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n925), .A2(new_n772), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n911), .B1(new_n923), .B2(new_n926), .ZN(G54));
  INV_X1    g741(.A(new_n911), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT121), .B1(KEYINPUT58), .B2(G475), .ZN(new_n929));
  AND3_X1   g743(.A1(KEYINPUT121), .A2(KEYINPUT58), .A3(G475), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n925), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n928), .B1(new_n931), .B2(new_n600), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n600), .B2(new_n931), .ZN(G60));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT59), .Z(new_n935));
  NOR2_X1   g749(.A1(new_n636), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n920), .B2(new_n921), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n938), .A3(new_n928), .ZN(new_n939));
  INV_X1    g753(.A(new_n936), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n857), .A2(new_n867), .A3(new_n883), .ZN(new_n941));
  INV_X1    g755(.A(new_n766), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n889), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n850), .A2(new_n861), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n878), .B1(new_n871), .B2(new_n877), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT54), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n940), .B1(new_n947), .B2(new_n892), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT122), .B1(new_n948), .B2(new_n911), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n935), .B1(new_n881), .B2(new_n892), .ZN(new_n950));
  INV_X1    g764(.A(new_n636), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT123), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n935), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n893), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n955), .A3(new_n636), .ZN(new_n956));
  AND4_X1   g770(.A1(new_n939), .A2(new_n949), .A3(new_n952), .A4(new_n956), .ZN(G63));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT60), .Z(new_n959));
  NAND2_X1  g773(.A1(new_n924), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n492), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n924), .A2(new_n660), .A3(new_n959), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n928), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(G66));
  OAI21_X1  g779(.A(G953), .B1(new_n610), .B2(new_n217), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n859), .B2(G953), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n284), .B(new_n285), .C1(G898), .C2(new_n319), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G69));
  OAI21_X1  g783(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(new_n592), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n751), .A2(new_n847), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n862), .B1(new_n782), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n795), .A3(new_n803), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n671), .A2(new_n706), .A3(new_n747), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT124), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n319), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT125), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n668), .A2(G953), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n978), .B2(new_n980), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n971), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n832), .A2(new_n853), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n693), .A2(new_n984), .A3(new_n801), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n451), .A3(new_n506), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n795), .A2(new_n803), .A3(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n698), .A2(new_n700), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT62), .B1(new_n988), .B2(new_n976), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT62), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n701), .A2(new_n977), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n987), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n971), .A2(G953), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(G227), .A2(G900), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(G953), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n983), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n978), .A2(new_n980), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(KEYINPUT125), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1001), .A2(G953), .A3(new_n995), .A4(new_n971), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n997), .A2(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(new_n433), .A2(new_n402), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT126), .ZN(new_n1005));
  INV_X1    g819(.A(new_n859), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n974), .A2(new_n977), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1005), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n679), .A2(KEYINPUT127), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(new_n435), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n870), .A2(new_n880), .A3(new_n1009), .A4(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1011), .A2(new_n928), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1009), .B1(new_n992), .B2(new_n1006), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n433), .A2(new_n402), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(G57));
endmodule


