//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G227), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT78), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT12), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT64), .A2(G143), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT64), .A2(G143), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n193), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT66), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n193), .A2(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n196), .A2(new_n198), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT3), .A3(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT79), .B(G101), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n210), .A2(G104), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT83), .B1(new_n210), .B2(G104), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT82), .B1(new_n208), .B2(G107), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n208), .A3(G107), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT82), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(new_n210), .A3(G104), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n217), .A2(new_n218), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G101), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n206), .B1(new_n216), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT64), .ZN(new_n226));
  INV_X1    g040(.A(G143), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT64), .A2(G143), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(G146), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n204), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n230), .A2(new_n234), .A3(new_n204), .A4(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n225), .A2(KEYINPUT86), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT86), .B1(new_n225), .B2(new_n236), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n224), .A2(new_n216), .ZN(new_n239));
  AOI21_X1  g053(.A(G146), .B1(new_n228), .B2(new_n229), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n241));
  OAI21_X1  g055(.A(G128), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n230), .A2(new_n204), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n239), .B1(new_n236), .B2(new_n244), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n237), .A2(new_n238), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(G137), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT11), .A3(G134), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G131), .ZN(new_n254));
  INV_X1    g068(.A(G131), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n249), .A2(new_n251), .A3(new_n255), .A4(new_n252), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT85), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n192), .B1(new_n246), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n225), .A2(new_n236), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT86), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n204), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n194), .A2(new_n195), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(G146), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n234), .B1(new_n266), .B2(new_n231), .ZN(new_n267));
  INV_X1    g081(.A(new_n235), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n244), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n214), .B1(new_n209), .B2(new_n211), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n223), .A2(G101), .B1(new_n270), .B2(new_n213), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n225), .A2(KEYINPUT86), .A3(new_n236), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n263), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n259), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(KEYINPUT12), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n260), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n206), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(new_n267), .B2(new_n268), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT84), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n224), .A2(KEYINPUT10), .A3(new_n216), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n206), .B1(new_n233), .B2(new_n235), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT84), .B1(new_n284), .B2(new_n281), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT10), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n283), .A2(new_n285), .B1(new_n272), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G101), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(new_n212), .B2(new_n215), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT4), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT80), .ZN(new_n292));
  NOR4_X1   g106(.A1(new_n270), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n288), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n296));
  AND2_X1   g110(.A1(KEYINPUT0), .A2(G128), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n230), .A2(new_n204), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT0), .B(G128), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(new_n196), .B2(new_n198), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n216), .B(KEYINPUT4), .C1(new_n288), .C2(new_n270), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n295), .A2(new_n296), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT80), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n289), .B2(new_n290), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n301), .B(new_n302), .C1(new_n305), .C2(new_n293), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT81), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n254), .A2(new_n256), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n287), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n191), .B1(new_n277), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n306), .B(new_n296), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n233), .A2(new_n235), .B1(new_n242), .B2(new_n243), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n286), .B1(new_n313), .B2(new_n239), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n280), .B1(new_n279), .B2(new_n282), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n284), .A2(KEYINPUT84), .A3(new_n281), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n257), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n318), .A2(new_n191), .A3(new_n310), .ZN(new_n319));
  INV_X1    g133(.A(G469), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n311), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G902), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT87), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n274), .A2(KEYINPUT12), .A3(new_n275), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT12), .B1(new_n274), .B2(new_n275), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n310), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n191), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n320), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n318), .A2(new_n191), .A3(new_n310), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT87), .ZN(new_n332));
  INV_X1    g146(.A(new_n323), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n287), .A2(new_n308), .A3(new_n309), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n309), .B1(new_n287), .B2(new_n308), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n328), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n191), .B(new_n310), .C1(new_n325), .C2(new_n326), .ZN(new_n338));
  AOI21_X1  g152(.A(G902), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n320), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n324), .A2(new_n334), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G221), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT9), .B(G234), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n342), .B1(new_n344), .B2(new_n322), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT77), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G237), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n187), .A3(G214), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n228), .A3(new_n229), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n348), .A2(new_n187), .A3(G143), .A4(G214), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G131), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT17), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n255), .A3(new_n351), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G140), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT16), .B1(new_n357), .B2(G125), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT75), .ZN(new_n359));
  INV_X1    g173(.A(G125), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n359), .B1(new_n360), .B2(G140), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(KEYINPUT75), .A3(G125), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(G140), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI211_X1 g178(.A(G146), .B(new_n358), .C1(new_n364), .C2(KEYINPUT16), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(KEYINPUT16), .ZN(new_n367));
  INV_X1    g181(.A(new_n358), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G146), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n255), .B1(new_n350), .B2(new_n351), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT17), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n356), .A2(new_n366), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G113), .B(G122), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(new_n208), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n364), .A2(G146), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n357), .A2(G125), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n363), .A3(new_n193), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT18), .A2(G131), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n352), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n352), .A2(new_n380), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n373), .A2(new_n375), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT90), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n350), .A2(new_n255), .A3(new_n351), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(new_n371), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n353), .A2(KEYINPUT90), .A3(new_n355), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n364), .A2(KEYINPUT19), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n377), .A2(new_n363), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n390), .B(new_n193), .C1(KEYINPUT19), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n370), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(KEYINPUT91), .B(new_n383), .C1(new_n389), .C2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n375), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n387), .A2(new_n388), .A3(new_n370), .A4(new_n392), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT91), .B1(new_n397), .B2(new_n383), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n384), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n400));
  NOR2_X1   g214(.A1(G475), .A2(G902), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT92), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n401), .ZN(new_n404));
  XOR2_X1   g218(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT92), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n399), .A2(new_n408), .A3(new_n400), .A4(new_n401), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n403), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n373), .A2(new_n383), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n395), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n384), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n322), .ZN(new_n414));
  XOR2_X1   g228(.A(KEYINPUT93), .B(G475), .Z(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n187), .A2(G952), .ZN(new_n419));
  INV_X1    g233(.A(G234), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(new_n348), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(G898), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(KEYINPUT96), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AOI211_X1 g239(.A(new_n322), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G214), .B1(G237), .B2(G902), .ZN(new_n429));
  INV_X1    g243(.A(G116), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G119), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT5), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(KEYINPUT67), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G116), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n436), .A3(G119), .ZN(new_n437));
  INV_X1    g251(.A(new_n431), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(G113), .B(new_n433), .C1(new_n439), .C2(new_n432), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT2), .B(G113), .Z(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n437), .A3(new_n438), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT68), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT68), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT67), .B(G116), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n431), .B1(new_n445), .B2(G119), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n446), .B2(new_n441), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n271), .B(new_n440), .C1(new_n443), .C2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G122), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n302), .B1(new_n305), .B2(new_n293), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n441), .B1(new_n438), .B2(new_n437), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n442), .A2(KEYINPUT68), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n446), .A2(new_n444), .A3(new_n441), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n448), .B(new_n449), .C1(new_n450), .C2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G224), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(G953), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT7), .ZN(new_n459));
  AOI211_X1 g273(.A(G125), .B(new_n206), .C1(new_n233), .C2(new_n235), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n230), .A2(new_n204), .A3(new_n297), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT64), .B(G143), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n197), .B1(new_n462), .B2(new_n193), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n461), .B1(new_n463), .B2(new_n299), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G125), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n459), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n284), .A2(new_n360), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n468), .A2(KEYINPUT7), .A3(new_n458), .A4(new_n465), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n455), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n452), .A2(new_n453), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n440), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n239), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(new_n448), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(KEYINPUT88), .A3(new_n239), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n449), .B(KEYINPUT8), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(G902), .B1(new_n470), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n448), .B1(new_n450), .B2(new_n454), .ZN(new_n480));
  INV_X1    g294(.A(new_n449), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n457), .B1(new_n460), .B2(new_n466), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n468), .A2(new_n458), .A3(new_n465), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n480), .A2(new_n487), .A3(new_n481), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G210), .B1(G237), .B2(G902), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n479), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n479), .B2(new_n489), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n428), .B(new_n429), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G217), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n343), .A2(new_n494), .A3(G953), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT66), .B(G128), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G143), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n228), .A2(G128), .A3(new_n229), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n248), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n445), .A2(G122), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n430), .A2(G122), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n210), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n210), .B1(new_n501), .B2(new_n502), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT13), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n265), .A2(KEYINPUT13), .A3(G128), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n498), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G134), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT94), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n513), .A3(G134), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n506), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n498), .A2(new_n248), .A3(new_n499), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n248), .B1(new_n498), .B2(new_n499), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n503), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT14), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n445), .A2(new_n519), .A3(G122), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT95), .B1(new_n501), .B2(KEYINPUT14), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n522));
  AOI211_X1 g336(.A(new_n522), .B(new_n519), .C1(new_n445), .C2(G122), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n502), .B(new_n520), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n518), .B1(G107), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n496), .B1(new_n515), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n505), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n516), .B1(new_n527), .B2(new_n503), .ZN(new_n528));
  INV_X1    g342(.A(new_n514), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n513), .B1(new_n510), .B2(G134), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n517), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n504), .B1(new_n532), .B2(new_n500), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n520), .A2(new_n502), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n501), .A2(KEYINPUT14), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n522), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n501), .A2(KEYINPUT95), .A3(KEYINPUT14), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n533), .B1(new_n538), .B2(new_n210), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n539), .A3(new_n495), .ZN(new_n540));
  AOI21_X1  g354(.A(G902), .B1(new_n526), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G478), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  AOI211_X1 g359(.A(G902), .B(new_n543), .C1(new_n526), .C2(new_n540), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n418), .A2(new_n493), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n341), .A2(new_n347), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT25), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT22), .B(G137), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n342), .A2(new_n420), .A3(G953), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n553), .B(new_n554), .Z(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT23), .B1(new_n199), .B2(G119), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n199), .A2(G119), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n200), .A2(new_n202), .A3(G119), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT23), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n558), .B1(new_n497), .B2(G119), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT24), .B(G110), .Z(new_n564));
  OAI22_X1  g378(.A1(new_n562), .A2(G110), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n370), .A2(new_n565), .A3(new_n378), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n562), .A2(G110), .B1(new_n563), .B2(new_n564), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n358), .B1(new_n364), .B2(KEYINPUT16), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(new_n193), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n567), .B1(new_n569), .B2(new_n365), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n556), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n570), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT76), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT76), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n566), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n571), .B1(new_n576), .B2(new_n556), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n552), .B1(new_n577), .B2(G902), .ZN(new_n578));
  INV_X1    g392(.A(new_n575), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n574), .B1(new_n566), .B2(new_n570), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n556), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n571), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(KEYINPUT25), .A3(new_n322), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n494), .B1(G234), .B2(new_n322), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(G902), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n585), .A2(new_n586), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT69), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n309), .B2(new_n464), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n301), .A2(KEYINPUT69), .A3(new_n257), .ZN(new_n592));
  INV_X1    g406(.A(new_n252), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n248), .A2(G137), .ZN(new_n594));
  OAI21_X1  g408(.A(G131), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n256), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n591), .B(new_n592), .C1(new_n284), .C2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT30), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT70), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n309), .A2(new_n464), .A3(new_n590), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT69), .B1(new_n301), .B2(new_n257), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT70), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n279), .A2(new_n256), .A3(new_n595), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT30), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  OAI22_X1  g420(.A1(new_n284), .A2(new_n596), .B1(new_n309), .B2(new_n464), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n598), .ZN(new_n608));
  OAI22_X1  g422(.A1(new_n443), .A2(new_n447), .B1(new_n446), .B2(new_n441), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT73), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT71), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n454), .B(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n597), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT26), .B(G101), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n348), .A2(new_n187), .A3(G210), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n612), .A2(new_n613), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n610), .B1(new_n599), .B2(new_n605), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n454), .B(KEYINPUT71), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n604), .A3(new_n602), .ZN(new_n626));
  INV_X1    g440(.A(new_n621), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT73), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n623), .A2(KEYINPUT31), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n624), .A2(new_n628), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT31), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT28), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n615), .B2(new_n607), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n625), .A2(KEYINPUT28), .A3(new_n604), .A4(new_n602), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n607), .A2(new_n609), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n631), .A2(new_n632), .B1(new_n621), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(G472), .A2(G902), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n640), .B(KEYINPUT74), .Z(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT32), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n615), .A2(new_n597), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT28), .B1(new_n647), .B2(new_n616), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n648), .A2(KEYINPUT29), .A3(new_n627), .A4(new_n634), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n627), .B1(new_n612), .B2(new_n626), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT29), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n637), .B2(new_n621), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n649), .B(new_n322), .C1(new_n650), .C2(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n639), .A2(new_n646), .B1(new_n653), .B2(G472), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n589), .B1(new_n645), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n551), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT97), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n213), .ZN(G3));
  AOI21_X1  g472(.A(new_n641), .B1(new_n630), .B2(new_n638), .ZN(new_n659));
  INV_X1    g473(.A(G472), .ZN(new_n660));
  AOI21_X1  g474(.A(G902), .B1(new_n630), .B2(new_n638), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n639), .A2(new_n322), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT98), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n659), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AOI211_X1 g480(.A(G469), .B(G902), .C1(new_n337), .C2(new_n338), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n331), .A2(new_n333), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n668), .B2(KEYINPUT87), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n346), .B1(new_n669), .B2(new_n334), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n666), .A2(new_n670), .A3(new_n588), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n515), .A2(new_n525), .A3(new_n496), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n495), .B1(new_n531), .B2(new_n539), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT99), .B1(new_n531), .B2(new_n539), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT33), .ZN(new_n675));
  OAI22_X1  g489(.A1(new_n672), .A2(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n515), .B2(new_n525), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n526), .A2(new_n678), .A3(KEYINPUT33), .A4(new_n540), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(G478), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n542), .A2(new_n322), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n541), .B2(new_n542), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n410), .B2(new_n417), .ZN(new_n685));
  INV_X1    g499(.A(new_n493), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n671), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT34), .B(G104), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G6));
  NAND3_X1  g504(.A1(new_n399), .A2(new_n401), .A3(new_n405), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n405), .B1(new_n399), .B2(new_n401), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n414), .A2(KEYINPUT100), .A3(new_n416), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT100), .ZN(new_n696));
  AOI21_X1  g510(.A(G902), .B1(new_n412), .B2(new_n384), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n696), .B1(new_n697), .B2(new_n415), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n695), .B(new_n698), .C1(new_n545), .C2(new_n546), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n493), .A2(new_n694), .A3(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n666), .A2(new_n670), .A3(new_n588), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT101), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT35), .B(G107), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G9));
  AOI21_X1  g518(.A(KEYINPUT25), .B1(new_n583), .B2(new_n322), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n552), .B(G902), .C1(new_n581), .C2(new_n582), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n586), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n556), .A2(KEYINPUT36), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n576), .B(new_n708), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n587), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n639), .A2(new_n662), .A3(new_n322), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G472), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n661), .A2(new_n662), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n643), .B(new_n711), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n666), .A2(KEYINPUT102), .A3(new_n711), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n718), .A3(new_n551), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT37), .B(G110), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G12));
  NAND2_X1  g535(.A1(new_n639), .A2(new_n646), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n653), .A2(G472), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n722), .B(new_n723), .C1(KEYINPUT32), .C2(new_n659), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n695), .A2(new_n698), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n407), .A2(new_n691), .ZN(new_n726));
  INV_X1    g540(.A(G900), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n422), .B1(new_n426), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n548), .A2(new_n725), .A3(new_n726), .A4(new_n729), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n585), .A2(new_n586), .B1(new_n587), .B2(new_n709), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n429), .B1(new_n491), .B2(new_n492), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n724), .A2(new_n341), .A3(new_n347), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G128), .ZN(G30));
  XOR2_X1   g549(.A(new_n728), .B(KEYINPUT39), .Z(new_n736));
  NAND2_X1  g550(.A1(new_n670), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT103), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT40), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(KEYINPUT40), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n621), .B1(new_n647), .B2(new_n616), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n623), .A2(new_n629), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(G472), .B1(new_n742), .B2(G902), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n743), .B(new_n722), .C1(KEYINPUT32), .C2(new_n659), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n731), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n491), .A2(new_n492), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT38), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n410), .A2(new_n417), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n547), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n429), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n745), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n739), .A2(new_n740), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n462), .ZN(G45));
  INV_X1    g567(.A(new_n684), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n418), .A2(new_n754), .A3(new_n729), .ZN(new_n755));
  INV_X1    g569(.A(new_n429), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n479), .A2(new_n489), .ZN(new_n757));
  INV_X1    g571(.A(new_n490), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n479), .A2(new_n489), .A3(new_n490), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n756), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n711), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n755), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(new_n724), .A3(new_n347), .A4(new_n341), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G146), .ZN(G48));
  NAND2_X1  g579(.A1(new_n337), .A2(new_n338), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n322), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(G469), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n340), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n345), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n655), .A2(new_n686), .A3(new_n685), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(KEYINPUT41), .B(G113), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G15));
  NAND3_X1  g587(.A1(new_n655), .A2(new_n700), .A3(new_n770), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G116), .ZN(G18));
  INV_X1    g589(.A(new_n345), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n768), .A2(new_n776), .A3(new_n761), .A4(new_n340), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n427), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n418), .A2(new_n731), .A3(new_n548), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n724), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G119), .ZN(G21));
  NAND2_X1  g595(.A1(new_n648), .A2(new_n634), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n782), .A2(new_n621), .B1(new_n631), .B2(new_n632), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n641), .B1(new_n783), .B2(new_n630), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT104), .B(G472), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n784), .B1(new_n664), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n778), .A2(new_n588), .A3(new_n749), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(KEYINPUT105), .B(G122), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(G24));
  INV_X1    g603(.A(new_n777), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n418), .A2(new_n754), .A3(new_n729), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(new_n786), .A3(new_n711), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G125), .ZN(G27));
  INV_X1    g607(.A(KEYINPUT42), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n724), .A2(new_n588), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n759), .A2(new_n429), .A3(new_n760), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n345), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n323), .B1(new_n339), .B2(new_n320), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT106), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n330), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT106), .B1(new_n327), .B2(new_n328), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n800), .B1(new_n801), .B2(new_n330), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n798), .B1(new_n802), .B2(new_n320), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n791), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n794), .B1(new_n795), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n801), .A2(new_n330), .ZN(new_n806));
  INV_X1    g620(.A(new_n800), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n320), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n340), .A2(new_n333), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n797), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n755), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n655), .A3(KEYINPUT42), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n805), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G131), .ZN(G33));
  INV_X1    g628(.A(new_n810), .ZN(new_n815));
  INV_X1    g629(.A(new_n730), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n655), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G134), .ZN(G36));
  NAND2_X1  g632(.A1(new_n748), .A2(new_n754), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT43), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(new_n666), .A3(new_n731), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT44), .Z(new_n822));
  AOI22_X1  g636(.A1(new_n329), .A2(new_n330), .B1(KEYINPUT45), .B2(G469), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT107), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT45), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n824), .B1(new_n825), .B2(new_n802), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n823), .A2(KEYINPUT107), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n333), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT46), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n667), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n830), .B1(new_n829), .B2(new_n828), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n776), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n796), .B(KEYINPUT108), .Z(new_n834));
  NAND4_X1  g648(.A1(new_n822), .A2(new_n736), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G137), .ZN(G39));
  NOR4_X1   g650(.A1(new_n724), .A2(new_n588), .A3(new_n755), .A4(new_n796), .ZN(new_n837));
  XNOR2_X1  g651(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n833), .A2(new_n838), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g655(.A(KEYINPUT110), .B(G140), .Z(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(G42));
  AND3_X1   g657(.A1(new_n747), .A2(new_n347), .A3(new_n429), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n744), .A2(new_n589), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n769), .A2(KEYINPUT49), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n819), .B1(KEYINPUT49), .B2(new_n769), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n729), .A2(new_n776), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n311), .A2(new_n319), .A3(KEYINPUT106), .ZN(new_n850));
  OAI21_X1  g664(.A(G469), .B1(new_n850), .B2(new_n800), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n849), .B1(new_n851), .B2(new_n798), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n418), .A2(new_n548), .A3(new_n761), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n744), .A2(new_n852), .A3(new_n731), .A4(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n764), .A2(new_n854), .A3(new_n792), .A4(new_n734), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n694), .A2(new_n699), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n711), .A3(new_n761), .A4(new_n729), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n645), .B2(new_n654), .ZN(new_n859));
  INV_X1    g673(.A(new_n785), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n639), .B2(new_n322), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n861), .A2(new_n731), .A3(new_n784), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n777), .A2(new_n755), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n859), .A2(new_n670), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n865), .A3(new_n764), .A4(new_n854), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n856), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n687), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n418), .A2(new_n547), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n686), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT111), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n588), .A3(new_n670), .A4(new_n666), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n719), .A2(new_n656), .A3(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n805), .A2(new_n812), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n771), .A2(new_n774), .A3(new_n787), .A4(new_n780), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n725), .A2(new_n726), .A3(new_n547), .A4(new_n729), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n879), .A2(new_n731), .A3(new_n796), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n670), .A2(new_n724), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n817), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT112), .ZN(new_n883));
  INV_X1    g697(.A(new_n784), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n884), .B(new_n711), .C1(new_n661), .C2(new_n860), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n804), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n811), .A2(KEYINPUT112), .A3(new_n862), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n867), .A2(new_n875), .A3(new_n878), .A4(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT54), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n771), .A2(new_n780), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n774), .A2(new_n787), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n893), .A3(new_n813), .A4(KEYINPUT53), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n856), .A2(new_n866), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT113), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n856), .A2(new_n866), .A3(KEYINPUT113), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n719), .A2(new_n874), .A3(new_n656), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n887), .A2(new_n886), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n817), .A3(new_n881), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT114), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n874), .A2(new_n656), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT114), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n888), .A2(new_n904), .A3(new_n905), .A4(new_n719), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n899), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n891), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n889), .A2(KEYINPUT53), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n875), .A2(new_n878), .A3(new_n888), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n911), .A2(KEYINPUT53), .ZN(new_n912));
  INV_X1    g726(.A(new_n898), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT113), .B1(new_n856), .B2(new_n866), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n910), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n909), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT115), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n820), .ZN(new_n921));
  AND4_X1   g735(.A1(new_n588), .A2(new_n921), .A3(new_n422), .A4(new_n786), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(new_n756), .A3(new_n747), .A4(new_n770), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT50), .Z(new_n924));
  NOR4_X1   g738(.A1(new_n769), .A2(new_n345), .A3(new_n421), .A4(new_n796), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n845), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n926), .A2(new_n418), .A3(new_n754), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n921), .A2(new_n925), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n929), .B2(new_n862), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n769), .A2(new_n347), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n839), .A2(new_n840), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n922), .A2(new_n834), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT51), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n931), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n931), .B2(new_n935), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n928), .A2(new_n795), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT48), .Z(new_n940));
  INV_X1    g754(.A(new_n685), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n419), .B1(new_n926), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n922), .B2(new_n790), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n938), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n920), .A2(new_n937), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(G952), .A2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n848), .B1(new_n945), .B2(new_n946), .ZN(G75));
  OAI21_X1  g761(.A(new_n890), .B1(new_n911), .B2(new_n895), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n903), .A2(new_n906), .ZN(new_n949));
  INV_X1    g763(.A(new_n894), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n913), .B2(new_n914), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n948), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n952), .A2(G210), .A3(G902), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n483), .A2(new_n488), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n486), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT55), .ZN(new_n956));
  XOR2_X1   g770(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n957));
  NOR3_X1   g771(.A1(new_n953), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n187), .A2(G952), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n956), .B1(new_n953), .B2(KEYINPUT56), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT117), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n960), .A2(KEYINPUT117), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(G51));
  AOI22_X1  g780(.A1(new_n899), .A2(new_n907), .B1(new_n889), .B2(new_n890), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT119), .B1(new_n967), .B2(new_n917), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT119), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n952), .A2(new_n969), .A3(KEYINPUT54), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT118), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n891), .A2(new_n908), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n891), .B2(new_n908), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n968), .B(new_n970), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n323), .B(KEYINPUT57), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT120), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n974), .A2(KEYINPUT120), .A3(new_n975), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n766), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n967), .A2(new_n322), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n826), .A2(new_n827), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n959), .B1(new_n980), .B2(new_n983), .ZN(G54));
  NAND3_X1  g798(.A1(new_n981), .A2(KEYINPUT58), .A3(G475), .ZN(new_n985));
  INV_X1    g799(.A(new_n399), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n987), .A2(new_n988), .A3(new_n959), .ZN(G60));
  XOR2_X1   g803(.A(new_n682), .B(KEYINPUT59), .Z(new_n990));
  NAND4_X1  g804(.A1(new_n974), .A2(new_n676), .A3(new_n679), .A4(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n959), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n920), .A2(new_n990), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(new_n680), .ZN(G63));
  NOR3_X1   g809(.A1(new_n494), .A2(new_n322), .A3(KEYINPUT60), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT60), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(G217), .B2(G902), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n967), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n959), .B1(new_n999), .B2(new_n709), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n577), .B(KEYINPUT121), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g817(.A(G953), .B1(new_n425), .B2(new_n456), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n900), .A2(new_n877), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT122), .Z(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT123), .ZN(new_n1008));
  INV_X1    g822(.A(G898), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n954), .B1(new_n1009), .B2(G953), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1008), .B(new_n1010), .ZN(G69));
  NAND2_X1  g825(.A1(new_n606), .A2(new_n608), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n390), .B1(KEYINPUT19), .B2(new_n391), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1012), .B(new_n1013), .Z(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(G900), .B2(G953), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n833), .A2(new_n655), .A3(new_n736), .A4(new_n853), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT125), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n864), .A2(new_n764), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  AND3_X1   g833(.A1(new_n1019), .A2(new_n813), .A3(new_n817), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1017), .A2(new_n835), .A3(new_n841), .A4(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1015), .B1(new_n1021), .B2(G953), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(KEYINPUT126), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT126), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n1024), .B(new_n1015), .C1(new_n1021), .C2(G953), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n752), .A2(new_n1019), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT62), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n870), .A2(new_n685), .ZN(new_n1028));
  OR4_X1    g842(.A1(new_n795), .A2(new_n738), .A3(new_n796), .A4(new_n1028), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n841), .A2(new_n835), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1014), .B1(new_n1031), .B2(G953), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1023), .A2(new_n1025), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1032), .A2(KEYINPUT124), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1034), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT124), .ZN(new_n1038));
  OAI211_X1 g852(.A(new_n1038), .B(new_n1014), .C1(new_n1031), .C2(G953), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1036), .A2(new_n1037), .A3(new_n1022), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1035), .A2(new_n1040), .ZN(G72));
  NAND3_X1  g855(.A1(new_n612), .A2(new_n626), .A3(new_n621), .ZN(new_n1042));
  OR3_X1    g856(.A1(new_n1021), .A2(new_n900), .A3(new_n877), .ZN(new_n1043));
  XNOR2_X1  g857(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n660), .A2(new_n322), .ZN(new_n1045));
  XNOR2_X1  g859(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1042), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n627), .B1(new_n624), .B2(new_n616), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1031), .A2(new_n1005), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1048), .B1(new_n1049), .B2(new_n1046), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n623), .A2(new_n629), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1046), .B1(new_n1051), .B2(new_n650), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n992), .B1(new_n916), .B2(new_n1052), .ZN(new_n1053));
  NOR3_X1   g867(.A1(new_n1047), .A2(new_n1050), .A3(new_n1053), .ZN(G57));
endmodule


