//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G236), .A3(G238), .A4(G235), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(G125), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n457), .C1(new_n458), .C2(new_n459), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n462), .A2(new_n467), .ZN(G160));
  NOR2_X1   g043(.A1(new_n458), .A2(new_n459), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G136), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n469), .A2(new_n457), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n457), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n471), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G162));
  NAND2_X1  g052(.A1(KEYINPUT4), .A2(G138), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n464), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(G102), .A2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n457), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G126), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n480), .B2(new_n481), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n457), .C1(new_n458), .C2(new_n459), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n485), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G50), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n496), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT68), .A3(G50), .ZN(new_n506));
  XOR2_X1   g081(.A(KEYINPUT5), .B(G543), .Z(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(new_n499), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n503), .A2(new_n506), .B1(G88), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n511), .A2(KEYINPUT69), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n511), .A2(KEYINPUT69), .B1(G75), .B2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n509), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n500), .A2(new_n510), .ZN(new_n520));
  INV_X1    g095(.A(G89), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT70), .B(G51), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n505), .A2(new_n525), .B1(new_n510), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n527), .B1(new_n522), .B2(new_n523), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n524), .A2(new_n528), .ZN(G168));
  NAND2_X1  g104(.A1(new_n505), .A2(G52), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n531), .B2(new_n520), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  NAND2_X1  g111(.A1(new_n505), .A2(G43), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n520), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n534), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT72), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  NAND2_X1  g123(.A1(G78), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G65), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n507), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G651), .B1(new_n508), .B2(G91), .ZN(new_n552));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(KEYINPUT73), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n554), .B(G543), .C1(new_n498), .C2(new_n497), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G299));
  INV_X1    g132(.A(G171), .ZN(G301));
  INV_X1    g133(.A(G168), .ZN(G286));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n560));
  INV_X1    g135(.A(G87), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n520), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n508), .A2(KEYINPUT74), .A3(G87), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n505), .A2(G49), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  AOI22_X1  g142(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n534), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n508), .A2(G86), .B1(new_n505), .B2(G48), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT75), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(new_n505), .A2(G47), .ZN(new_n577));
  INV_X1    g152(.A(G85), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n520), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n534), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n508), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n507), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n505), .B2(G54), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n584), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n584), .B1(new_n593), .B2(G868), .ZN(G321));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(G299), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G168), .B2(new_n596), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(G168), .B2(new_n596), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n603), .A2(KEYINPUT77), .B1(G868), .B2(new_n542), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(KEYINPUT77), .B2(new_n603), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT78), .Z(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g182(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n608));
  INV_X1    g183(.A(G111), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G2105), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n472), .A2(G123), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  AOI211_X1 g188(.A(new_n610), .B(new_n613), .C1(G135), .C2(new_n470), .ZN(new_n614));
  INV_X1    g189(.A(G2096), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n480), .A2(new_n481), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n465), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT80), .B(G2100), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND4_X1  g200(.A1(new_n616), .A2(new_n617), .A3(new_n624), .A4(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(G2427), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(KEYINPUT14), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n632), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n637), .A2(KEYINPUT82), .A3(new_n638), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n637), .A2(new_n638), .ZN(new_n644));
  INV_X1    g219(.A(G14), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n643), .A2(KEYINPUT83), .A3(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(KEYINPUT83), .B1(new_n643), .B2(new_n646), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(G401));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT84), .ZN(new_n652));
  NOR2_X1   g227(.A1(G2072), .A2(G2078), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n442), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2084), .B(G2090), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n654), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n654), .B(KEYINPUT17), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n658), .B(new_n655), .C1(new_n652), .C2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n655), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n652), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n657), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n615), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT85), .B(G2100), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT86), .ZN(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n674), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  OAI221_X1 g255(.A(new_n676), .B1(new_n674), .B2(new_n672), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT88), .ZN(new_n687));
  OR3_X1    g262(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n687), .B1(new_n684), .B2(new_n685), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n689), .B1(new_n688), .B2(new_n690), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G24), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n582), .B2(new_n694), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT90), .B(G1986), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n470), .A2(G131), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n472), .A2(G119), .ZN(new_n700));
  OR2_X1    g275(.A1(G95), .A2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n701), .B(G2104), .C1(G107), .C2(new_n457), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT89), .B(G29), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G25), .B(new_n703), .S(new_n705), .Z(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n698), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n575), .A2(G16), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT91), .ZN(new_n711));
  NOR2_X1   g286(.A1(G6), .A2(G16), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n694), .B1(new_n573), .B2(new_n574), .ZN(new_n715));
  OAI21_X1  g290(.A(KEYINPUT91), .B1(new_n715), .B2(new_n712), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT32), .B(G1981), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n714), .A2(new_n718), .A3(new_n716), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n694), .A2(G23), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n566), .A2(new_n565), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n562), .B2(new_n563), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n723), .B1(new_n725), .B2(new_n694), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT92), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(new_n723), .C1(new_n725), .C2(new_n694), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT33), .B(G1976), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT93), .Z(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n727), .A2(new_n732), .A3(new_n729), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n694), .A2(G22), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G303), .B2(G16), .ZN(new_n737));
  INV_X1    g312(.A(G1971), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n734), .A2(new_n735), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n722), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT34), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n709), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI211_X1 g319(.A(KEYINPUT94), .B(KEYINPUT34), .C1(new_n722), .C2(new_n741), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  AND3_X1   g321(.A1(new_n740), .A2(new_n735), .A3(new_n739), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n747), .A2(new_n720), .A3(new_n734), .A4(new_n721), .ZN(new_n748));
  AOI21_X1  g323(.A(KEYINPUT94), .B1(new_n748), .B2(KEYINPUT34), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n744), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(KEYINPUT36), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n744), .B(new_n752), .C1(new_n746), .C2(new_n749), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT31), .B(G11), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT30), .B(G28), .Z(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT24), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(G34), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(G34), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n704), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G160), .ZN(new_n762));
  INV_X1    g337(.A(G29), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT98), .B(G2084), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n757), .B(new_n766), .C1(new_n614), .C2(new_n705), .ZN(new_n767));
  NAND2_X1  g342(.A1(G162), .A2(new_n705), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n705), .A2(G35), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT29), .B(G2090), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n771), .A2(new_n772), .B1(new_n764), .B2(new_n765), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n694), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n694), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  INV_X1    g352(.A(new_n772), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n776), .A2(new_n777), .B1(new_n770), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n470), .A2(G140), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n472), .A2(G128), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n457), .A2(G116), .ZN(new_n782));
  OAI21_X1  g357(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n780), .B(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G29), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n704), .A2(G26), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G2067), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n767), .A2(new_n773), .A3(new_n779), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G19), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n542), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT95), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1341), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G168), .A2(new_n694), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n694), .B2(G21), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT26), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G129), .B2(new_n472), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n470), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT99), .Z(new_n806));
  MUX2_X1   g381(.A(G32), .B(new_n806), .S(G29), .Z(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT27), .B(G1996), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT100), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n800), .A2(G1966), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G29), .A2(G33), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n618), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(new_n457), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT25), .ZN(new_n815));
  NAND2_X1  g390(.A1(G103), .A2(G2104), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(G2105), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n457), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n470), .A2(G139), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n812), .B1(new_n820), .B2(G29), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT97), .B(G2072), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  AOI211_X1 g399(.A(new_n823), .B(new_n824), .C1(G1961), .C2(new_n775), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n811), .B(new_n825), .C1(new_n807), .C2(new_n810), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n694), .A2(G4), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n593), .B2(new_n694), .ZN(new_n828));
  INV_X1    g403(.A(G1348), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(G1966), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n799), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n694), .A2(G20), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT101), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT23), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G299), .B2(G16), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT102), .B(G1956), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n705), .A2(G27), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G164), .B2(new_n705), .ZN(new_n840));
  INV_X1    g415(.A(G2078), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n830), .A2(new_n832), .A3(new_n838), .A4(new_n842), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n797), .A2(new_n826), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT103), .B1(new_n754), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n846));
  INV_X1    g421(.A(new_n844), .ZN(new_n847));
  AOI211_X1 g422(.A(new_n846), .B(new_n847), .C1(new_n751), .C2(new_n753), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n845), .A2(new_n848), .ZN(G311));
  NAND2_X1  g424(.A1(new_n754), .A2(new_n844), .ZN(G150));
  NAND2_X1  g425(.A1(new_n593), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n508), .A2(G93), .B1(new_n505), .B2(G55), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT104), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n855), .A2(new_n534), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n541), .B2(new_n539), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n542), .A3(new_n856), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n852), .B(new_n860), .Z(new_n861));
  AND2_X1   g436(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(KEYINPUT39), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n862), .A2(new_n863), .A3(G860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(G860), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT37), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n864), .A2(new_n866), .ZN(G145));
  XNOR2_X1  g442(.A(new_n762), .B(new_n476), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n614), .B(new_n868), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n470), .A2(G142), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n472), .A2(G130), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n457), .A2(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n870), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT107), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n703), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n784), .B(new_n494), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n620), .B(KEYINPUT106), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n876), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n820), .B1(new_n805), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT105), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n806), .A2(new_n820), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n880), .A2(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n869), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  INV_X1    g465(.A(new_n869), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n891), .A3(new_n886), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n889), .A2(new_n892), .A3(KEYINPUT108), .A4(new_n893), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n896), .A2(KEYINPUT40), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT40), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(G395));
  XNOR2_X1  g475(.A(new_n860), .B(new_n602), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n592), .A2(G299), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n592), .A2(G299), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT41), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n909));
  NAND2_X1  g484(.A1(G305), .A2(G290), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n575), .A2(new_n582), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(G303), .B(new_n725), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(G303), .B(G288), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(new_n910), .B2(new_n911), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(KEYINPUT109), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT110), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n906), .A2(new_n920), .A3(new_n907), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n909), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n909), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(G868), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n857), .A2(new_n596), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(G295));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n925), .ZN(G331));
  NAND2_X1  g502(.A1(G286), .A2(G301), .ZN(new_n928));
  NAND2_X1  g503(.A1(G168), .A2(G171), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n860), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n904), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n858), .A2(new_n928), .A3(new_n859), .A4(new_n929), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n933), .A2(KEYINPUT111), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(KEYINPUT111), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n935), .A2(new_n936), .B1(new_n860), .B2(new_n930), .ZN(new_n937));
  INV_X1    g512(.A(new_n905), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n934), .B(new_n917), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n939), .A2(new_n893), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n917), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT43), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n938), .B1(new_n931), .B2(new_n933), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n931), .A2(new_n932), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n935), .B2(new_n936), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n943), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AND4_X1   g524(.A1(KEYINPUT43), .A2(new_n949), .A3(new_n893), .A4(new_n939), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT44), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(new_n940), .B2(new_n944), .ZN(new_n954));
  AND4_X1   g529(.A1(new_n953), .A2(new_n949), .A3(new_n893), .A4(new_n939), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n956), .ZN(G397));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n494), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(G160), .A2(G40), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1996), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT46), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n965), .B(KEYINPUT126), .Z(new_n966));
  INV_X1    g541(.A(new_n963), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n784), .B(new_n790), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI211_X1 g544(.A(new_n805), .B(new_n969), .C1(KEYINPUT46), .C2(new_n964), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n966), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n963), .A2(new_n964), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(new_n806), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n974), .B(KEYINPUT113), .Z(new_n975));
  NOR2_X1   g550(.A1(new_n967), .A2(new_n968), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n963), .A2(G1996), .A3(new_n805), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n977), .B(KEYINPUT114), .Z(new_n978));
  NOR3_X1   g553(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n707), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n703), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n703), .A2(new_n980), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n963), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n967), .A2(G1986), .A3(G290), .ZN(new_n985));
  XOR2_X1   g560(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n986));
  XNOR2_X1  g561(.A(new_n985), .B(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n972), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n979), .A2(new_n982), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(G2067), .B2(new_n784), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n990), .A2(KEYINPUT125), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n967), .B1(new_n990), .B2(KEYINPUT125), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n582), .B(G1986), .Z(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n963), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n979), .A2(new_n995), .A3(new_n983), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(G288), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n998), .A2(KEYINPUT116), .ZN(new_n999));
  INV_X1    g574(.A(G40), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n462), .A2(new_n467), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(new_n494), .A3(new_n958), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1002), .A2(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n725), .A2(G1976), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n998), .A2(KEYINPUT116), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n999), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n571), .A2(G1981), .ZN(new_n1007));
  INV_X1    g582(.A(G1981), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n569), .A2(new_n570), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(KEYINPUT49), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT117), .B(KEYINPUT49), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1011), .A2(KEYINPUT118), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT118), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1003), .B(new_n1010), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT52), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1006), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n958), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n1001), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT45), .B1(new_n494), .B2(new_n958), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n738), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n959), .A2(KEYINPUT50), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n494), .A2(new_n1025), .A3(new_n958), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1001), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1023), .B1(G2090), .B2(new_n1027), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1028), .A2(G8), .ZN(new_n1029));
  NOR2_X1   g604(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1030));
  AND2_X1   g605(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1031));
  OAI211_X1 g606(.A(G303), .B(G8), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G166), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1032), .B1(new_n1034), .B2(new_n1031), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1029), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1019), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1029), .A2(new_n1035), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1021), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1042), .A2(KEYINPUT53), .A3(new_n841), .A4(new_n961), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n961), .A2(new_n841), .A3(new_n1001), .A4(new_n1020), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1027), .A2(new_n777), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(G171), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1045), .A2(KEYINPUT123), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1044), .A2(new_n1050), .B1(new_n1027), .B2(new_n777), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1044), .A2(new_n1050), .ZN(new_n1052));
  AOI21_X1  g627(.A(G301), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1041), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(new_n1033), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n831), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1058));
  INV_X1    g633(.A(G2084), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1024), .A2(new_n1059), .A3(new_n1001), .A4(new_n1026), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G168), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1058), .A2(G286), .A3(new_n1060), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1057), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1058), .A2(G168), .A3(new_n1060), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT51), .B1(new_n1065), .B2(G8), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1048), .A2(G171), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1051), .A2(new_n1052), .A3(G301), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(KEYINPUT54), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1054), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n962), .B1(new_n959), .B2(KEYINPUT50), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1348), .B1(new_n1072), .B2(new_n1026), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1002), .A2(KEYINPUT121), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1001), .A2(new_n494), .A3(new_n1075), .A4(new_n958), .ZN(new_n1076));
  AOI21_X1  g651(.A(G2067), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1073), .A2(new_n1077), .A3(KEYINPUT122), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n790), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1027), .A2(new_n829), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT60), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(new_n1082), .A3(new_n1079), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT122), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(new_n593), .A3(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  NAND3_X1  g665(.A1(new_n1074), .A2(new_n1076), .A3(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n961), .A2(new_n964), .A3(new_n1001), .A4(new_n1020), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n542), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT59), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1096), .A3(new_n542), .ZN(new_n1097));
  XNOR2_X1  g672(.A(G299), .B(KEYINPUT57), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1956), .B1(new_n1072), .B2(new_n1026), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1021), .A2(new_n1022), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1098), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  XNOR2_X1  g679(.A(G299), .B(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n961), .A2(new_n1001), .A3(new_n1020), .A4(new_n1100), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1024), .A2(new_n1001), .A3(new_n1026), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1105), .B(new_n1106), .C1(new_n1107), .C2(G1956), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1095), .A2(new_n1097), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT60), .B(new_n592), .C1(new_n1078), .C2(new_n1083), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1103), .A2(new_n1108), .A3(KEYINPUT61), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1089), .A2(new_n1111), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1103), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1078), .A2(new_n1083), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1108), .A2(new_n593), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1071), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1063), .ZN(new_n1122));
  AOI21_X1  g697(.A(G286), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1056), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1066), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(KEYINPUT62), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1121), .A2(new_n1126), .A3(new_n1053), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1040), .B1(new_n1119), .B2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1009), .B(KEYINPUT120), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G288), .A2(G1976), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1129), .B1(new_n1016), .B2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1003), .B(KEYINPUT119), .Z(new_n1132));
  OAI22_X1  g707(.A1(new_n1038), .A2(new_n1019), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1006), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1029), .A2(new_n1035), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1062), .A2(new_n1033), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1038), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1037), .A2(KEYINPUT63), .A3(new_n1038), .A4(new_n1136), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1133), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g716(.A(KEYINPUT124), .B(new_n996), .C1(new_n1128), .C2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1112), .A2(new_n1144), .A3(new_n1145), .A4(new_n1113), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1088), .A2(new_n593), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1087), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1118), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1071), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1127), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1141), .B1(new_n1152), .B2(new_n1039), .ZN(new_n1153));
  INV_X1    g728(.A(new_n996), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1143), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n993), .B1(new_n1142), .B2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g731(.A1(new_n666), .A2(G319), .A3(new_n667), .ZN(new_n1158));
  NOR3_X1   g732(.A1(new_n691), .A2(new_n692), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g733(.A(new_n1159), .B1(new_n648), .B2(new_n649), .ZN(new_n1160));
  AOI21_X1  g734(.A(new_n1160), .B1(new_n896), .B2(new_n897), .ZN(new_n1161));
  INV_X1    g735(.A(new_n944), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n939), .A2(new_n893), .ZN(new_n1163));
  OAI21_X1  g737(.A(KEYINPUT43), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n940), .A2(new_n953), .A3(new_n949), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AND2_X1   g740(.A1(new_n1161), .A2(new_n1166), .ZN(G308));
  NAND2_X1  g741(.A1(new_n1161), .A2(new_n1166), .ZN(G225));
endmodule


