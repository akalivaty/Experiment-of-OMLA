//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1175, new_n1176,
    new_n1177, new_n1179, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1239,
    new_n1240, new_n1241;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(G355));
  AOI22_X1  g0003(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT67), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G50), .A2(G226), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g0009(.A(new_n209), .B1(G77), .B2(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n205), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT68), .Z(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(G58), .A2(G68), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT66), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(KEYINPUT66), .A2(G20), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n224), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n218), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n221), .A2(new_n231), .A3(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n216), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  OAI21_X1  g0051(.A(G20), .B1(new_n223), .B2(G50), .ZN(new_n252));
  INV_X1    g0052(.A(G150), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n229), .A2(G33), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n252), .B1(new_n253), .B2(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n230), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  INV_X1    g0061(.A(G13), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n262), .A2(new_n226), .A3(G1), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n258), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n260), .B1(new_n265), .B2(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n264), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT69), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT9), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G222), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n272), .B(new_n274), .C1(new_n275), .C2(new_n273), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n276), .B(new_n279), .C1(G77), .C2(new_n272), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n281), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G226), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n280), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(G200), .B2(new_n288), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n271), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n288), .A2(G179), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n268), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT14), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n284), .B1(new_n285), .B2(new_n208), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT70), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G97), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n212), .A2(G1698), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(G226), .B2(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G33), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n302), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n279), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n301), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT13), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT13), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n301), .A2(new_n314), .A3(new_n311), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n299), .B1(new_n316), .B2(G169), .ZN(new_n317));
  AOI211_X1 g0117(.A(KEYINPUT14), .B(new_n295), .C1(new_n313), .C2(new_n315), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT71), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n313), .A2(new_n321), .A3(new_n315), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n301), .A2(KEYINPUT71), .A3(new_n314), .A4(new_n311), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n254), .A2(G50), .B1(G20), .B2(new_n207), .ZN(new_n327));
  INV_X1    g0127(.A(G77), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n256), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n260), .ZN(new_n330));
  XOR2_X1   g0130(.A(new_n330), .B(KEYINPUT11), .Z(new_n331));
  NOR2_X1   g0131(.A1(new_n267), .A2(new_n207), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n265), .A2(new_n207), .A3(G13), .A4(G20), .ZN(new_n333));
  XOR2_X1   g0133(.A(new_n333), .B(KEYINPUT12), .Z(new_n334));
  NOR3_X1   g0134(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n326), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n316), .A2(G200), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n335), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n289), .B1(new_n322), .B2(new_n323), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n257), .ZN(new_n343));
  AND2_X1   g0143(.A1(KEYINPUT66), .A2(G20), .ZN(new_n344));
  NOR2_X1   g0144(.A1(KEYINPUT66), .A2(G20), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n343), .A2(new_n254), .B1(new_n346), .B2(G77), .ZN(new_n347));
  XOR2_X1   g0147(.A(KEYINPUT15), .B(G87), .Z(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n347), .B1(new_n256), .B2(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n260), .B1(new_n328), .B2(new_n263), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n328), .B2(new_n267), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G238), .A2(G1698), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n272), .B(new_n353), .C1(new_n212), .C2(G1698), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n354), .B(new_n279), .C1(G107), .C2(new_n272), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n286), .A2(G244), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n284), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n352), .B1(G190), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(G200), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT73), .ZN(new_n364));
  AOI21_X1  g0164(.A(G20), .B1(new_n306), .B2(new_n308), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(KEYINPUT7), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  OAI211_X1 g0167(.A(KEYINPUT73), .B(new_n367), .C1(new_n272), .C2(G20), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g0169(.A1(KEYINPUT72), .A2(G33), .ZN(new_n370));
  NAND2_X1  g0170(.A1(KEYINPUT72), .A2(G33), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n305), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n346), .B1(new_n372), .B2(new_n308), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT7), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n207), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n211), .A2(new_n207), .ZN(new_n376));
  OAI21_X1  g0176(.A(G20), .B1(new_n376), .B2(new_n222), .ZN(new_n377));
  INV_X1    g0177(.A(G159), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(new_n255), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n363), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n260), .ZN(new_n381));
  INV_X1    g0181(.A(new_n306), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT72), .B(G33), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(KEYINPUT3), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT7), .B1(new_n384), .B2(G20), .ZN(new_n385));
  AND2_X1   g0185(.A1(KEYINPUT72), .A2(G33), .ZN(new_n386));
  NOR2_X1   g0186(.A1(KEYINPUT72), .A2(G33), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT3), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n306), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT7), .B1(new_n227), .B2(new_n228), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n207), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n379), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n381), .B1(new_n392), .B2(KEYINPUT16), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n380), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n283), .B1(new_n286), .B2(G232), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G226), .A2(G1698), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n275), .B2(G1698), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n388), .A2(new_n306), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT74), .B1(new_n400), .B2(new_n279), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT74), .ZN(new_n402));
  AOI211_X1 g0202(.A(new_n402), .B(new_n278), .C1(new_n398), .C2(new_n399), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n289), .B(new_n395), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(new_n279), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n395), .ZN(new_n406));
  INV_X1    g0206(.A(G200), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n343), .A2(new_n263), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n267), .B2(new_n343), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n394), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n413), .A2(KEYINPUT77), .A3(KEYINPUT17), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(KEYINPUT76), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n411), .B1(new_n380), .B2(new_n393), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT76), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(new_n409), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(KEYINPUT77), .A3(new_n409), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n414), .B1(new_n420), .B2(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n394), .A2(new_n412), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n320), .B(new_n395), .C1(new_n401), .C2(new_n403), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n406), .A2(new_n295), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT75), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT75), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n422), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT18), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n421), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n357), .A2(G179), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n295), .B2(new_n357), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n352), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NOR4_X1   g0235(.A1(new_n298), .A2(new_n342), .A3(new_n362), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n263), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(G116), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AOI211_X1 g0239(.A(new_n260), .B(new_n263), .C1(new_n265), .C2(G33), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G116), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT84), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n260), .B1(new_n226), .B2(G116), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n307), .A2(G97), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G283), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n447), .B(new_n448), .C1(new_n344), .C2(new_n345), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT83), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n229), .A2(KEYINPUT83), .A3(new_n448), .A4(new_n447), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n445), .B1(new_n453), .B2(KEYINPUT20), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(KEYINPUT20), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n453), .A2(new_n445), .A3(KEYINPUT20), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n439), .B(new_n444), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n384), .B1(G264), .B2(new_n273), .ZN(new_n459));
  NOR2_X1   g0259(.A1(G257), .A2(G1698), .ZN(new_n460));
  INV_X1    g0260(.A(G303), .ZN(new_n461));
  OAI22_X1  g0261(.A1(new_n459), .A2(new_n460), .B1(new_n461), .B2(new_n272), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n279), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G1), .ZN(new_n465));
  NOR2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  AND2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n465), .B(G274), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n465), .B1(new_n467), .B2(new_n466), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n469), .A2(new_n278), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G270), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n463), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n458), .A2(new_n473), .A3(G179), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n458), .A2(G169), .A3(new_n472), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT21), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT21), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n458), .A2(new_n478), .A3(G169), .A4(new_n472), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n475), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n454), .A2(new_n455), .ZN(new_n481));
  INV_X1    g0281(.A(new_n457), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n443), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n472), .A2(G200), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n462), .A2(new_n279), .B1(G270), .B2(new_n470), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G190), .A3(new_n468), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n483), .A2(new_n484), .A3(new_n439), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT85), .ZN(new_n488));
  INV_X1    g0288(.A(new_n458), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT85), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(new_n484), .A4(new_n486), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n229), .A2(G33), .A3(G97), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT19), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G87), .ZN(new_n496));
  INV_X1    g0296(.A(G97), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(new_n215), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n302), .A2(new_n494), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n346), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n388), .A2(new_n229), .A3(G68), .A4(new_n306), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n495), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(new_n260), .B1(new_n263), .B2(new_n349), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n440), .A2(new_n348), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n503), .A2(KEYINPUT81), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT81), .B1(new_n503), .B2(new_n504), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n465), .A2(new_n282), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n508), .B(new_n278), .C1(G250), .C2(new_n465), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n386), .A2(new_n387), .A3(new_n442), .ZN(new_n510));
  NOR2_X1   g0310(.A1(G238), .A2(G1698), .ZN(new_n511));
  INV_X1    g0311(.A(G244), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(G1698), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n510), .B1(new_n384), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n509), .B1(new_n514), .B2(new_n278), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G169), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n320), .B2(new_n515), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n515), .A2(new_n289), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(G200), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n440), .A2(G87), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n519), .A2(new_n503), .A3(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n507), .A2(new_n517), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n254), .A2(G77), .ZN(new_n523));
  XNOR2_X1  g0323(.A(G97), .B(G107), .ZN(new_n524));
  NOR2_X1   g0324(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(KEYINPUT6), .A2(G107), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(KEYINPUT78), .B2(KEYINPUT6), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n346), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n366), .A2(new_n368), .B1(new_n373), .B2(KEYINPUT7), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n523), .B(new_n530), .C1(new_n531), .C2(new_n215), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n260), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n437), .A2(G97), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n441), .A2(new_n497), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n533), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n469), .A2(G257), .A3(new_n278), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n468), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT79), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT79), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n542), .A3(new_n468), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n388), .A2(G244), .A3(new_n306), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n309), .A2(new_n512), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(G1698), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G250), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT4), .B1(new_n309), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n279), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n544), .A2(new_n554), .A3(new_n320), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT80), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n278), .B1(new_n549), .B2(new_n552), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n541), .A2(new_n543), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(KEYINPUT80), .A3(new_n320), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n544), .A2(new_n554), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n295), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n538), .A2(new_n557), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n544), .A2(new_n554), .A3(G190), .ZN(new_n565));
  OAI21_X1  g0365(.A(G200), .B1(new_n558), .B2(new_n559), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI211_X1 g0367(.A(new_n534), .B(new_n536), .C1(new_n532), .C2(new_n260), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT82), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n522), .A2(new_n564), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n480), .A2(new_n492), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n550), .A2(new_n273), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n384), .B(new_n573), .C1(G257), .C2(new_n273), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n370), .A2(G294), .A3(new_n371), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n278), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n468), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n469), .A2(G264), .A3(new_n278), .ZN(new_n579));
  XNOR2_X1  g0379(.A(new_n579), .B(KEYINPUT88), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n576), .A2(new_n579), .A3(new_n577), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n581), .A2(new_n320), .B1(new_n582), .B2(new_n295), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT87), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n584), .A2(KEYINPUT25), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n437), .B2(G107), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n440), .A2(G107), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT22), .ZN(new_n588));
  OAI21_X1  g0388(.A(G87), .B1(new_n344), .B2(new_n345), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(new_n309), .ZN(new_n590));
  NAND2_X1  g0390(.A1(KEYINPUT23), .A2(G107), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT23), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n346), .A2(new_n592), .A3(new_n215), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(KEYINPUT86), .A2(KEYINPUT24), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n226), .B1(new_n510), .B2(KEYINPUT23), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n384), .A2(KEYINPUT22), .A3(G87), .A4(new_n229), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n594), .A2(new_n596), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n597), .A2(new_n590), .A3(new_n591), .A4(new_n593), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n389), .A2(new_n588), .A3(new_n589), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n599), .A2(new_n602), .B1(KEYINPUT86), .B2(KEYINPUT24), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n586), .B(new_n587), .C1(new_n603), .C2(new_n381), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n584), .A2(KEYINPUT25), .ZN(new_n605));
  NOR4_X1   g0405(.A1(new_n437), .A2(G107), .A3(new_n605), .A4(new_n585), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n583), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n604), .A2(new_n606), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n581), .A2(new_n407), .B1(new_n582), .B2(new_n289), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT80), .B1(new_n560), .B2(new_n320), .ZN(new_n611));
  NOR4_X1   g0411(.A1(new_n558), .A2(new_n559), .A3(new_n556), .A4(G179), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n536), .B1(new_n532), .B2(new_n260), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n614), .A2(new_n535), .B1(new_n295), .B2(new_n562), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n613), .A2(new_n615), .B1(new_n568), .B2(new_n567), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n570), .B1(new_n616), .B2(new_n522), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n572), .A2(new_n610), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n436), .A2(new_n618), .ZN(G372));
  NAND2_X1  g0419(.A1(new_n503), .A2(new_n504), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n521), .A2(new_n518), .B1(new_n517), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n564), .A2(new_n569), .A3(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n604), .A2(new_n609), .A3(new_n606), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n480), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n607), .A2(KEYINPUT89), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT89), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n627), .B(new_n583), .C1(new_n604), .C2(new_n606), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n624), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n517), .A2(new_n620), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n503), .A2(new_n520), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n518), .A3(new_n519), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n631), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n564), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT90), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n564), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .A3(new_n522), .ZN(new_n640));
  OAI211_X1 g0440(.A(KEYINPUT90), .B(new_n632), .C1(new_n564), .C2(new_n635), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n630), .A2(new_n631), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n436), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n297), .ZN(new_n645));
  INV_X1    g0445(.A(new_n430), .ZN(new_n646));
  INV_X1    g0446(.A(new_n434), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n336), .A2(new_n326), .B1(new_n341), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n646), .B1(new_n648), .B2(new_n421), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n645), .B1(new_n649), .B2(new_n293), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n644), .A2(new_n650), .ZN(G369));
  NAND2_X1  g0451(.A1(new_n229), .A2(G13), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT27), .B1(new_n652), .B2(G1), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n346), .A2(new_n262), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(new_n265), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n653), .A2(new_n656), .A3(G213), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G343), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT91), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n489), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n625), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n480), .A2(new_n492), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n661), .ZN(new_n664));
  XOR2_X1   g0464(.A(KEYINPUT92), .B(G330), .Z(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n608), .A2(new_n659), .ZN(new_n668));
  OAI22_X1  g0468(.A1(new_n668), .A2(new_n610), .B1(new_n607), .B2(new_n660), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n480), .A2(new_n659), .ZN(new_n671));
  INV_X1    g0471(.A(new_n610), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n629), .B2(new_n660), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n670), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n232), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n498), .A2(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n224), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT29), .B1(new_n643), .B2(new_n660), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT93), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT26), .B1(new_n564), .B2(new_n635), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n631), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n477), .A2(new_n479), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(new_n607), .A3(new_n474), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n687), .B1(new_n689), .B2(new_n624), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n639), .A2(new_n632), .A3(new_n522), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(KEYINPUT29), .A3(new_n660), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n643), .A2(new_n660), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(KEYINPUT93), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n685), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n618), .A2(new_n660), .ZN(new_n698));
  INV_X1    g0498(.A(new_n581), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n515), .A2(new_n320), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n699), .A2(new_n560), .A3(new_n700), .A4(new_n485), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n699), .A2(G179), .A3(new_n560), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n515), .A3(new_n472), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n659), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n698), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n665), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n697), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n683), .B1(new_n715), .B2(G1), .ZN(G364));
  NAND2_X1  g0516(.A1(new_n654), .A2(G45), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n718), .A2(new_n265), .A3(new_n678), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n667), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n665), .B2(new_n664), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n230), .B1(G20), .B2(new_n295), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n229), .A2(G190), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n407), .A2(G179), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G179), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(G283), .A2(new_n728), .B1(new_n731), .B2(G329), .ZN(new_n732));
  INV_X1    g0532(.A(G311), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n725), .A2(new_n320), .A3(G200), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n732), .B(new_n309), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n727), .A2(new_n226), .A3(new_n289), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n461), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n725), .A2(new_n320), .A3(new_n407), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(KEYINPUT33), .B(G317), .Z(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n729), .A2(G190), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n346), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G294), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR4_X1   g0547(.A1(new_n736), .A2(new_n739), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n346), .A2(G179), .A3(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n407), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G326), .ZN(new_n751));
  INV_X1    g0551(.A(G322), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n749), .A2(G200), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n748), .B(new_n751), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT95), .ZN(new_n756));
  INV_X1    g0556(.A(new_n750), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n735), .A2(new_n328), .B1(new_n261), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n730), .A2(new_n378), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT32), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n745), .B(KEYINPUT94), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G97), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n309), .B1(new_n737), .B2(G87), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n760), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n758), .B(new_n765), .C1(G68), .C2(new_n740), .ZN(new_n766));
  INV_X1    g0566(.A(new_n728), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n766), .B1(new_n211), .B2(new_n754), .C1(new_n215), .C2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n723), .B1(new_n756), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n722), .ZN(new_n773));
  NAND3_X1  g0573(.A1(G355), .A2(new_n232), .A3(new_n272), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n247), .A2(new_n464), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n384), .A2(new_n677), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G45), .B2(new_n224), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n774), .B1(G116), .B2(new_n232), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n769), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n772), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n779), .B(new_n719), .C1(new_n664), .C2(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n721), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  NAND2_X1  g0583(.A1(new_n659), .A2(new_n352), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(KEYINPUT96), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT96), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n659), .A2(new_n786), .A3(new_n352), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n785), .A2(new_n361), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n434), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n434), .A2(new_n659), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n694), .B(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(new_n714), .ZN(new_n794));
  INV_X1    g0594(.A(new_n719), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n792), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n770), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n722), .A2(new_n770), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n328), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n767), .A2(new_n496), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n763), .B1(new_n461), .B2(new_n757), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n801), .B(new_n802), .C1(G294), .C2(new_n753), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n309), .B1(new_n741), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G311), .B2(new_n731), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n803), .B(new_n806), .C1(new_n215), .C2(new_n738), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(G116), .B2(new_n734), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n740), .A2(G150), .B1(G143), .B2(new_n753), .ZN(new_n809));
  INV_X1    g0609(.A(G137), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n810), .B2(new_n757), .C1(new_n378), .C2(new_n735), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT34), .Z(new_n812));
  OAI221_X1 g0612(.A(new_n384), .B1(new_n745), .B2(new_n211), .C1(new_n738), .C2(new_n261), .ZN(new_n813));
  INV_X1    g0613(.A(G132), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n730), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n767), .A2(new_n207), .ZN(new_n816));
  NOR4_X1   g0616(.A1(new_n812), .A2(new_n813), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n722), .B1(new_n808), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n798), .A2(new_n719), .A3(new_n800), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n796), .A2(new_n819), .ZN(G384));
  NAND2_X1  g0620(.A1(new_n422), .A2(new_n657), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n429), .A2(new_n413), .A3(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(KEYINPUT37), .B(new_n822), .C1(new_n431), .C2(new_n821), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT38), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n429), .A2(new_n821), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n415), .A2(new_n418), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n393), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n392), .A2(KEYINPUT16), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n412), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n657), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n421), .B2(new_n430), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n832), .A2(new_n427), .A3(new_n428), .ZN(new_n836));
  AND4_X1   g0636(.A1(new_n417), .A2(new_n394), .A3(new_n409), .A4(new_n412), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n417), .B1(new_n416), .B2(new_n409), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n834), .B1(new_n839), .B2(KEYINPUT100), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT100), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n826), .A2(new_n841), .A3(new_n836), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n827), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n828), .A2(new_n825), .ZN(new_n844));
  OAI211_X1 g0644(.A(KEYINPUT38), .B(new_n835), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n829), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n339), .A2(new_n340), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n336), .B(new_n659), .C1(new_n326), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n336), .A2(new_n659), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n324), .A2(new_n317), .A3(new_n318), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n341), .B(new_n849), .C1(new_n850), .C2(new_n335), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n792), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n713), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT40), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n846), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n711), .B1(new_n618), .B2(new_n660), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n853), .B1(new_n858), .B2(new_n710), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n839), .A2(KEYINPUT100), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(new_n842), .A3(new_n833), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n844), .B1(new_n861), .B2(KEYINPUT37), .ZN(new_n862));
  INV_X1    g0662(.A(new_n421), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n833), .B1(new_n863), .B2(new_n646), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n824), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT101), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(new_n866), .A3(new_n845), .ZN(new_n867));
  OAI211_X1 g0667(.A(KEYINPUT101), .B(new_n824), .C1(new_n862), .C2(new_n864), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n859), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n856), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT103), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n869), .A2(KEYINPUT103), .A3(new_n856), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n857), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n436), .A2(new_n713), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n665), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT104), .ZN(new_n878));
  INV_X1    g0678(.A(new_n874), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n868), .ZN(new_n881));
  XNOR2_X1  g0681(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n829), .A2(new_n845), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n337), .A2(new_n659), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n791), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n694), .B2(new_n790), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n888), .A2(new_n867), .A3(new_n868), .A4(new_n852), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n646), .B2(new_n657), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n685), .A2(new_n436), .A3(new_n693), .A4(new_n696), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n892), .A2(new_n650), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n891), .B(new_n893), .Z(new_n894));
  XNOR2_X1  g0694(.A(new_n880), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n265), .B2(new_n654), .ZN(new_n896));
  OAI21_X1  g0696(.A(G77), .B1(new_n211), .B2(new_n207), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n224), .A2(new_n897), .B1(G50), .B2(new_n207), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(G1), .A3(new_n262), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT99), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n529), .B(KEYINPUT97), .Z(new_n901));
  INV_X1    g0701(.A(KEYINPUT35), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n230), .B(new_n229), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(G116), .C1(new_n902), .C2(new_n901), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT98), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT36), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n896), .A2(new_n900), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT105), .ZN(G367));
  INV_X1    g0708(.A(new_n776), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n243), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n773), .B1(new_n232), .B2(new_n349), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n767), .A2(new_n497), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n735), .A2(new_n804), .B1(new_n745), .B2(new_n215), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT110), .Z(new_n914));
  OR3_X1    g0714(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n442), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT46), .B1(new_n738), .B2(new_n442), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n915), .A2(new_n916), .B1(G317), .B2(new_n731), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n914), .B(new_n917), .C1(new_n733), .C2(new_n757), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n912), .B(new_n918), .C1(G303), .C2(new_n753), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(new_n389), .C1(new_n746), .C2(new_n741), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT111), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n767), .A2(new_n328), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(G68), .B2(new_n762), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n923), .B1(new_n211), .B2(new_n738), .C1(new_n253), .C2(new_n754), .ZN(new_n924));
  AOI22_X1  g0724(.A1(G50), .A2(new_n734), .B1(new_n740), .B2(G159), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT112), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n309), .B1(new_n750), .B2(G143), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n810), .B2(new_n730), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n924), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n921), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT47), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n719), .B1(new_n910), .B2(new_n911), .C1(new_n931), .C2(new_n723), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT113), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n660), .A2(new_n633), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n517), .A3(new_n620), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n635), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n933), .B1(new_n780), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n718), .A2(new_n265), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n616), .B1(new_n568), .B2(new_n660), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n564), .B2(new_n660), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n675), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT45), .Z(new_n943));
  NOR2_X1   g0743(.A1(new_n675), .A2(new_n941), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT44), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n670), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT109), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n674), .A2(new_n949), .B1(new_n669), .B2(new_n671), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n674), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(new_n666), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n715), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n715), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n678), .B(KEYINPUT41), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n939), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n947), .A2(new_n941), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT108), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n674), .A2(new_n616), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT106), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n564), .B1(new_n940), .B2(new_n607), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n963), .A2(KEYINPUT42), .B1(new_n660), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT107), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n966), .A2(new_n967), .B1(KEYINPUT43), .B2(new_n936), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n961), .B(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n937), .B1(new_n957), .B2(new_n969), .ZN(G387));
  OR2_X1    g0770(.A1(new_n715), .A2(new_n952), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(new_n678), .A3(new_n953), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n952), .A2(new_n939), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n669), .A2(new_n780), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n384), .B1(new_n730), .B2(new_n253), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n975), .B(new_n912), .C1(G77), .C2(new_n737), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT115), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n761), .A2(new_n349), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G50), .B2(new_n753), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n977), .B(new_n979), .C1(new_n257), .C2(new_n741), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(G159), .B2(new_n750), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n207), .B2(new_n735), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT116), .Z(new_n983));
  AOI22_X1  g0783(.A1(new_n740), .A2(G311), .B1(G317), .B2(new_n753), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n461), .B2(new_n735), .C1(new_n752), .C2(new_n757), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT48), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n804), .B2(new_n745), .C1(new_n746), .C2(new_n738), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT49), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n728), .A2(G116), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n731), .A2(G326), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n989), .A2(new_n389), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n988), .B2(new_n987), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n722), .B1(new_n983), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n680), .B(KEYINPUT114), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n343), .A2(new_n261), .ZN(new_n996));
  AOI21_X1  g0796(.A(G45), .B1(new_n996), .B2(KEYINPUT50), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n995), .B(new_n997), .C1(new_n207), .C2(new_n328), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n776), .B1(new_n240), .B2(new_n464), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n272), .A2(new_n232), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(G107), .B2(new_n232), .C1(new_n680), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n773), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n994), .A2(new_n719), .A3(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n972), .B(new_n973), .C1(new_n974), .C2(new_n1004), .ZN(G393));
  AOI21_X1  g0805(.A(new_n679), .B1(new_n948), .B2(new_n953), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n954), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n941), .A2(new_n780), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G150), .A2(new_n750), .B1(new_n753), .B2(G159), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT117), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT51), .Z(new_n1011));
  NOR2_X1   g0811(.A1(new_n761), .A2(new_n328), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n389), .B1(new_n731), .B2(G143), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n767), .B2(new_n496), .C1(new_n735), .C2(new_n257), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1012), .B(new_n1014), .C1(G50), .C2(new_n740), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1011), .B(new_n1015), .C1(new_n207), .C2(new_n738), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G311), .A2(new_n753), .B1(new_n750), .B2(G317), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT52), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n309), .B1(new_n804), .B2(new_n738), .C1(new_n767), .C2(new_n215), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n746), .A2(new_n735), .B1(new_n741), .B2(new_n461), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n442), .B2(new_n745), .C1(new_n752), .C2(new_n730), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n723), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n773), .B1(new_n909), .B2(new_n250), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G97), .B2(new_n677), .ZN(new_n1025));
  OR4_X1    g0825(.A1(new_n795), .A2(new_n1008), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n948), .B2(new_n938), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1007), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(G390));
  NAND3_X1  g0829(.A1(new_n881), .A2(new_n770), .A3(new_n883), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n799), .A2(new_n257), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n754), .A2(new_n442), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1032), .B(new_n1012), .C1(G283), .C2(new_n750), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n731), .A2(G294), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n816), .B1(G87), .B2(new_n737), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n497), .A2(new_n735), .B1(new_n741), .B2(new_n215), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1036), .A2(new_n272), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n731), .A2(G125), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n814), .B2(new_n754), .C1(new_n741), .C2(new_n810), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G159), .B2(new_n762), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n750), .A2(G128), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n272), .B1(new_n767), .B2(new_n261), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT54), .B(G143), .Z(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(new_n734), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n737), .A2(G150), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT53), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1038), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n722), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1030), .A2(new_n719), .A3(new_n1031), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT118), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n659), .B(new_n790), .C1(new_n690), .C2(new_n691), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n791), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n692), .A2(new_n660), .A3(new_n789), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(KEYINPUT118), .A3(new_n887), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n852), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n885), .B1(new_n829), .B2(new_n845), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n885), .B1(new_n888), .B2(new_n852), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n884), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(G330), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n858), .B2(new_n710), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n854), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT119), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n713), .A2(new_n665), .A3(new_n792), .A4(new_n852), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT119), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1061), .A2(new_n1071), .A3(new_n1065), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1067), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1051), .B1(new_n1073), .B2(new_n938), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n1061), .A2(new_n1071), .A3(new_n1065), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1071), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n713), .A2(G330), .A3(new_n792), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n852), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n1082), .A3(new_n1068), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT120), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1080), .B1(new_n714), .B2(new_n797), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n1064), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n888), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT120), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1081), .A2(new_n1088), .A3(new_n1082), .A4(new_n1068), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1084), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n892), .B(new_n650), .C1(new_n1062), .C2(new_n875), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n679), .B1(new_n1078), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1073), .A2(new_n1093), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1074), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(G378));
  OAI21_X1  g0898(.A(new_n1092), .B1(new_n1073), .B2(new_n1093), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1100));
  XNOR2_X1  g0900(.A(new_n298), .B(new_n1100), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n270), .A2(new_n657), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1101), .B(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n874), .A2(G330), .A3(new_n1104), .ZN(new_n1105));
  OR3_X1    g0905(.A1(new_n846), .A2(new_n856), .A3(new_n855), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n869), .A2(KEYINPUT103), .A3(new_n856), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT103), .B1(new_n869), .B2(new_n856), .ZN(new_n1108));
  OAI211_X1 g0908(.A(G330), .B(new_n1106), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1103), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1105), .A2(new_n1110), .A3(new_n891), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n891), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1104), .B1(new_n874), .B2(G330), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1109), .A2(new_n1103), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1099), .A2(KEYINPUT57), .A3(new_n1111), .A4(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1116), .A2(new_n678), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT57), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1111), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1091), .B1(new_n1078), .B2(new_n1094), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT122), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1123), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1117), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1119), .A2(new_n938), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n799), .A2(new_n261), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(G33), .A2(G41), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT121), .Z(new_n1129));
  OAI211_X1 g0929(.A(new_n1129), .B(new_n261), .C1(new_n384), .C2(G41), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n728), .A2(G58), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n804), .B2(new_n730), .C1(new_n735), .C2(new_n349), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G68), .B2(new_n762), .ZN(new_n1133));
  AOI211_X1 g0933(.A(G41), .B(new_n384), .C1(new_n740), .C2(G97), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G77), .B2(new_n737), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n215), .B2(new_n754), .C1(new_n442), .C2(new_n757), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT58), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n734), .A2(G137), .B1(G128), .B2(new_n753), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n750), .A2(G125), .B1(new_n737), .B2(new_n1044), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n814), .B2(new_n741), .C1(new_n253), .C2(new_n761), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT59), .Z(new_n1145));
  AOI21_X1  g0945(.A(new_n1129), .B1(new_n731), .B2(G124), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n378), .C2(new_n767), .ZN(new_n1147));
  AND4_X1   g0947(.A1(new_n1130), .A2(new_n1139), .A3(new_n1140), .A4(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1127), .B1(new_n1148), .B2(new_n723), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n795), .B(new_n1149), .C1(new_n1104), .C2(new_n770), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1126), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1125), .A2(new_n1151), .ZN(G375));
  AOI211_X1 g0952(.A(new_n922), .B(new_n978), .C1(G283), .C2(new_n753), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n734), .A2(G107), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n731), .A2(G303), .B1(G97), .B2(new_n737), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT123), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n309), .B1(new_n741), .B2(new_n442), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G294), .B2(new_n750), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1131), .B1(new_n378), .B2(new_n738), .C1(new_n757), .C2(new_n814), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G50), .B2(new_n762), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n740), .A2(new_n1044), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n753), .A2(G137), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n389), .B1(new_n731), .B2(G128), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n735), .A2(new_n253), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1159), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n722), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n719), .B(new_n1168), .C1(new_n852), .C2(new_n771), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n207), .B2(new_n799), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1090), .B2(new_n939), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1091), .A2(new_n1084), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n956), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1094), .B2(new_n1173), .ZN(G381));
  NOR2_X1   g0974(.A1(G375), .A2(G378), .ZN(new_n1175));
  NOR4_X1   g0975(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(G387), .A2(G390), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(G407));
  INV_X1    g0978(.A(new_n1175), .ZN(new_n1179));
  OAI211_X1 g0979(.A(G407), .B(G213), .C1(G343), .C2(new_n1179), .ZN(G409));
  INV_X1    g0980(.A(KEYINPUT62), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1097), .B1(new_n1125), .B2(new_n1151), .ZN(new_n1182));
  INV_X1    g0982(.A(G213), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1183), .A2(G343), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1099), .A2(new_n956), .A3(new_n1111), .A4(new_n1115), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1151), .A2(new_n1097), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT124), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1189), .A2(KEYINPUT60), .A3(new_n1087), .A4(new_n1091), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT60), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1172), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1190), .A2(new_n678), .A3(new_n1192), .A4(new_n1093), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1193), .A2(G384), .A3(new_n1171), .ZN(new_n1194));
  AOI21_X1  g0994(.A(G384), .B1(new_n1193), .B2(new_n1171), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1188), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1171), .ZN(new_n1197));
  INV_X1    g0997(.A(G384), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1193), .A2(G384), .A3(new_n1171), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(KEYINPUT124), .A3(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1196), .A2(new_n1201), .ZN(new_n1202));
  NOR4_X1   g1002(.A1(new_n1182), .A2(new_n1184), .A3(new_n1187), .A4(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT127), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1181), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT61), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(G375), .A2(G378), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1184), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n1208), .A3(new_n1186), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1202), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1184), .A2(G2897), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1213), .A2(new_n1211), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1209), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1207), .A2(new_n1208), .A3(new_n1186), .A4(new_n1210), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1205), .A2(new_n1206), .A3(new_n1215), .A4(new_n1217), .ZN(new_n1218));
  OR2_X1    g1018(.A1(G387), .A2(new_n1028), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G387), .A2(new_n1028), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(KEYINPUT125), .A3(new_n1220), .ZN(new_n1221));
  OR3_X1    g1021(.A1(G387), .A2(KEYINPUT125), .A3(new_n1028), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(G393), .B(new_n782), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT126), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1220), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(G387), .A2(KEYINPUT126), .A3(new_n1028), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1223), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1226), .A2(new_n1219), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1224), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1218), .A2(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1216), .B(KEYINPUT63), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1234), .A2(new_n1186), .B1(new_n1211), .B2(new_n1210), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT61), .B1(new_n1235), .B2(new_n1214), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1230), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1232), .A2(new_n1237), .ZN(G405));
  NOR2_X1   g1038(.A1(new_n1175), .A2(new_n1182), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1210), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1213), .B2(new_n1239), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(new_n1231), .ZN(G402));
endmodule


