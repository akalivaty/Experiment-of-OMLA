//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n454), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n455), .A2(KEYINPUT66), .A3(G567), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT67), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n472), .A2(new_n476), .A3(new_n473), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n480), .B1(new_n470), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n470), .A2(KEYINPUT68), .ZN(new_n486));
  XNOR2_X1  g061(.A(KEYINPUT3), .B(G2104), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(new_n489), .A3(new_n473), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT69), .ZN(new_n493));
  OR2_X1    g068(.A1(G100), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n486), .A2(new_n489), .A3(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G124), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  NAND4_X1  g074(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n473), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(new_n466), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n505), .B1(new_n487), .B2(G126), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n503), .B1(new_n506), .B2(new_n473), .ZN(new_n507));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n508), .B1(KEYINPUT70), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n487), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(G102), .A2(G2104), .ZN(new_n513));
  AOI21_X1  g088(.A(G2105), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n507), .A2(new_n514), .ZN(G164));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT5), .B1(new_n519), .B2(KEYINPUT71), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n518), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(G75), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G62), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n531), .A2(new_n532), .A3(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(new_n531), .B2(G651), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n521), .B(new_n528), .C1(new_n533), .C2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XOR2_X1   g112(.A(new_n537), .B(KEYINPUT7), .Z(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(G63), .A2(G651), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n518), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n522), .A2(new_n525), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n520), .A2(G51), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n539), .A2(new_n544), .A3(new_n545), .ZN(G168));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n526), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT73), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n527), .A2(G90), .ZN(new_n552));
  INV_X1    g127(.A(G52), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n516), .A2(new_n517), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G543), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n551), .B(new_n552), .C1(new_n553), .C2(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  AOI22_X1  g132(.A1(new_n527), .A2(G81), .B1(new_n520), .B2(G43), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT74), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n543), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G651), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND3_X1  g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(new_n527), .A2(G91), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n543), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  NOR3_X1   g150(.A1(new_n555), .A2(KEYINPUT9), .A3(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n520), .B2(G53), .ZN(new_n578));
  OAI221_X1 g153(.A(new_n573), .B1(new_n574), .B2(new_n561), .C1(new_n576), .C2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G168), .ZN(G286));
  INV_X1    g155(.A(G74), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n561), .B1(new_n526), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(G49), .B2(new_n520), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n527), .A2(G87), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(new_n543), .A2(new_n554), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT77), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n527), .A2(new_n589), .A3(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n520), .A2(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n526), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(KEYINPUT76), .B1(new_n595), .B2(G651), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n595), .A2(KEYINPUT76), .A3(G651), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n591), .B(new_n592), .C1(new_n596), .C2(new_n597), .ZN(G305));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n586), .A2(new_n599), .B1(new_n555), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n543), .A2(G60), .ZN(new_n602));
  NAND2_X1  g177(.A1(G72), .A2(G543), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n561), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n601), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n520), .A2(G54), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n543), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  AND3_X1   g183(.A1(new_n527), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  AOI21_X1  g184(.A(KEYINPUT10), .B1(new_n527), .B2(G92), .ZN(new_n610));
  OAI221_X1 g185(.A(new_n607), .B1(new_n561), .B2(new_n608), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT78), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n606), .B1(new_n612), .B2(G868), .ZN(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G299), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n615), .B2(G168), .ZN(G297));
  XNOR2_X1  g192(.A(G297), .B(KEYINPUT79), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  NOR2_X1   g195(.A1(new_n564), .A2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n612), .A2(new_n619), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT80), .Z(G323));
  XNOR2_X1  g199(.A(KEYINPUT81), .B(KEYINPUT11), .ZN(new_n625));
  XNOR2_X1  g200(.A(G323), .B(new_n625), .ZN(G282));
  NOR2_X1   g201(.A1(new_n466), .A2(G2105), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n487), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  NAND2_X1  g205(.A1(KEYINPUT82), .A2(G2100), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n491), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n496), .A2(G123), .ZN(new_n634));
  OR2_X1    g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n635), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  OAI211_X1 g213(.A(new_n632), .B(new_n638), .C1(KEYINPUT82), .C2(G2100), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT83), .Z(G156));
  XOR2_X1   g215(.A(KEYINPUT85), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT15), .B(G2435), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT14), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2443), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT86), .Z(new_n661));
  XOR2_X1   g236(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n661), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n664), .B1(new_n666), .B2(new_n659), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n659), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n667), .ZN(new_n669));
  INV_X1    g244(.A(new_n659), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n661), .A2(new_n670), .A3(new_n664), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT88), .ZN(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n681), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n677), .A2(KEYINPUT20), .A3(new_n678), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  OAI221_X1 g261(.A(new_n683), .B1(KEYINPUT20), .B2(new_n684), .C1(new_n686), .C2(new_n681), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1981), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT89), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n689), .B(new_n693), .ZN(G229));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT91), .B(G16), .Z(new_n696));
  NAND2_X1  g271(.A1(G290), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G24), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n695), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n695), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(G1986), .Z(new_n702));
  NOR2_X1   g277(.A1(G16), .A2(G23), .ZN(new_n703));
  NOR2_X1   g278(.A1(G288), .A2(KEYINPUT93), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT93), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n583), .B2(new_n584), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n703), .B1(new_n707), .B2(G16), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT33), .B(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n698), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n698), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT94), .B(G1971), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(G6), .B(G305), .S(G16), .Z(new_n715));
  XOR2_X1   g290(.A(KEYINPUT32), .B(G1981), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n710), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n702), .B1(new_n718), .B2(KEYINPUT34), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n491), .A2(G131), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n496), .A2(G119), .ZN(new_n721));
  OR2_X1    g296(.A1(G95), .A2(G2105), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n722), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT90), .ZN(new_n725));
  MUX2_X1   g300(.A(G25), .B(new_n725), .S(G29), .Z(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT35), .B(G1991), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n726), .B(new_n727), .Z(new_n728));
  OAI211_X1 g303(.A(new_n719), .B(new_n728), .C1(KEYINPUT34), .C2(new_n718), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT36), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n487), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(new_n473), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n627), .A2(G103), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT25), .Z(new_n734));
  INV_X1    g309(.A(G139), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n732), .B(new_n734), .C1(new_n490), .C2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT97), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G29), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G29), .B2(G33), .ZN(new_n739));
  INV_X1    g314(.A(G2072), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G35), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G162), .B2(new_n742), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT29), .ZN(new_n745));
  INV_X1    g320(.A(G2090), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n612), .A2(G16), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT95), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G4), .B2(G16), .ZN(new_n750));
  OR3_X1    g325(.A1(new_n749), .A2(G4), .A3(G16), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G29), .A2(G32), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n627), .A2(G105), .ZN(new_n756));
  INV_X1    g331(.A(G141), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n490), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n496), .A2(G129), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT98), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n496), .A2(KEYINPUT98), .A3(G129), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT26), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n755), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT27), .B(G1996), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n747), .A2(new_n754), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n564), .A2(new_n698), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G19), .B2(new_n698), .ZN(new_n773));
  INV_X1    g348(.A(G1341), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT23), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n698), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  NAND2_X1  g356(.A1(G171), .A2(G16), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G5), .B2(G16), .ZN(new_n783));
  INV_X1    g358(.A(G1961), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n739), .A2(new_n740), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n775), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT31), .B(G11), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n752), .A2(new_n753), .ZN(new_n789));
  AND2_X1   g364(.A1(KEYINPUT24), .A2(G34), .ZN(new_n790));
  NOR2_X1   g365(.A1(KEYINPUT24), .A2(G34), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n790), .A2(new_n791), .A3(G29), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n484), .B2(G29), .ZN(new_n793));
  INV_X1    g368(.A(G2084), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n637), .A2(new_n742), .ZN(new_n796));
  NAND2_X1  g371(.A1(G168), .A2(G16), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G16), .B2(G21), .ZN(new_n798));
  INV_X1    g373(.A(G1966), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT99), .ZN(new_n801));
  INV_X1    g376(.A(G28), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n801), .A2(new_n802), .A3(KEYINPUT30), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(KEYINPUT30), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n801), .B1(new_n802), .B2(KEYINPUT30), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n803), .A2(new_n742), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n800), .B(new_n806), .C1(new_n799), .C2(new_n798), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n742), .A2(G27), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G164), .B2(new_n742), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G2078), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n795), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n787), .A2(new_n788), .A3(new_n789), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n742), .A2(G26), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n491), .A2(G140), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT96), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(G104), .A2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n496), .A2(G128), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n813), .B1(new_n820), .B2(new_n742), .ZN(new_n821));
  MUX2_X1   g396(.A(new_n813), .B(new_n821), .S(KEYINPUT28), .Z(new_n822));
  INV_X1    g397(.A(G2067), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n773), .A2(new_n774), .B1(new_n783), .B2(new_n784), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n771), .A2(new_n812), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n730), .A2(new_n741), .A3(new_n827), .ZN(G150));
  INV_X1    g403(.A(G150), .ZN(G311));
  AOI22_X1  g404(.A1(new_n543), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(new_n561), .ZN(new_n831));
  INV_X1    g406(.A(G93), .ZN(new_n832));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n586), .A2(new_n832), .B1(new_n555), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(KEYINPUT102), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(KEYINPUT102), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n831), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n612), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  OR3_X1    g418(.A1(new_n563), .A2(new_n837), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n837), .A2(new_n843), .ZN(new_n845));
  OAI211_X1 g420(.A(KEYINPUT103), .B(new_n831), .C1(new_n835), .C2(new_n836), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n563), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n842), .B(new_n848), .Z(new_n849));
  OAI21_X1  g424(.A(new_n839), .B1(new_n849), .B2(G860), .ZN(G145));
  NAND2_X1  g425(.A1(new_n491), .A2(G142), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n496), .A2(G130), .ZN(new_n852));
  NOR2_X1   g427(.A1(G106), .A2(G2105), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n498), .B(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n484), .B(new_n637), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G126), .ZN(new_n860));
  OAI22_X1  g435(.A1(new_n470), .A2(new_n860), .B1(new_n504), .B2(new_n466), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n861), .A2(G2105), .B1(new_n502), .B2(new_n500), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n512), .A2(new_n513), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n473), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT104), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n507), .A2(new_n514), .A3(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n765), .A3(new_n763), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n868), .B1(new_n763), .B2(new_n765), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n820), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n865), .A2(new_n867), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n766), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n875), .A3(new_n869), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n737), .B(KEYINPUT105), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n629), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT97), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n736), .B(new_n881), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n872), .A2(KEYINPUT105), .A3(new_n882), .A4(new_n876), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n879), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n880), .B1(new_n879), .B2(new_n883), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n884), .A2(new_n885), .A3(new_n724), .ZN(new_n886));
  INV_X1    g461(.A(new_n724), .ZN(new_n887));
  INV_X1    g462(.A(new_n883), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n882), .B(KEYINPUT105), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n876), .B2(new_n872), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n629), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n879), .A2(new_n880), .A3(new_n883), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n859), .B1(new_n886), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n724), .B1(new_n884), .B2(new_n885), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n887), .A3(new_n892), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n858), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g475(.A1(new_n837), .A2(new_n615), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n611), .A2(G299), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n611), .A2(G299), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n848), .B(new_n622), .ZN(new_n907));
  MUX2_X1   g482(.A(new_n906), .B(new_n904), .S(new_n907), .Z(new_n908));
  XNOR2_X1  g483(.A(G166), .B(G305), .ZN(new_n909));
  INV_X1    g484(.A(G290), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(G305), .B(G303), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(G290), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n707), .ZN(new_n915));
  INV_X1    g490(.A(new_n707), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT42), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n908), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n901), .B1(new_n920), .B2(new_n615), .ZN(G295));
  OAI21_X1  g496(.A(new_n901), .B1(new_n920), .B2(new_n615), .ZN(G331));
  INV_X1    g497(.A(new_n918), .ZN(new_n923));
  NAND2_X1  g498(.A1(G171), .A2(G286), .ZN(new_n924));
  NAND2_X1  g499(.A1(G301), .A2(G168), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n848), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n844), .A2(new_n924), .A3(new_n847), .A4(new_n925), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n906), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n927), .A2(new_n928), .B1(new_n903), .B2(new_n902), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n923), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n927), .A2(new_n928), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n904), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n935), .A2(new_n918), .A3(new_n930), .A4(new_n929), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n936), .A3(new_n895), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n933), .A2(new_n936), .A3(new_n939), .A4(new_n895), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n941), .B(KEYINPUT44), .Z(G397));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n873), .B2(G1384), .ZN(new_n944));
  INV_X1    g519(.A(G40), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n482), .B2(G2105), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n475), .A2(new_n946), .A3(new_n477), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1996), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT107), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n875), .B(new_n823), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n949), .B2(new_n767), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n952), .A2(new_n767), .B1(new_n948), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n724), .B(new_n727), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(G290), .A2(G1986), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n948), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT48), .Z(new_n962));
  INV_X1    g537(.A(new_n948), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n725), .A2(new_n727), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n955), .A2(new_n964), .B1(new_n823), .B2(new_n820), .ZN(new_n965));
  OAI22_X1  g540(.A1(new_n959), .A2(new_n962), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n953), .B2(new_n767), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n951), .A2(KEYINPUT46), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n951), .A2(KEYINPUT46), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n971));
  XNOR2_X1  g546(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n966), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n507), .B2(new_n514), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT109), .B(new_n974), .C1(new_n507), .C2(new_n514), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n943), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n862), .B2(new_n864), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n947), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n799), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n977), .A2(new_n978), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n980), .B2(new_n987), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n975), .A2(KEYINPUT110), .A3(KEYINPUT50), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n947), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n988), .A2(new_n992), .A3(new_n794), .A4(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n982), .A2(KEYINPUT115), .A3(new_n799), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n985), .A2(G168), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G8), .ZN(new_n997));
  NAND2_X1  g572(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT120), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n985), .A2(new_n994), .A3(new_n995), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1003), .A2(G8), .A3(G286), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .A4(G8), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT45), .B(new_n974), .C1(new_n865), .C2(new_n867), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n975), .A2(new_n943), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n993), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1971), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n988), .A2(new_n992), .A3(new_n993), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(G2090), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G303), .A2(G8), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n1015), .B(KEYINPUT55), .Z(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(G8), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n986), .A2(new_n993), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1018), .A2(G8), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n707), .A2(KEYINPUT111), .A3(G1976), .ZN(new_n1020));
  OAI21_X1  g595(.A(G1976), .B1(new_n704), .B2(new_n706), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1019), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT52), .ZN(new_n1025));
  OR2_X1    g600(.A1(G305), .A2(G1981), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n595), .A2(G651), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1027), .B(new_n592), .C1(new_n587), .C2(new_n586), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G1981), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(KEYINPUT49), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(G305), .B2(G1981), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1030), .B(new_n1019), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1019), .A2(new_n1020), .A3(new_n1023), .A4(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1017), .A2(new_n1025), .A3(new_n1036), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1016), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n980), .A2(new_n987), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n993), .B(new_n1042), .C1(new_n986), .C2(new_n987), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n746), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1012), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G8), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1040), .B1(new_n1041), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n1010), .B2(G2078), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1052), .B(KEYINPUT121), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1013), .A2(new_n784), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1051), .A2(G2078), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1053), .B(new_n1054), .C1(new_n1055), .C2(new_n982), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1056), .A2(G171), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT62), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1002), .A2(new_n1058), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1007), .A2(new_n1050), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT124), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1059), .A2(new_n1050), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT124), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1062), .A2(new_n1063), .A3(new_n1057), .A4(new_n1007), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(G301), .B(KEYINPUT54), .Z(new_n1066));
  NAND2_X1  g641(.A1(new_n479), .A2(KEYINPUT122), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT122), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1055), .B1(new_n478), .B2(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n944), .A2(new_n1070), .A3(new_n946), .A4(new_n1008), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1066), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1066), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1056), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1050), .A2(new_n1075), .A3(new_n1077), .A4(new_n1006), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT58), .B(G1341), .Z(new_n1079));
  NAND2_X1  g654(.A1(new_n1018), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1008), .A2(new_n949), .A3(new_n993), .A4(new_n1009), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n564), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT117), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1085), .A3(new_n564), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(KEYINPUT59), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1085), .B1(new_n1082), .B2(new_n564), .ZN(new_n1089));
  AOI211_X1 g664(.A(KEYINPUT117), .B(new_n563), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1956), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1043), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(G299), .B(KEYINPUT57), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1008), .A2(new_n993), .A3(new_n1009), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1096), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n1102));
  NOR4_X1   g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(KEYINPUT61), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1095), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1104), .A2(new_n1105), .B1(new_n1107), .B2(new_n1099), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1092), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1018), .A2(G2067), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1013), .B2(new_n753), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n612), .A2(KEYINPUT60), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1113), .B(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(KEYINPUT60), .B2(new_n612), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1092), .B(KEYINPUT119), .C1(new_n1103), .C2(new_n1108), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1111), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1100), .A2(new_n1113), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1101), .B1(new_n1119), .B2(new_n612), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1078), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  OR2_X1    g696(.A1(KEYINPUT116), .A2(KEYINPUT63), .ZN(new_n1122));
  NAND2_X1  g697(.A1(KEYINPUT116), .A2(KEYINPUT63), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1049), .A2(new_n1041), .ZN(new_n1124));
  AND4_X1   g699(.A1(new_n1017), .A2(new_n1025), .A3(new_n1036), .A4(new_n1039), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1003), .A2(G8), .A3(G168), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1122), .B(new_n1123), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1016), .B1(new_n1014), .B2(G8), .ZN(new_n1130));
  OR4_X1    g705(.A1(new_n1129), .A2(new_n1040), .A3(new_n1127), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1026), .B1(new_n1133), .B2(G288), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1019), .B(KEYINPUT113), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1025), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1017), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1134), .A2(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1132), .A2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1065), .A2(new_n1121), .A3(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(G290), .A2(G1986), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n948), .B1(new_n960), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n958), .A2(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT108), .Z(new_n1144));
  OAI21_X1  g719(.A(new_n973), .B1(new_n1140), .B2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g720(.A1(G227), .A2(new_n463), .ZN(new_n1147));
  NAND2_X1  g721(.A1(new_n657), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n1149));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g724(.A1(new_n657), .A2(KEYINPUT126), .A3(new_n1147), .ZN(new_n1151));
  AOI21_X1  g725(.A(G229), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n899), .A2(new_n941), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n1154));
  XNOR2_X1  g728(.A(new_n1153), .B(new_n1154), .ZN(G308));
  XNOR2_X1  g729(.A(new_n1153), .B(KEYINPUT127), .ZN(G225));
endmodule


