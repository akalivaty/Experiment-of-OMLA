//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1197, new_n1198, new_n1199, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1264, new_n1265, new_n1266;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n206), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n214), .A2(new_n217), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n213), .ZN(G361));
  XOR2_X1   g0026(.A(G226), .B(G232), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT67), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n230), .B(new_n231), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n220), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n221), .A2(G33), .ZN(new_n251));
  OAI22_X1  g0051(.A1(new_n251), .A2(new_n203), .B1(new_n221), .B2(G68), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n246), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT11), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT71), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT71), .A2(G1), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n257), .A2(G13), .A3(G20), .A4(new_n258), .ZN(new_n259));
  OR3_X1    g0059(.A1(new_n259), .A2(KEYINPUT12), .A3(G68), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT12), .B1(new_n259), .B2(G68), .ZN(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT71), .A2(G1), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT71), .A2(G1), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n246), .B1(new_n264), .B2(G20), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n260), .A2(new_n261), .B1(G68), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n254), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n256), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT70), .ZN(new_n275));
  AND2_X1   g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n220), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n273), .A2(new_n280), .A3(new_n256), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n275), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n277), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n272), .A2(new_n268), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT72), .B1(new_n264), .B2(new_n284), .ZN(new_n285));
  AND4_X1   g0085(.A1(KEYINPUT72), .A2(new_n257), .A3(new_n284), .A4(new_n258), .ZN(new_n286));
  OAI211_X1 g0086(.A(G238), .B(new_n283), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT13), .ZN(new_n288));
  INV_X1    g0088(.A(G232), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  AND2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n290), .B1(G226), .B2(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G97), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n277), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n282), .A2(new_n287), .A3(new_n288), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT75), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n283), .B1(new_n293), .B2(new_n294), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n257), .A2(new_n284), .A3(new_n258), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT72), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n257), .A2(new_n284), .A3(KEYINPUT72), .A4(new_n258), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n277), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n299), .B1(new_n304), .B2(G238), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT75), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n305), .A2(new_n306), .A3(new_n288), .A4(new_n282), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n282), .A2(new_n287), .A3(new_n296), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT13), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n298), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT14), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(G169), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n309), .A2(G179), .A3(new_n297), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n311), .B1(new_n310), .B2(G169), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n267), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n309), .A2(G190), .A3(new_n297), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT76), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n309), .A2(KEYINPUT76), .A3(G190), .A4(new_n297), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n267), .B1(new_n310), .B2(G200), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n321), .A2(KEYINPUT77), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT77), .B1(new_n321), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n316), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OR2_X1    g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NAND2_X1  g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(G223), .A3(G1698), .ZN(new_n329));
  INV_X1    g0129(.A(G1698), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(G222), .A3(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n329), .B(new_n331), .C1(new_n203), .C2(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n277), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n304), .A2(G226), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(new_n282), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n335), .A2(G179), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n202), .A2(new_n221), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT8), .B(G58), .ZN(new_n338));
  INV_X1    g0138(.A(G150), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n338), .A2(new_n251), .B1(new_n339), .B2(new_n248), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n246), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n259), .A2(G50), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(G50), .B2(new_n265), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n335), .A2(new_n345), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n336), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT9), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n335), .A2(G200), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n333), .A2(new_n334), .A3(G190), .A4(new_n282), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n341), .A2(KEYINPUT9), .A3(new_n343), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n349), .A2(new_n350), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT10), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(KEYINPUT10), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n347), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n328), .A2(G223), .A3(new_n330), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n328), .A2(G226), .A3(G1698), .ZN(new_n361));
  INV_X1    g0161(.A(G33), .ZN(new_n362));
  INV_X1    g0162(.A(G87), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n360), .B(new_n361), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n277), .ZN(new_n365));
  OAI211_X1 g0165(.A(G232), .B(new_n283), .C1(new_n285), .C2(new_n286), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n282), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G200), .ZN(new_n368));
  AND2_X1   g0168(.A1(G58), .A2(G68), .ZN(new_n369));
  NOR2_X1   g0169(.A1(G58), .A2(G68), .ZN(new_n370));
  OAI21_X1  g0170(.A(G20), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT79), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n247), .A2(G159), .ZN(new_n374));
  OAI211_X1 g0174(.A(KEYINPUT79), .B(G20), .C1(new_n369), .C2(new_n370), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT7), .B1(new_n328), .B2(G20), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n291), .A2(new_n292), .ZN(new_n379));
  AND2_X1   g0179(.A1(KEYINPUT78), .A2(KEYINPUT7), .ZN(new_n380));
  NOR2_X1   g0180(.A1(KEYINPUT78), .A2(KEYINPUT7), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n382), .A3(new_n221), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(new_n383), .A3(G68), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n377), .A2(KEYINPUT16), .A3(new_n384), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n386));
  INV_X1    g0186(.A(G68), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n382), .B1(new_n328), .B2(G20), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n379), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n386), .B1(new_n390), .B2(new_n376), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n385), .A2(new_n391), .A3(new_n246), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n259), .A2(new_n338), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n265), .B2(new_n338), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n365), .A2(new_n282), .A3(G190), .A4(new_n366), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n368), .A2(new_n392), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n367), .A2(G169), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n365), .A2(new_n282), .A3(G179), .A4(new_n366), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n392), .A2(new_n394), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT18), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(new_n400), .B2(new_n401), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(G244), .B(new_n283), .C1(new_n285), .C2(new_n286), .ZN(new_n406));
  OAI211_X1 g0206(.A(G238), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n326), .A2(G107), .A3(new_n327), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(G232), .B(new_n330), .C1(new_n291), .C2(new_n292), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT73), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n328), .A2(KEYINPUT73), .A3(G232), .A4(new_n330), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n282), .B(new_n406), .C1(new_n414), .C2(new_n283), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n345), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n412), .A2(new_n413), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n277), .B1(new_n417), .B2(new_n409), .ZN(new_n418));
  INV_X1    g0218(.A(G179), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(new_n419), .A3(new_n282), .A4(new_n406), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n338), .A2(new_n248), .B1(new_n221), .B2(new_n203), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT15), .B(G87), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n251), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n246), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n259), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n203), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n265), .A2(G77), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n416), .A2(new_n420), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G200), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n282), .A2(new_n406), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(new_n418), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT74), .B1(new_n432), .B2(new_n428), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n428), .B1(new_n415), .B2(G200), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT74), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n431), .A2(G190), .A3(new_n418), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n397), .A2(new_n405), .A3(new_n429), .A4(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n325), .A2(new_n359), .A3(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(G244), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n441));
  OAI211_X1 g0241(.A(G238), .B(new_n330), .C1(new_n291), .C2(new_n292), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G116), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n257), .A2(G45), .A3(new_n258), .ZN(new_n445));
  INV_X1    g0245(.A(G250), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n277), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n264), .A2(G45), .A3(new_n278), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n277), .A2(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n449), .A2(G169), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT19), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n221), .B1(new_n294), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(G97), .A2(G107), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n363), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n221), .B(G68), .C1(new_n291), .C2(new_n292), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n451), .B1(new_n251), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT84), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT84), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n455), .A2(new_n456), .A3(new_n461), .A4(new_n458), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n246), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n246), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n257), .A2(G33), .A3(new_n258), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n259), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT82), .ZN(new_n467));
  INV_X1    g0267(.A(new_n422), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT82), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n259), .A2(new_n464), .A3(new_n465), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n425), .A2(new_n422), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n463), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n449), .A2(new_n419), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n450), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G244), .B(new_n330), .C1(new_n291), .C2(new_n292), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G250), .A2(G1698), .ZN(new_n481));
  NAND2_X1  g0281(.A1(KEYINPUT4), .A2(G244), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(G1698), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n328), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n277), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT5), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G41), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n257), .A2(new_n488), .A3(G45), .A4(new_n258), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT83), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n264), .A2(new_n491), .A3(G45), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n493), .B(G274), .C1(new_n276), .C2(new_n220), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n490), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n493), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n283), .B(G257), .C1(new_n489), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n486), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n345), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n283), .B1(new_n478), .B2(new_n484), .ZN(new_n501));
  INV_X1    g0301(.A(new_n498), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n419), .A3(new_n496), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n388), .A2(new_n389), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G107), .ZN(new_n506));
  INV_X1    g0306(.A(G107), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(G97), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT81), .ZN(new_n509));
  NAND2_X1  g0309(.A1(KEYINPUT6), .A2(G97), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(G107), .ZN(new_n511));
  AND2_X1   g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(new_n453), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n508), .B(new_n511), .C1(new_n513), .C2(KEYINPUT6), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(G20), .B1(G77), .B2(new_n247), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n464), .B1(new_n506), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n467), .A2(G97), .A3(new_n470), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n425), .A2(new_n457), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n500), .B(new_n504), .C1(new_n516), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n499), .A2(G200), .ZN(new_n521));
  INV_X1    g0321(.A(new_n516), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n517), .A2(new_n518), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n486), .A2(G190), .A3(new_n496), .A4(new_n498), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n521), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n467), .A2(G87), .A3(new_n470), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT85), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n467), .A2(KEYINPUT85), .A3(G87), .A4(new_n470), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n444), .A2(new_n277), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n447), .A2(new_n448), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n531), .A2(G190), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n430), .B1(new_n531), .B2(new_n532), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n463), .A2(new_n472), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AND4_X1   g0337(.A1(new_n475), .A2(new_n520), .A3(new_n525), .A4(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT22), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n221), .A2(KEYINPUT86), .A3(G87), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n379), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n540), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n328), .A2(new_n542), .A3(KEYINPUT22), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n443), .A2(G20), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT23), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n221), .B2(G107), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n507), .A2(KEYINPUT23), .A3(G20), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n541), .A2(new_n543), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT24), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT24), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n541), .A2(new_n543), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n464), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n467), .A2(G107), .A3(new_n470), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n425), .A2(KEYINPUT25), .A3(new_n507), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT25), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n259), .B2(G107), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(G257), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n561));
  OAI211_X1 g0361(.A(G250), .B(new_n330), .C1(new_n291), .C2(new_n292), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G294), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n277), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n283), .B(G264), .C1(new_n489), .C2(new_n497), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n496), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G200), .ZN(new_n568));
  INV_X1    g0368(.A(new_n489), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n277), .B1(new_n569), .B2(new_n493), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(G264), .B1(new_n277), .B2(new_n564), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(G190), .A3(new_n496), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n560), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n419), .A3(new_n496), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n567), .A2(new_n345), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n574), .B(new_n575), .C1(new_n553), .C2(new_n559), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(G116), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n245), .A2(new_n220), .B1(G20), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n479), .B(new_n221), .C1(G33), .C2(new_n457), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT20), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(KEYINPUT20), .A3(new_n580), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n425), .A2(new_n578), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n259), .A2(new_n464), .A3(new_n465), .A4(G116), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(G264), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n589));
  OAI211_X1 g0389(.A(G257), .B(new_n330), .C1(new_n291), .C2(new_n292), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n326), .A2(G303), .A3(new_n327), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n277), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n283), .B(G270), .C1(new_n489), .C2(new_n497), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n496), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n588), .A2(new_n595), .A3(G169), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(G200), .ZN(new_n599));
  INV_X1    g0399(.A(new_n588), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n593), .A2(new_n496), .A3(G190), .A4(new_n594), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n496), .A2(new_n594), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n419), .B1(new_n592), .B2(new_n277), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n588), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n588), .A2(new_n595), .A3(KEYINPUT21), .A4(G169), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n598), .A2(new_n602), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n577), .A2(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n440), .A2(new_n538), .A3(new_n608), .ZN(G372));
  NAND2_X1  g0409(.A1(new_n356), .A2(new_n357), .ZN(new_n610));
  INV_X1    g0410(.A(new_n397), .ZN(new_n611));
  INV_X1    g0411(.A(new_n429), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n323), .B2(new_n324), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n611), .B1(new_n613), .B2(new_n316), .ZN(new_n614));
  INV_X1    g0414(.A(new_n405), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n347), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n537), .A2(new_n475), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(new_n520), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n516), .A2(new_n519), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n499), .A2(G179), .ZN(new_n622));
  AOI21_X1  g0422(.A(G169), .B1(new_n503), .B2(new_n496), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(KEYINPUT26), .A3(new_n475), .A4(new_n537), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n520), .A2(new_n525), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n537), .A2(new_n475), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n576), .A2(new_n598), .A3(new_n605), .A4(new_n606), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .A4(new_n573), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n626), .A2(new_n475), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n440), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n616), .A2(new_n617), .A3(new_n632), .ZN(G369));
  NAND3_X1  g0433(.A1(new_n598), .A2(new_n605), .A3(new_n606), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n221), .A2(G13), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n264), .A2(new_n635), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(G343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n600), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n607), .B2(new_n643), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(G330), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n560), .A2(new_n642), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n577), .A2(new_n647), .B1(new_n576), .B2(new_n642), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n634), .A2(new_n642), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n577), .ZN(new_n651));
  INV_X1    g0451(.A(new_n576), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n642), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(new_n653), .ZN(G399));
  INV_X1    g0454(.A(new_n215), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n454), .A2(G116), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G1), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n218), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT28), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT29), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n631), .A2(new_n662), .A3(new_n642), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n631), .B2(new_n642), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n608), .A2(new_n538), .A3(new_n642), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT87), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n603), .A2(new_n571), .A3(new_n449), .A4(new_n604), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n503), .A2(KEYINPUT30), .A3(new_n496), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n531), .A2(new_n565), .A3(new_n532), .A4(new_n566), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n593), .A2(new_n496), .A3(G179), .A4(new_n594), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n499), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n674), .A2(KEYINPUT87), .A3(new_n675), .A4(KEYINPUT30), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n449), .A2(G179), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(new_n499), .A3(new_n567), .A4(new_n595), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n499), .A2(new_n672), .A3(new_n673), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(KEYINPUT30), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n641), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT31), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g0484(.A(KEYINPUT31), .B(new_n641), .C1(new_n677), .C2(new_n681), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n667), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n666), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n661), .B1(new_n689), .B2(G1), .ZN(G364));
  AOI21_X1  g0490(.A(new_n256), .B1(new_n635), .B2(G45), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n656), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n646), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(G330), .B2(new_n645), .ZN(new_n695));
  INV_X1    g0495(.A(new_n693), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n220), .B1(G20), .B2(new_n345), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n221), .A2(new_n419), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(G190), .A3(new_n430), .ZN(new_n700));
  INV_X1    g0500(.A(G58), .ZN(new_n701));
  NOR2_X1   g0501(.A1(G190), .A2(G200), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  OAI22_X1  g0503(.A1(new_n700), .A2(new_n701), .B1(new_n703), .B2(new_n203), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n699), .A2(G200), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G190), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n221), .A2(G179), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n702), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G159), .ZN(new_n711));
  XOR2_X1   g0511(.A(KEYINPUT89), .B(KEYINPUT32), .Z(new_n712));
  OAI22_X1  g0512(.A1(new_n707), .A2(new_n387), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G190), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n714), .A2(G179), .A3(G200), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n221), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI211_X1 g0517(.A(new_n704), .B(new_n713), .C1(G97), .C2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n705), .A2(new_n714), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G50), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n708), .A2(new_n714), .A3(G200), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n711), .A2(new_n712), .B1(G107), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n708), .A2(G190), .A3(G200), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G87), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n328), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT90), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n718), .A2(new_n720), .A3(new_n723), .A4(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G322), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n700), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G311), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n379), .B1(new_n703), .B2(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n731), .B(new_n733), .C1(G329), .C2(new_n710), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n719), .A2(G326), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT33), .B(G317), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n706), .A2(new_n736), .B1(new_n725), .B2(G303), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n717), .A2(G294), .B1(new_n722), .B2(G283), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n734), .A2(new_n735), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n698), .B1(new_n729), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n697), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n328), .A2(G355), .A3(new_n215), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(G116), .B2(new_n215), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT88), .Z(new_n747));
  NOR2_X1   g0547(.A1(new_n655), .A2(new_n328), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n269), .A2(new_n271), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n748), .B1(new_n219), .B2(new_n749), .C1(new_n243), .C2(new_n268), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n696), .B(new_n740), .C1(new_n744), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n743), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(new_n645), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n695), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(G396));
  NAND2_X1  g0556(.A1(new_n641), .A2(new_n428), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n437), .B1(new_n434), .B2(new_n435), .ZN(new_n758));
  AOI211_X1 g0558(.A(KEYINPUT74), .B(new_n428), .C1(new_n415), .C2(G200), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT93), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n429), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n428), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n415), .B2(new_n345), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(KEYINPUT93), .A3(new_n420), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(KEYINPUT94), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  AND4_X1   g0567(.A1(KEYINPUT93), .A2(new_n416), .A3(new_n420), .A4(new_n428), .ZN(new_n768));
  AOI21_X1  g0568(.A(KEYINPUT93), .B1(new_n764), .B2(new_n420), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT94), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n770), .A2(new_n771), .A3(new_n438), .A4(new_n757), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(new_n631), .A3(new_n642), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n631), .A2(new_n642), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n767), .B(new_n772), .C1(new_n429), .C2(new_n642), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n693), .B1(new_n777), .B2(new_n688), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n688), .B2(new_n777), .ZN(new_n779));
  INV_X1    g0579(.A(new_n719), .ZN(new_n780));
  INV_X1    g0580(.A(G303), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n781), .B1(new_n721), .B2(new_n363), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(G107), .B2(new_n725), .ZN(new_n783));
  INV_X1    g0583(.A(G294), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n700), .A2(new_n784), .B1(new_n703), .B2(new_n578), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n328), .B(new_n785), .C1(G311), .C2(new_n710), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G97), .A2(new_n717), .B1(new_n706), .B2(G283), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n783), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G137), .A2(new_n719), .B1(new_n706), .B2(G150), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT91), .Z(new_n790));
  INV_X1    g0590(.A(new_n700), .ZN(new_n791));
  INV_X1    g0591(.A(new_n703), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n791), .A2(G143), .B1(new_n792), .B2(G159), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT92), .B(KEYINPUT34), .Z(new_n794));
  NAND3_X1  g0594(.A1(new_n790), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n722), .A2(G68), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n379), .B1(new_n710), .B2(G132), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n717), .A2(G58), .B1(new_n725), .B2(G50), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n795), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n794), .B1(new_n790), .B2(new_n793), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n788), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n697), .A2(new_n741), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n801), .A2(new_n697), .B1(new_n203), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n776), .B2(new_n742), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n693), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n779), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT95), .Z(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G384));
  INV_X1    g0608(.A(KEYINPUT40), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n267), .A2(new_n641), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n325), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n316), .B(new_n810), .C1(new_n323), .C2(new_n324), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT97), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n686), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n667), .A2(new_n684), .A3(KEYINPUT97), .A4(new_n685), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n814), .A2(new_n776), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT38), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT37), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n400), .A2(new_n401), .ZN(new_n821));
  INV_X1    g0621(.A(new_n639), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n401), .A2(new_n822), .ZN(new_n823));
  AND4_X1   g0623(.A1(new_n820), .A2(new_n821), .A3(new_n823), .A4(new_n396), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n385), .A2(new_n246), .ZN(new_n825));
  INV_X1    g0625(.A(new_n386), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n377), .B2(new_n384), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n394), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n822), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT96), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n828), .A2(KEYINPUT96), .A3(new_n822), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n400), .A2(new_n828), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n831), .A2(new_n396), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n824), .B1(KEYINPUT37), .B2(new_n834), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n828), .A2(KEYINPUT96), .A3(new_n822), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT96), .B1(new_n828), .B2(new_n822), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n397), .B2(new_n405), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n819), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n821), .A2(KEYINPUT18), .ZN(new_n841));
  INV_X1    g0641(.A(new_n401), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n842), .A2(KEYINPUT17), .A3(new_n395), .A4(new_n368), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT17), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n396), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n841), .A2(new_n843), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n831), .A2(new_n832), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n833), .A2(new_n396), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n820), .B1(new_n838), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n849), .B(KEYINPUT38), .C1(new_n851), .C2(new_n824), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n840), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n809), .B1(new_n818), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n812), .A2(new_n813), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n816), .A2(new_n776), .A3(new_n817), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n821), .A2(new_n823), .A3(new_n396), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(new_n820), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n823), .B1(new_n397), .B2(new_n405), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n819), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n809), .B1(new_n862), .B2(new_n852), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n855), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n816), .A2(new_n817), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n866), .A2(new_n440), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n865), .A2(new_n867), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n868), .A2(G330), .A3(new_n869), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n840), .A2(KEYINPUT39), .A3(new_n852), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT39), .B1(new_n862), .B2(new_n852), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n316), .A2(new_n641), .ZN(new_n873));
  OR3_X1    g0673(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n766), .A2(new_n642), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n774), .A2(new_n875), .B1(new_n812), .B2(new_n813), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n853), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n615), .A2(new_n639), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n874), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n440), .B1(new_n663), .B2(new_n664), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n616), .A3(new_n617), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n879), .B(new_n881), .Z(new_n882));
  OAI22_X1  g0682(.A1(new_n870), .A2(new_n882), .B1(new_n264), .B2(new_n635), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n882), .B2(new_n870), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n578), .B(new_n223), .C1(new_n514), .C2(KEYINPUT35), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(KEYINPUT35), .B2(new_n514), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n886), .B(KEYINPUT36), .Z(new_n887));
  OR3_X1    g0687(.A1(new_n218), .A2(new_n369), .A3(new_n203), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n249), .A2(G68), .ZN(new_n889));
  AOI211_X1 g0689(.A(G13), .B(new_n264), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  OR3_X1    g0690(.A1(new_n884), .A2(new_n887), .A3(new_n890), .ZN(G367));
  AOI21_X1  g0691(.A(new_n642), .B1(new_n530), .B2(new_n536), .ZN(new_n892));
  INV_X1    g0692(.A(new_n475), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n619), .B2(new_n892), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n753), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n235), .A2(new_n748), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n897), .B(new_n744), .C1(new_n215), .C2(new_n422), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT103), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n696), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n898), .ZN(new_n901));
  INV_X1    g0701(.A(G283), .ZN(new_n902));
  INV_X1    g0702(.A(G317), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n703), .A2(new_n902), .B1(new_n709), .B2(new_n903), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n328), .B(new_n904), .C1(G303), .C2(new_n791), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n725), .A2(G116), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT46), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n719), .A2(G311), .B1(new_n722), .B2(G97), .ZN(new_n908));
  AOI22_X1  g0708(.A1(G107), .A2(new_n717), .B1(new_n706), .B2(G294), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n905), .A2(new_n907), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT104), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n716), .A2(new_n387), .B1(new_n700), .B2(new_n339), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n912), .B(KEYINPUT105), .Z(new_n913));
  INV_X1    g0713(.A(G159), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n707), .A2(new_n914), .B1(new_n724), .B2(new_n701), .ZN(new_n915));
  INV_X1    g0715(.A(G143), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n780), .A2(new_n916), .B1(new_n721), .B2(new_n203), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n379), .B1(new_n710), .B2(G137), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n249), .B2(new_n703), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n915), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n911), .B1(new_n913), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT47), .Z(new_n922));
  AOI211_X1 g0722(.A(new_n896), .B(new_n901), .C1(new_n922), .C2(new_n697), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n656), .B(KEYINPUT41), .Z(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  MUX2_X1   g0725(.A(new_n577), .B(new_n648), .S(new_n650), .Z(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(new_n646), .Z(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n687), .A3(new_n665), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT102), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n689), .A2(KEYINPUT102), .A3(new_n927), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n627), .B1(new_n621), .B2(new_n642), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n624), .A2(new_n641), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(KEYINPUT100), .A2(KEYINPUT44), .ZN(new_n935));
  OR3_X1    g0735(.A1(new_n653), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n653), .B2(new_n934), .ZN(new_n937));
  NAND2_X1  g0737(.A1(KEYINPUT100), .A2(KEYINPUT44), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n653), .A2(new_n934), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT99), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT99), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n653), .A2(new_n942), .A3(new_n934), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n941), .A2(KEYINPUT45), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n649), .A2(KEYINPUT101), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT45), .B1(new_n941), .B2(new_n943), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n945), .A2(new_n948), .B1(KEYINPUT101), .B2(new_n649), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n930), .A2(new_n931), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n689), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n925), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n691), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n646), .A2(new_n648), .A3(new_n934), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT98), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n895), .A2(KEYINPUT43), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n934), .A2(new_n651), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n520), .B1(new_n932), .B2(new_n576), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n961), .A2(KEYINPUT42), .B1(new_n963), .B2(new_n642), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n962), .A2(new_n964), .B1(KEYINPUT43), .B2(new_n895), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OR3_X1    g0766(.A1(new_n959), .A2(new_n960), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n966), .B1(new_n959), .B2(new_n960), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n923), .B1(new_n955), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(G387));
  AND2_X1   g0772(.A1(new_n928), .A2(new_n656), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n689), .B2(new_n927), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n927), .A2(new_n692), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n658), .A2(new_n379), .A3(new_n655), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n507), .B2(new_n655), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT106), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n232), .B1(new_n269), .B2(new_n271), .ZN(new_n979));
  INV_X1    g0779(.A(new_n338), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n249), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT50), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n658), .B(new_n268), .C1(new_n387), .C2(new_n203), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n748), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n978), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n696), .B1(new_n985), .B2(new_n744), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n468), .A2(new_n717), .B1(new_n706), .B2(new_n980), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n203), .B2(new_n724), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n328), .B1(new_n700), .B2(new_n249), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n703), .A2(new_n387), .B1(new_n709), .B2(new_n339), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n780), .A2(new_n914), .B1(new_n721), .B2(new_n457), .ZN(new_n991));
  NOR4_X1   g0791(.A1(new_n988), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n791), .A2(G317), .B1(new_n792), .B2(G303), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n780), .B2(new_n730), .C1(new_n732), .C2(new_n707), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT48), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n717), .A2(G283), .B1(new_n725), .B2(G294), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT49), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n1000), .A2(KEYINPUT107), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n328), .B1(new_n710), .B2(G326), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n578), .B2(new_n721), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n1000), .B2(KEYINPUT107), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n992), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n986), .B1(new_n648), .B2(new_n753), .C1(new_n1005), .C2(new_n698), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n975), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n974), .A2(new_n1007), .ZN(G393));
  INV_X1    g0808(.A(KEYINPUT108), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n649), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n646), .A2(KEYINPUT108), .A3(new_n648), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n946), .A2(new_n949), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1009), .B(new_n649), .C1(new_n945), .C2(new_n948), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n691), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n932), .A2(new_n743), .A3(new_n933), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n240), .A2(new_n748), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n744), .B1(new_n457), .B2(new_n215), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n693), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n780), .A2(new_n903), .B1(new_n732), .B2(new_n700), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT52), .Z(new_n1020));
  OAI221_X1 g0820(.A(new_n379), .B1(new_n709), .B2(new_n730), .C1(new_n784), .C2(new_n703), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n707), .A2(new_n781), .B1(new_n721), .B2(new_n507), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n716), .A2(new_n578), .B1(new_n724), .B2(new_n902), .ZN(new_n1023));
  OR4_X1    g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT110), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n780), .A2(new_n339), .B1(new_n914), .B2(new_n700), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT51), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n724), .A2(new_n387), .B1(new_n709), .B2(new_n916), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(KEYINPUT109), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(KEYINPUT109), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n716), .A2(new_n203), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n328), .B1(new_n703), .B2(new_n338), .C1(new_n363), .C2(new_n721), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(G50), .C2(new_n706), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1024), .A2(KEYINPUT110), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1025), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1018), .B1(new_n1036), .B2(new_n697), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1014), .B1(new_n1015), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n931), .A2(new_n930), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n950), .A2(new_n951), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n657), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1012), .A2(new_n928), .A3(new_n1013), .ZN(new_n1042));
  AND3_X1   g0842(.A1(new_n1041), .A2(KEYINPUT111), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT111), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1038), .B1(new_n1043), .B2(new_n1044), .ZN(G390));
  AND4_X1   g0845(.A1(G330), .A2(new_n816), .A3(new_n776), .A4(new_n817), .ZN(new_n1046));
  AND4_X1   g0846(.A1(new_n774), .A2(new_n812), .A3(new_n813), .A4(new_n875), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1046), .B1(new_n1047), .B2(new_n876), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n774), .A2(new_n875), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n814), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n688), .A2(new_n776), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n774), .A2(new_n812), .A3(new_n813), .A4(new_n875), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n440), .A2(new_n816), .A3(G330), .A4(new_n817), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1055), .A2(new_n880), .A3(new_n616), .A4(new_n617), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1054), .A2(KEYINPUT113), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT113), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1046), .A2(new_n814), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n873), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n871), .A2(new_n872), .B1(new_n876), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT112), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n862), .A2(new_n852), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1050), .A2(new_n1064), .A3(new_n873), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n876), .A2(new_n1062), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1064), .B1(new_n1068), .B2(new_n1065), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1061), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1050), .A2(new_n873), .A3(new_n1065), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(KEYINPUT112), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n814), .A2(new_n688), .A3(new_n776), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1072), .A2(new_n1073), .A3(new_n1063), .A4(new_n1066), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1060), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n657), .B1(new_n1078), .B2(new_n1075), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n741), .B1(new_n871), .B2(new_n872), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n802), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n693), .B1(new_n1082), .B2(new_n980), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n703), .A2(new_n457), .B1(new_n709), .B2(new_n784), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n328), .B(new_n1084), .C1(G116), .C2(new_n791), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n726), .A3(new_n796), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1031), .B1(G283), .B2(new_n719), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n507), .B2(new_n707), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n724), .A2(new_n339), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G159), .A2(new_n717), .B1(new_n719), .B2(G128), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n379), .B1(new_n791), .B2(G132), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n792), .A2(new_n1095), .B1(new_n710), .B2(G125), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n706), .A2(G137), .B1(new_n722), .B2(G50), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1092), .A2(new_n1093), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1086), .A2(new_n1088), .B1(new_n1091), .B2(new_n1098), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n698), .B1(new_n1099), .B2(KEYINPUT115), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1083), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1076), .A2(new_n692), .B1(new_n1081), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1080), .A2(new_n1103), .ZN(G378));
  NAND2_X1  g0904(.A1(new_n344), .A2(new_n822), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n358), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n358), .A2(new_n1105), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OR3_X1    g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n741), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n693), .B1(new_n1082), .B2(G50), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n780), .A2(new_n578), .B1(new_n721), .B2(new_n701), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G97), .B2(new_n706), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n379), .A2(new_n272), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G283), .B2(new_n710), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n791), .A2(G107), .B1(new_n792), .B2(new_n468), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n717), .A2(G68), .B1(new_n725), .B2(G77), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT58), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1120), .B(new_n249), .C1(G33), .C2(G41), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n706), .A2(G132), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n780), .B2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n791), .A2(G128), .B1(new_n792), .B2(G137), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n724), .B2(new_n1094), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(G150), .C2(new_n717), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n722), .A2(G159), .ZN(new_n1138));
  AOI211_X1 g0938(.A(G33), .B(G41), .C1(new_n710), .C2(G124), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1128), .B1(new_n1125), .B2(new_n1124), .C1(new_n1136), .C2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1117), .B1(new_n1141), .B2(new_n697), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1115), .A2(new_n1142), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT117), .Z(new_n1144));
  INV_X1    g0944(.A(KEYINPUT118), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT40), .B1(new_n858), .B2(new_n853), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1065), .A2(KEYINPUT40), .ZN(new_n1147));
  OAI21_X1  g0947(.A(G330), .B1(new_n818), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1145), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n855), .A2(new_n864), .A3(KEYINPUT118), .A4(G330), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n1150), .A3(new_n1113), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(KEYINPUT118), .A3(new_n1114), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n879), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n879), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1151), .A2(new_n1156), .A3(new_n1153), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1144), .B1(new_n1158), .B2(new_n691), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1057), .B1(new_n1078), .B2(new_n1075), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n1157), .A3(new_n1155), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT57), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n657), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1151), .A2(new_n1156), .A3(new_n1153), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1156), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(KEYINPUT57), .A3(new_n1160), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1159), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(G375));
  NAND2_X1  g0969(.A1(new_n856), .A2(new_n741), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n693), .B1(new_n1082), .B2(G68), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n716), .A2(new_n249), .B1(new_n724), .B2(new_n914), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G132), .B2(new_n719), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n379), .B1(new_n710), .B2(G128), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n791), .A2(G137), .B1(new_n792), .B2(G150), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n706), .A2(new_n1095), .B1(new_n722), .B2(G58), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n707), .A2(new_n578), .B1(new_n721), .B2(new_n203), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n780), .A2(new_n784), .B1(new_n724), .B2(new_n457), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n379), .B1(new_n709), .B2(new_n781), .C1(new_n507), .C2(new_n703), .ZN(new_n1180));
  OR3_X1    g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n716), .A2(new_n422), .B1(new_n700), .B2(new_n902), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT119), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1177), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1171), .B1(new_n1184), .B2(new_n697), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1054), .A2(new_n692), .B1(new_n1170), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1056), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n925), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1186), .B1(new_n1060), .B2(new_n1188), .ZN(G381));
  NAND3_X1  g0989(.A1(new_n974), .A2(new_n755), .A3(new_n1007), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n971), .A2(new_n807), .A3(new_n1191), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1192), .A2(G390), .A3(G381), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT120), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(G375), .A2(G378), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(G407));
  NAND2_X1  g0996(.A1(new_n640), .A2(G213), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(G407), .A2(G213), .A3(new_n1199), .ZN(G409));
  NAND2_X1  g1000(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1159), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(G378), .A3(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1166), .A2(new_n692), .B1(new_n1115), .B2(new_n1142), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1166), .A2(new_n925), .A3(new_n1160), .ZN(new_n1205));
  AOI21_X1  g1005(.A(G378), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1203), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1060), .A2(new_n1187), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT123), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT122), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1187), .A2(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT60), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n657), .B1(new_n1212), .B2(KEYINPUT60), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1209), .A2(new_n1210), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1187), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1078), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT123), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1186), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(G384), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n807), .A3(new_n1186), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1208), .A2(new_n1197), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT62), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT61), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1198), .A2(G2897), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1224), .B(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1206), .B1(new_n1168), .B2(G378), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(new_n1198), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1226), .B(new_n1227), .C1(new_n1229), .C2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT121), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1208), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1203), .A2(KEYINPUT121), .A3(new_n1207), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1234), .A2(new_n1197), .A3(new_n1224), .A4(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(KEYINPUT62), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n755), .B1(new_n974), .B2(new_n1007), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1191), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n969), .B1(new_n954), .B2(new_n691), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1038), .B1(new_n1043), .B2(new_n1044), .C1(new_n1241), .C2(new_n923), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n971), .A2(G390), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1240), .B1(new_n1244), .B2(KEYINPUT127), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT127), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1246), .B(new_n1239), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n1232), .A2(new_n1237), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1208), .A2(KEYINPUT63), .A3(new_n1197), .A4(new_n1224), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1245), .A2(new_n1247), .A3(KEYINPUT61), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1236), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1197), .B1(new_n1230), .B2(KEYINPUT121), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1203), .A2(KEYINPUT121), .A3(new_n1207), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1234), .A2(KEYINPUT125), .A3(new_n1197), .A4(new_n1235), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1229), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1253), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  AOI211_X1 g1061(.A(KEYINPUT126), .B(new_n1229), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1248), .B1(new_n1261), .B2(new_n1262), .ZN(G405));
  NOR2_X1   g1063(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(new_n1224), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1168), .B(G378), .Z(new_n1266));
  XNOR2_X1  g1066(.A(new_n1265), .B(new_n1266), .ZN(G402));
endmodule


