

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U556 ( .A1(n527), .A2(G2104), .ZN(n888) );
  AND2_X2 U557 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  OR2_X2 U558 ( .A1(n750), .A2(n737), .ZN(n743) );
  OR2_X1 U559 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X2 U560 ( .A1(G2104), .A2(n527), .ZN(n891) );
  NOR2_X2 U561 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  INV_X1 U562 ( .A(KEYINPUT90), .ZN(n701) );
  XNOR2_X2 U563 ( .A(KEYINPUT1), .B(n542), .ZN(n590) );
  XOR2_X1 U564 ( .A(KEYINPUT39), .B(n824), .Z(n522) );
  NAND2_X1 U565 ( .A1(n809), .A2(n757), .ZN(n523) );
  NOR2_X1 U566 ( .A1(n738), .A2(n691), .ZN(n693) );
  INV_X1 U567 ( .A(KEYINPUT92), .ZN(n712) );
  INV_X1 U568 ( .A(KEYINPUT95), .ZN(n744) );
  XNOR2_X1 U569 ( .A(KEYINPUT32), .B(KEYINPUT96), .ZN(n747) );
  INV_X1 U570 ( .A(n929), .ZN(n758) );
  NOR2_X1 U571 ( .A1(n815), .A2(n758), .ZN(n759) );
  NAND2_X1 U572 ( .A1(n892), .A2(G114), .ZN(n528) );
  NOR2_X1 U573 ( .A1(G651), .A2(n640), .ZN(n655) );
  NOR2_X2 U574 ( .A1(n541), .A2(n540), .ZN(G160) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n524), .Z(n887) );
  NAND2_X1 U576 ( .A1(G138), .A2(n887), .ZN(n526) );
  INV_X1 U577 ( .A(G2105), .ZN(n527) );
  NAND2_X1 U578 ( .A1(G102), .A2(n888), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n534) );
  NAND2_X1 U580 ( .A1(G126), .A2(n891), .ZN(n530) );
  XNOR2_X1 U581 ( .A(n528), .B(KEYINPUT82), .ZN(n529) );
  NAND2_X1 U582 ( .A1(n530), .A2(n529), .ZN(n532) );
  INV_X1 U583 ( .A(KEYINPUT83), .ZN(n531) );
  XNOR2_X1 U584 ( .A(n532), .B(n531), .ZN(n533) );
  NOR2_X1 U585 ( .A1(n534), .A2(n533), .ZN(G164) );
  NAND2_X1 U586 ( .A1(n887), .A2(G137), .ZN(n537) );
  NAND2_X1 U587 ( .A1(G101), .A2(n888), .ZN(n535) );
  XOR2_X1 U588 ( .A(KEYINPUT23), .B(n535), .Z(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n541) );
  NAND2_X1 U590 ( .A1(G125), .A2(n891), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G113), .A2(n892), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U593 ( .A(KEYINPUT64), .B(G651), .Z(n549) );
  OR2_X1 U594 ( .A1(G543), .A2(n549), .ZN(n542) );
  NAND2_X1 U595 ( .A1(G63), .A2(n590), .ZN(n543) );
  XNOR2_X1 U596 ( .A(KEYINPUT71), .B(n543), .ZN(n546) );
  XOR2_X1 U597 ( .A(G543), .B(KEYINPUT0), .Z(n640) );
  NAND2_X1 U598 ( .A1(n655), .A2(G51), .ZN(n544) );
  XOR2_X1 U599 ( .A(KEYINPUT72), .B(n544), .Z(n545) );
  NOR2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U601 ( .A(n547), .B(KEYINPUT6), .ZN(n554) );
  NOR2_X1 U602 ( .A1(G651), .A2(G543), .ZN(n660) );
  NAND2_X1 U603 ( .A1(n660), .A2(G89), .ZN(n548) );
  XNOR2_X1 U604 ( .A(n548), .B(KEYINPUT4), .ZN(n551) );
  NOR2_X1 U605 ( .A1(n640), .A2(n549), .ZN(n659) );
  NAND2_X1 U606 ( .A1(G76), .A2(n659), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U608 ( .A(KEYINPUT5), .B(n552), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U610 ( .A(n555), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(n660), .A2(G91), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G65), .A2(n590), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n655), .A2(G53), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G78), .A2(n659), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n560) );
  OR2_X1 U618 ( .A1(n561), .A2(n560), .ZN(G299) );
  XOR2_X1 U619 ( .A(G2446), .B(G2430), .Z(n563) );
  XNOR2_X1 U620 ( .A(G2451), .B(G2454), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U622 ( .A(n564), .B(G2427), .Z(n566) );
  XNOR2_X1 U623 ( .A(G1341), .B(G1348), .ZN(n565) );
  XNOR2_X1 U624 ( .A(n566), .B(n565), .ZN(n570) );
  XOR2_X1 U625 ( .A(G2443), .B(KEYINPUT100), .Z(n568) );
  XNOR2_X1 U626 ( .A(G2438), .B(G2435), .ZN(n567) );
  XNOR2_X1 U627 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U628 ( .A(n570), .B(n569), .Z(n571) );
  AND2_X1 U629 ( .A1(G14), .A2(n571), .ZN(G401) );
  AND2_X1 U630 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  INV_X1 U632 ( .A(G132), .ZN(G219) );
  INV_X1 U633 ( .A(G82), .ZN(G220) );
  NAND2_X1 U634 ( .A1(n655), .A2(G52), .ZN(n573) );
  NAND2_X1 U635 ( .A1(G64), .A2(n590), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n579) );
  NAND2_X1 U637 ( .A1(G90), .A2(n660), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G77), .A2(n659), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT66), .B(n576), .Z(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT9), .B(n577), .ZN(n578) );
  NOR2_X1 U642 ( .A1(n579), .A2(n578), .ZN(G171) );
  INV_X1 U643 ( .A(G171), .ZN(G301) );
  NAND2_X1 U644 ( .A1(G88), .A2(n660), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G50), .A2(n655), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U647 ( .A1(G75), .A2(n659), .ZN(n582) );
  XNOR2_X1 U648 ( .A(KEYINPUT79), .B(n582), .ZN(n583) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G62), .A2(n590), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(G303) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n587), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U654 ( .A(G223), .ZN(n836) );
  NAND2_X1 U655 ( .A1(n836), .A2(G567), .ZN(n588) );
  XNOR2_X1 U656 ( .A(n588), .B(KEYINPUT11), .ZN(n589) );
  XNOR2_X1 U657 ( .A(KEYINPUT67), .B(n589), .ZN(G234) );
  NAND2_X1 U658 ( .A1(n590), .A2(G56), .ZN(n591) );
  XOR2_X1 U659 ( .A(KEYINPUT14), .B(n591), .Z(n597) );
  NAND2_X1 U660 ( .A1(n660), .A2(G81), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G68), .A2(n659), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U664 ( .A(KEYINPUT13), .B(n595), .Z(n596) );
  NOR2_X1 U665 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n655), .A2(G43), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n939) );
  INV_X1 U668 ( .A(G860), .ZN(n637) );
  OR2_X1 U669 ( .A1(n939), .A2(n637), .ZN(G153) );
  XNOR2_X1 U670 ( .A(KEYINPUT70), .B(KEYINPUT15), .ZN(n609) );
  NAND2_X1 U671 ( .A1(G92), .A2(n660), .ZN(n600) );
  XNOR2_X1 U672 ( .A(n600), .B(KEYINPUT68), .ZN(n607) );
  NAND2_X1 U673 ( .A1(n655), .A2(G54), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G66), .A2(n590), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U676 ( .A1(G79), .A2(n659), .ZN(n603) );
  XNOR2_X1 U677 ( .A(KEYINPUT69), .B(n603), .ZN(n604) );
  NOR2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n609), .B(n608), .ZN(n936) );
  BUF_X1 U681 ( .A(n936), .Z(n846) );
  INV_X1 U682 ( .A(G868), .ZN(n674) );
  AND2_X1 U683 ( .A1(n846), .A2(n674), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n674), .A2(G301), .ZN(n610) );
  NOR2_X1 U685 ( .A1(n611), .A2(n610), .ZN(G284) );
  NOR2_X1 U686 ( .A1(G868), .A2(G299), .ZN(n613) );
  NOR2_X1 U687 ( .A1(G286), .A2(n674), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U689 ( .A1(n637), .A2(G559), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n614), .A2(n846), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(KEYINPUT73), .ZN(n616) );
  XOR2_X1 U692 ( .A(KEYINPUT16), .B(n616), .Z(G148) );
  NOR2_X1 U693 ( .A1(G868), .A2(n939), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n846), .A2(G868), .ZN(n617) );
  NOR2_X1 U695 ( .A1(G559), .A2(n617), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(G282) );
  XNOR2_X1 U697 ( .A(G2100), .B(KEYINPUT75), .ZN(n629) );
  NAND2_X1 U698 ( .A1(n891), .A2(G123), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT18), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G135), .A2(n887), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U702 ( .A(KEYINPUT74), .B(n623), .ZN(n627) );
  NAND2_X1 U703 ( .A1(G111), .A2(n892), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G99), .A2(n888), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n958) );
  XNOR2_X1 U707 ( .A(n958), .B(G2096), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(G156) );
  NAND2_X1 U709 ( .A1(n660), .A2(G93), .ZN(n631) );
  NAND2_X1 U710 ( .A1(G67), .A2(n590), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n655), .A2(G55), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G80), .A2(n659), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n633), .A2(n632), .ZN(n634) );
  OR2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n673) );
  XNOR2_X1 U716 ( .A(n673), .B(KEYINPUT76), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n846), .A2(G559), .ZN(n636) );
  XOR2_X1 U718 ( .A(n939), .B(n636), .Z(n671) );
  NAND2_X1 U719 ( .A1(n671), .A2(n637), .ZN(n638) );
  XNOR2_X1 U720 ( .A(n639), .B(n638), .ZN(G145) );
  NAND2_X1 U721 ( .A1(G87), .A2(n640), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U724 ( .A1(n590), .A2(n643), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G49), .A2(n655), .ZN(n644) );
  XOR2_X1 U726 ( .A(KEYINPUT77), .B(n644), .Z(n645) );
  NAND2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U728 ( .A(KEYINPUT78), .B(n647), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G86), .A2(n660), .ZN(n649) );
  NAND2_X1 U730 ( .A1(G48), .A2(n655), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n659), .A2(G73), .ZN(n650) );
  XOR2_X1 U733 ( .A(KEYINPUT2), .B(n650), .Z(n651) );
  NOR2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U735 ( .A1(G61), .A2(n590), .ZN(n653) );
  NAND2_X1 U736 ( .A1(n654), .A2(n653), .ZN(G305) );
  NAND2_X1 U737 ( .A1(n655), .A2(G47), .ZN(n657) );
  NAND2_X1 U738 ( .A1(G60), .A2(n590), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U740 ( .A(KEYINPUT65), .B(n658), .ZN(n664) );
  NAND2_X1 U741 ( .A1(n659), .A2(G72), .ZN(n662) );
  NAND2_X1 U742 ( .A1(G85), .A2(n660), .ZN(n661) );
  AND2_X1 U743 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U744 ( .A1(n664), .A2(n663), .ZN(G290) );
  INV_X1 U745 ( .A(G303), .ZN(G166) );
  XOR2_X1 U746 ( .A(n673), .B(G305), .Z(n667) );
  XNOR2_X1 U747 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n665) );
  XNOR2_X1 U748 ( .A(n665), .B(G299), .ZN(n666) );
  XNOR2_X1 U749 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U750 ( .A(G288), .B(n668), .ZN(n670) );
  XNOR2_X1 U751 ( .A(G290), .B(G166), .ZN(n669) );
  XNOR2_X1 U752 ( .A(n670), .B(n669), .ZN(n843) );
  XNOR2_X1 U753 ( .A(n671), .B(n843), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n672), .A2(G868), .ZN(n676) );
  NAND2_X1 U755 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U761 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n681) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n681), .Z(n682) );
  NOR2_X1 U765 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U766 ( .A1(G96), .A2(n683), .ZN(n841) );
  NAND2_X1 U767 ( .A1(n841), .A2(G2106), .ZN(n687) );
  NAND2_X1 U768 ( .A1(G108), .A2(G120), .ZN(n684) );
  NOR2_X1 U769 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U770 ( .A1(G69), .A2(n685), .ZN(n842) );
  NAND2_X1 U771 ( .A1(n842), .A2(G567), .ZN(n686) );
  NAND2_X1 U772 ( .A1(n687), .A2(n686), .ZN(n922) );
  NAND2_X1 U773 ( .A1(G661), .A2(G483), .ZN(n688) );
  XOR2_X1 U774 ( .A(KEYINPUT81), .B(n688), .Z(n689) );
  NOR2_X1 U775 ( .A1(n922), .A2(n689), .ZN(n840) );
  NAND2_X1 U776 ( .A1(n840), .A2(G36), .ZN(G176) );
  NOR2_X2 U777 ( .A1(G164), .A2(G1384), .ZN(n766) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n765) );
  INV_X1 U779 ( .A(n765), .ZN(n690) );
  NAND2_X2 U780 ( .A1(n766), .A2(n690), .ZN(n738) );
  INV_X1 U781 ( .A(G1996), .ZN(n691) );
  XNOR2_X1 U782 ( .A(KEYINPUT26), .B(KEYINPUT89), .ZN(n692) );
  XNOR2_X1 U783 ( .A(n693), .B(n692), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n738), .A2(G1341), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X2 U786 ( .A1(n939), .A2(n696), .ZN(n703) );
  NAND2_X1 U787 ( .A1(n703), .A2(n936), .ZN(n700) );
  INV_X1 U788 ( .A(n738), .ZN(n719) );
  NOR2_X1 U789 ( .A1(n719), .A2(G1348), .ZN(n698) );
  NOR2_X1 U790 ( .A1(G2067), .A2(n738), .ZN(n697) );
  NOR2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n702) );
  XNOR2_X1 U793 ( .A(n702), .B(n701), .ZN(n705) );
  NOR2_X1 U794 ( .A1(n703), .A2(n936), .ZN(n704) );
  NOR2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U796 ( .A(KEYINPUT91), .B(n706), .ZN(n711) );
  NAND2_X1 U797 ( .A1(n719), .A2(G2072), .ZN(n707) );
  XOR2_X1 U798 ( .A(KEYINPUT27), .B(n707), .Z(n709) );
  NAND2_X1 U799 ( .A1(G1956), .A2(n738), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n714) );
  OR2_X1 U801 ( .A1(G299), .A2(n714), .ZN(n710) );
  AND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n713) );
  XNOR2_X1 U803 ( .A(n713), .B(n712), .ZN(n717) );
  NAND2_X1 U804 ( .A1(G299), .A2(n714), .ZN(n715) );
  XNOR2_X1 U805 ( .A(KEYINPUT28), .B(n715), .ZN(n716) );
  NAND2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U807 ( .A(n718), .B(KEYINPUT29), .ZN(n725) );
  NOR2_X1 U808 ( .A1(n719), .A2(G1961), .ZN(n720) );
  XOR2_X1 U809 ( .A(KEYINPUT87), .B(n720), .Z(n723) );
  XOR2_X1 U810 ( .A(G2078), .B(KEYINPUT25), .Z(n721) );
  XNOR2_X1 U811 ( .A(KEYINPUT88), .B(n721), .ZN(n1007) );
  NOR2_X1 U812 ( .A1(n738), .A2(n1007), .ZN(n722) );
  NOR2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n731) );
  NOR2_X1 U814 ( .A1(G301), .A2(n731), .ZN(n724) );
  NOR2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n736) );
  NAND2_X1 U816 ( .A1(G8), .A2(n738), .ZN(n815) );
  NOR2_X1 U817 ( .A1(G1966), .A2(n815), .ZN(n751) );
  NOR2_X1 U818 ( .A1(G2084), .A2(n738), .ZN(n749) );
  NOR2_X1 U819 ( .A1(n751), .A2(n749), .ZN(n726) );
  NAND2_X1 U820 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U821 ( .A(KEYINPUT94), .B(n727), .ZN(n729) );
  XOR2_X1 U822 ( .A(KEYINPUT30), .B(KEYINPUT93), .Z(n728) );
  XNOR2_X1 U823 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U824 ( .A1(G168), .A2(n730), .ZN(n733) );
  AND2_X1 U825 ( .A1(G301), .A2(n731), .ZN(n732) );
  NOR2_X1 U826 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U827 ( .A(n734), .B(KEYINPUT31), .ZN(n735) );
  NOR2_X1 U828 ( .A1(n736), .A2(n735), .ZN(n750) );
  INV_X1 U829 ( .A(G286), .ZN(n737) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n815), .ZN(n740) );
  NOR2_X1 U831 ( .A1(G2090), .A2(n738), .ZN(n739) );
  NOR2_X1 U832 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U833 ( .A1(n741), .A2(G303), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n743), .A2(n742), .ZN(n745) );
  XNOR2_X1 U835 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U836 ( .A1(n746), .A2(G8), .ZN(n748) );
  XNOR2_X1 U837 ( .A(n748), .B(n747), .ZN(n755) );
  NAND2_X1 U838 ( .A1(n749), .A2(G8), .ZN(n753) );
  NOR2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n809) );
  NOR2_X1 U842 ( .A1(G303), .A2(G1971), .ZN(n756) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n932) );
  NOR2_X1 U844 ( .A1(n756), .A2(n932), .ZN(n757) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n929) );
  NAND2_X1 U846 ( .A1(n523), .A2(n759), .ZN(n802) );
  INV_X1 U847 ( .A(KEYINPUT97), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n932), .A2(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n932), .A2(KEYINPUT97), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n815), .A2(n764), .ZN(n799) );
  XOR2_X1 U853 ( .A(G1981), .B(G305), .Z(n923) );
  XNOR2_X1 U854 ( .A(G1986), .B(G290), .ZN(n928) );
  NOR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n827) );
  NAND2_X1 U856 ( .A1(n928), .A2(n827), .ZN(n767) );
  XNOR2_X1 U857 ( .A(n767), .B(KEYINPUT84), .ZN(n786) );
  NAND2_X1 U858 ( .A1(G131), .A2(n887), .ZN(n769) );
  NAND2_X1 U859 ( .A1(G95), .A2(n888), .ZN(n768) );
  NAND2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n773) );
  NAND2_X1 U861 ( .A1(G119), .A2(n891), .ZN(n771) );
  NAND2_X1 U862 ( .A1(G107), .A2(n892), .ZN(n770) );
  NAND2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n900) );
  INV_X1 U865 ( .A(G1991), .ZN(n1002) );
  NOR2_X1 U866 ( .A1(n900), .A2(n1002), .ZN(n783) );
  NAND2_X1 U867 ( .A1(G105), .A2(n888), .ZN(n774) );
  XNOR2_X1 U868 ( .A(n774), .B(KEYINPUT38), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G117), .A2(n892), .ZN(n776) );
  NAND2_X1 U870 ( .A1(G141), .A2(n887), .ZN(n775) );
  NAND2_X1 U871 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U872 ( .A1(n891), .A2(G129), .ZN(n777) );
  XOR2_X1 U873 ( .A(KEYINPUT86), .B(n777), .Z(n778) );
  NOR2_X1 U874 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U875 ( .A1(n781), .A2(n780), .ZN(n904) );
  AND2_X1 U876 ( .A1(n904), .A2(G1996), .ZN(n782) );
  NOR2_X1 U877 ( .A1(n783), .A2(n782), .ZN(n966) );
  INV_X1 U878 ( .A(n827), .ZN(n784) );
  NOR2_X1 U879 ( .A1(n966), .A2(n784), .ZN(n822) );
  INV_X1 U880 ( .A(n822), .ZN(n785) );
  NAND2_X1 U881 ( .A1(n786), .A2(n785), .ZN(n817) );
  INV_X1 U882 ( .A(n817), .ZN(n810) );
  AND2_X1 U883 ( .A1(n923), .A2(n810), .ZN(n797) );
  XNOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NAND2_X1 U885 ( .A1(G140), .A2(n887), .ZN(n788) );
  NAND2_X1 U886 ( .A1(G104), .A2(n888), .ZN(n787) );
  NAND2_X1 U887 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U888 ( .A(KEYINPUT34), .B(n789), .ZN(n794) );
  NAND2_X1 U889 ( .A1(G128), .A2(n891), .ZN(n791) );
  NAND2_X1 U890 ( .A1(G116), .A2(n892), .ZN(n790) );
  NAND2_X1 U891 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U892 ( .A(n792), .B(KEYINPUT35), .Z(n793) );
  NOR2_X1 U893 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U894 ( .A(KEYINPUT36), .B(n795), .Z(n796) );
  XNOR2_X1 U895 ( .A(KEYINPUT85), .B(n796), .ZN(n908) );
  NOR2_X1 U896 ( .A1(n825), .A2(n908), .ZN(n965) );
  NAND2_X1 U897 ( .A1(n965), .A2(n827), .ZN(n831) );
  NAND2_X1 U898 ( .A1(n797), .A2(n831), .ZN(n798) );
  NOR2_X1 U899 ( .A1(n799), .A2(n798), .ZN(n803) );
  INV_X1 U900 ( .A(n803), .ZN(n800) );
  OR2_X1 U901 ( .A1(KEYINPUT97), .A2(n800), .ZN(n801) );
  NOR2_X1 U902 ( .A1(n802), .A2(n801), .ZN(n805) );
  AND2_X1 U903 ( .A1(n803), .A2(KEYINPUT33), .ZN(n804) );
  NOR2_X1 U904 ( .A1(n805), .A2(n804), .ZN(n833) );
  NOR2_X1 U905 ( .A1(G2090), .A2(G303), .ZN(n806) );
  XNOR2_X1 U906 ( .A(n806), .B(KEYINPUT98), .ZN(n807) );
  NAND2_X1 U907 ( .A1(n807), .A2(G8), .ZN(n808) );
  NAND2_X1 U908 ( .A1(n809), .A2(n808), .ZN(n812) );
  AND2_X1 U909 ( .A1(n815), .A2(n810), .ZN(n811) );
  NAND2_X1 U910 ( .A1(n812), .A2(n811), .ZN(n819) );
  NOR2_X1 U911 ( .A1(G1981), .A2(G305), .ZN(n813) );
  XOR2_X1 U912 ( .A(n813), .B(KEYINPUT24), .Z(n814) );
  OR2_X1 U913 ( .A1(n815), .A2(n814), .ZN(n816) );
  OR2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n829) );
  NOR2_X1 U916 ( .A1(G1996), .A2(n904), .ZN(n953) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n820) );
  AND2_X1 U918 ( .A1(n1002), .A2(n900), .ZN(n957) );
  NOR2_X1 U919 ( .A1(n820), .A2(n957), .ZN(n821) );
  NOR2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U921 ( .A1(n953), .A2(n823), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n825), .A2(n908), .ZN(n955) );
  NAND2_X1 U923 ( .A1(n522), .A2(n955), .ZN(n826) );
  AND2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n835) );
  XOR2_X1 U927 ( .A(KEYINPUT99), .B(KEYINPUT40), .Z(n834) );
  XNOR2_X1 U928 ( .A(n835), .B(n834), .ZN(G329) );
  NAND2_X1 U929 ( .A1(n836), .A2(G2106), .ZN(n837) );
  XOR2_X1 U930 ( .A(KEYINPUT101), .B(n837), .Z(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U932 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(G188) );
  XOR2_X1 U935 ( .A(G120), .B(KEYINPUT102), .Z(G236) );
  INV_X1 U937 ( .A(G108), .ZN(G238) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  NOR2_X1 U939 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U941 ( .A(n939), .B(n843), .ZN(n845) );
  XNOR2_X1 U942 ( .A(G286), .B(G171), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n847) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n848) );
  NOR2_X1 U945 ( .A1(G37), .A2(n848), .ZN(G397) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(G2090), .Z(n850) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2084), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n851), .B(G2096), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U952 ( .A(G2100), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT103), .B(G2678), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n857), .B(n856), .Z(G227) );
  XNOR2_X1 U956 ( .A(G1996), .B(KEYINPUT104), .ZN(n867) );
  XOR2_X1 U957 ( .A(G1971), .B(G1956), .Z(n859) );
  XNOR2_X1 U958 ( .A(G1991), .B(G1986), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U960 ( .A(G1976), .B(G1981), .Z(n861) );
  XNOR2_X1 U961 ( .A(G1961), .B(G1966), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U963 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U964 ( .A(KEYINPUT41), .B(G2474), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(G229) );
  NAND2_X1 U967 ( .A1(n891), .A2(G124), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n868), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G112), .A2(n892), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G136), .A2(n887), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G100), .A2(n888), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U974 ( .A1(n874), .A2(n873), .ZN(G162) );
  NAND2_X1 U975 ( .A1(n887), .A2(G142), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n875), .B(KEYINPUT106), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G106), .A2(n888), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n878), .B(KEYINPUT45), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G118), .A2(n892), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G130), .A2(n891), .ZN(n881) );
  XNOR2_X1 U983 ( .A(KEYINPUT105), .B(n881), .ZN(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n912) );
  XOR2_X1 U985 ( .A(KEYINPUT107), .B(KEYINPUT46), .Z(n885) );
  XNOR2_X1 U986 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U988 ( .A(n886), .B(KEYINPUT110), .Z(n902) );
  NAND2_X1 U989 ( .A1(G139), .A2(n887), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G103), .A2(n888), .ZN(n889) );
  NAND2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n898) );
  NAND2_X1 U992 ( .A1(G127), .A2(n891), .ZN(n894) );
  NAND2_X1 U993 ( .A1(G115), .A2(n892), .ZN(n893) );
  NAND2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U995 ( .A(KEYINPUT108), .B(n895), .Z(n896) );
  XNOR2_X1 U996 ( .A(KEYINPUT47), .B(n896), .ZN(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(KEYINPUT109), .B(n899), .Z(n948) );
  XNOR2_X1 U999 ( .A(n900), .B(n948), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(n903), .B(G162), .Z(n906) );
  XOR2_X1 U1002 ( .A(G160), .B(n904), .Z(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n958), .B(n907), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n908), .B(G164), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1007 ( .A(n912), .B(n911), .Z(n913) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(KEYINPUT112), .B(n914), .ZN(G395) );
  NOR2_X1 U1010 ( .A1(G401), .A2(n922), .ZN(n919) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n915) );
  XOR2_X1 U1012 ( .A(KEYINPUT113), .B(n915), .Z(n916) );
  XNOR2_X1 U1013 ( .A(n916), .B(KEYINPUT49), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(G397), .A2(n917), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(n920), .A2(G395), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n921), .B(KEYINPUT114), .ZN(G308) );
  INV_X1 U1018 ( .A(G308), .ZN(G225) );
  INV_X1 U1019 ( .A(n922), .ZN(G319) );
  INV_X1 U1020 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1021 ( .A(G16), .B(KEYINPUT56), .Z(n947) );
  XNOR2_X1 U1022 ( .A(G168), .B(G1966), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n925), .B(KEYINPUT120), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT57), .B(n926), .ZN(n934) );
  XNOR2_X1 U1026 ( .A(G1956), .B(G299), .ZN(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n945) );
  XNOR2_X1 U1031 ( .A(G166), .B(G1971), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(KEYINPUT121), .ZN(n938) );
  XOR2_X1 U1033 ( .A(G1348), .B(n936), .Z(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(G301), .B(G1961), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(n939), .B(G1341), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n1030) );
  INV_X1 U1041 ( .A(KEYINPUT55), .ZN(n1021) );
  XNOR2_X1 U1042 ( .A(KEYINPUT52), .B(KEYINPUT116), .ZN(n971) );
  XOR2_X1 U1043 ( .A(G2072), .B(n948), .Z(n950) );
  XOR2_X1 U1044 ( .A(G164), .B(G2078), .Z(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(KEYINPUT50), .B(n951), .ZN(n963) );
  XOR2_X1 U1047 ( .A(G2090), .B(G162), .Z(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1049 ( .A(KEYINPUT51), .B(n954), .Z(n956) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n961) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(KEYINPUT115), .B(n959), .ZN(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1054 ( .A1(n963), .A2(n962), .ZN(n969) );
  XOR2_X1 U1055 ( .A(G160), .B(G2084), .Z(n964) );
  NOR2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n967) );
  NAND2_X1 U1057 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1058 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1059 ( .A(n971), .B(n970), .ZN(n972) );
  NAND2_X1 U1060 ( .A1(n1021), .A2(n972), .ZN(n973) );
  NAND2_X1 U1061 ( .A1(n973), .A2(G29), .ZN(n1028) );
  XOR2_X1 U1062 ( .A(G4), .B(KEYINPUT123), .Z(n975) );
  XNOR2_X1 U1063 ( .A(G1348), .B(KEYINPUT59), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(n975), .B(n974), .ZN(n979) );
  XNOR2_X1 U1065 ( .A(G1341), .B(G19), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(G1981), .B(G6), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1069 ( .A(KEYINPUT122), .B(G1956), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(G20), .B(n980), .ZN(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(KEYINPUT60), .B(n983), .ZN(n987) );
  XNOR2_X1 U1073 ( .A(G1961), .B(G5), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G21), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n996) );
  XOR2_X1 U1077 ( .A(G1986), .B(G24), .Z(n992) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G22), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(G1976), .B(G23), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n990), .B(KEYINPUT124), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1083 ( .A(KEYINPUT58), .B(n993), .Z(n994) );
  XNOR2_X1 U1084 ( .A(KEYINPUT125), .B(n994), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1086 ( .A(n997), .B(KEYINPUT61), .Z(n998) );
  XNOR2_X1 U1087 ( .A(KEYINPUT126), .B(n998), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(G16), .A2(n999), .ZN(n1026) );
  XNOR2_X1 U1089 ( .A(KEYINPUT117), .B(G2090), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(n1000), .B(G35), .ZN(n1019) );
  XNOR2_X1 U1091 ( .A(G2084), .B(G34), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1001), .B(KEYINPUT54), .ZN(n1017) );
  XNOR2_X1 U1093 ( .A(n1002), .B(G25), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(G28), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(n1004), .B(KEYINPUT118), .ZN(n1013) );
  XNOR2_X1 U1096 ( .A(G1996), .B(G32), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(G33), .B(G2072), .ZN(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1007), .B(G27), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(G26), .B(G2067), .ZN(n1008) );
  NOR2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(KEYINPUT119), .B(n1014), .Z(n1015) );
  XNOR2_X1 U1105 ( .A(KEYINPUT53), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(n1021), .B(n1020), .ZN(n1023) );
  INV_X1 U1109 ( .A(G29), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(G11), .A2(n1024), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT127), .B(n1031), .Z(n1032) );
  XNOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1032), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

