

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783;

  NAND2_X1 U360 ( .A1(n422), .A2(n420), .ZN(n772) );
  AND2_X1 U361 ( .A1(n447), .A2(n445), .ZN(n422) );
  NOR2_X1 U362 ( .A1(n781), .A2(KEYINPUT44), .ZN(n389) );
  NAND2_X1 U363 ( .A1(n375), .A2(n373), .ZN(n783) );
  NAND2_X2 U364 ( .A1(n341), .A2(n398), .ZN(n624) );
  OR2_X1 U365 ( .A1(n685), .A2(n399), .ZN(n398) );
  AND2_X1 U366 ( .A1(n386), .A2(n385), .ZN(n384) );
  XNOR2_X1 U367 ( .A(n340), .B(n474), .ZN(n721) );
  XNOR2_X1 U368 ( .A(n771), .B(G146), .ZN(n340) );
  XNOR2_X1 U369 ( .A(n436), .B(n546), .ZN(n770) );
  XNOR2_X1 U370 ( .A(n469), .B(KEYINPUT64), .ZN(n470) );
  NAND2_X1 U371 ( .A1(n414), .A2(n413), .ZN(n594) );
  AND2_X2 U372 ( .A1(n412), .A2(n415), .ZN(n414) );
  XNOR2_X2 U373 ( .A(n339), .B(n559), .ZN(n561) );
  NAND2_X2 U374 ( .A1(n659), .A2(n639), .ZN(n339) );
  XNOR2_X1 U375 ( .A(n512), .B(n513), .ZN(n515) );
  XNOR2_X2 U376 ( .A(n419), .B(n418), .ZN(n608) );
  OR2_X2 U377 ( .A1(n755), .A2(G902), .ZN(n518) );
  INV_X1 U378 ( .A(n342), .ZN(n341) );
  NAND2_X1 U379 ( .A1(n394), .A2(n396), .ZN(n342) );
  NOR2_X1 U380 ( .A1(n679), .A2(n507), .ZN(n459) );
  XNOR2_X1 U381 ( .A(G104), .B(G113), .ZN(n491) );
  INV_X1 U382 ( .A(G953), .ZN(n773) );
  AND2_X2 U383 ( .A1(n357), .A2(n637), .ZN(n393) );
  NAND2_X2 U384 ( .A1(n616), .A2(n615), .ZN(n358) );
  AND2_X2 U385 ( .A1(n625), .A2(n620), .ZN(n621) );
  XNOR2_X2 U386 ( .A(n358), .B(KEYINPUT106), .ZN(n714) );
  XNOR2_X2 U387 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n469) );
  NOR2_X1 U388 ( .A1(n629), .A2(n697), .ZN(n627) );
  NAND2_X2 U389 ( .A1(n614), .A2(n690), .ZN(n686) );
  AND2_X2 U390 ( .A1(n717), .A2(n715), .ZN(n754) );
  AND2_X1 U391 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U392 ( .A(n440), .B(n439), .ZN(n598) );
  XNOR2_X1 U393 ( .A(n451), .B(n520), .ZN(n540) );
  XNOR2_X1 U394 ( .A(n486), .B(G146), .ZN(n546) );
  XNOR2_X1 U395 ( .A(n452), .B(G116), .ZN(n451) );
  NAND2_X1 U396 ( .A1(n414), .A2(n413), .ZN(n343) );
  BUF_X1 U397 ( .A(n619), .Z(n629) );
  XNOR2_X2 U398 ( .A(n528), .B(n473), .ZN(n771) );
  XNOR2_X2 U399 ( .A(n543), .B(n472), .ZN(n528) );
  XOR2_X1 U400 ( .A(G137), .B(G134), .Z(n471) );
  OR2_X1 U401 ( .A1(n609), .A2(n737), .ZN(n450) );
  INV_X1 U402 ( .A(G125), .ZN(n486) );
  XNOR2_X1 U403 ( .A(n498), .B(n644), .ZN(n441) );
  INV_X1 U404 ( .A(KEYINPUT1), .ZN(n443) );
  OR2_X1 U405 ( .A1(n435), .A2(n668), .ZN(n434) );
  INV_X1 U406 ( .A(n384), .ZN(n380) );
  NAND2_X1 U407 ( .A1(n377), .A2(n354), .ZN(n376) );
  NAND2_X1 U408 ( .A1(n381), .A2(n378), .ZN(n377) );
  INV_X1 U409 ( .A(n598), .ZN(n378) );
  OR2_X1 U410 ( .A1(n534), .A2(n408), .ZN(n601) );
  BUF_X1 U411 ( .A(n561), .Z(n605) );
  NOR2_X1 U412 ( .A1(G237), .A2(G953), .ZN(n492) );
  INV_X1 U413 ( .A(n772), .ZN(n456) );
  INV_X1 U414 ( .A(n579), .ZN(n580) );
  NAND2_X1 U415 ( .A1(n363), .A2(n360), .ZN(n366) );
  AND2_X1 U416 ( .A1(n364), .A2(n365), .ZN(n363) );
  NAND2_X1 U417 ( .A1(n686), .A2(KEYINPUT109), .ZN(n364) );
  NAND2_X1 U418 ( .A1(n453), .A2(KEYINPUT22), .ZN(n406) );
  XNOR2_X1 U419 ( .A(n518), .B(n458), .ZN(n575) );
  XNOR2_X1 U420 ( .A(G110), .B(G119), .ZN(n509) );
  XOR2_X1 U421 ( .A(G137), .B(G128), .Z(n510) );
  XNOR2_X1 U422 ( .A(n427), .B(n425), .ZN(n514) );
  XNOR2_X1 U423 ( .A(KEYINPUT78), .B(KEYINPUT8), .ZN(n427) );
  NOR2_X1 U424 ( .A1(n426), .A2(G953), .ZN(n425) );
  INV_X1 U425 ( .A(G234), .ZN(n426) );
  XNOR2_X1 U426 ( .A(G107), .B(G116), .ZN(n479) );
  INV_X1 U427 ( .A(KEYINPUT9), .ZN(n478) );
  XNOR2_X1 U428 ( .A(KEYINPUT7), .B(G134), .ZN(n432) );
  XNOR2_X1 U429 ( .A(G122), .B(KEYINPUT100), .ZN(n476) );
  XOR2_X1 U430 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n477) );
  XOR2_X1 U431 ( .A(G143), .B(G122), .Z(n490) );
  XNOR2_X1 U432 ( .A(n487), .B(G140), .ZN(n436) );
  XOR2_X1 U433 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n487) );
  XNOR2_X1 U434 ( .A(G131), .B(KEYINPUT12), .ZN(n488) );
  XOR2_X1 U435 ( .A(KEYINPUT11), .B(KEYINPUT96), .Z(n489) );
  NAND2_X1 U436 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U437 ( .A1(n400), .A2(n401), .ZN(n399) );
  AND2_X1 U438 ( .A1(n397), .A2(n623), .ZN(n396) );
  NAND2_X1 U439 ( .A1(n629), .A2(KEYINPUT34), .ZN(n397) );
  XNOR2_X1 U440 ( .A(n531), .B(n530), .ZN(n693) );
  INV_X1 U441 ( .A(KEYINPUT103), .ZN(n439) );
  INV_X1 U442 ( .A(n586), .ZN(n362) );
  NAND2_X1 U443 ( .A1(n674), .A2(n372), .ZN(n371) );
  NOR2_X1 U444 ( .A1(n344), .A2(n351), .ZN(n372) );
  INV_X1 U445 ( .A(n707), .ZN(n368) );
  NAND2_X1 U446 ( .A1(n438), .A2(n442), .ZN(n437) );
  XNOR2_X1 U447 ( .A(n602), .B(KEYINPUT36), .ZN(n438) );
  INV_X1 U448 ( .A(n639), .ZN(n457) );
  XNOR2_X1 U449 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n545) );
  NAND2_X1 U450 ( .A1(G234), .A2(G237), .ZN(n502) );
  INV_X1 U451 ( .A(G237), .ZN(n535) );
  NAND2_X1 U452 ( .A1(n586), .A2(KEYINPUT109), .ZN(n365) );
  XNOR2_X1 U453 ( .A(n499), .B(n536), .ZN(n639) );
  XNOR2_X1 U454 ( .A(KEYINPUT83), .B(KEYINPUT15), .ZN(n499) );
  NAND2_X1 U455 ( .A1(n455), .A2(n569), .ZN(n453) );
  NAND2_X1 U456 ( .A1(n721), .A2(n536), .ZN(n433) );
  XOR2_X1 U457 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n522) );
  XNOR2_X1 U458 ( .A(G101), .B(G146), .ZN(n521) );
  XNOR2_X1 U459 ( .A(KEYINPUT16), .B(G122), .ZN(n539) );
  NAND2_X1 U460 ( .A1(n604), .A2(n428), .ZN(n679) );
  INV_X1 U461 ( .A(n741), .ZN(n409) );
  NAND2_X1 U462 ( .A1(n588), .A2(KEYINPUT19), .ZN(n415) );
  NAND2_X1 U463 ( .A1(n421), .A2(n448), .ZN(n420) );
  NOR2_X1 U464 ( .A1(n450), .A2(KEYINPUT48), .ZN(n448) );
  INV_X1 U465 ( .A(KEYINPUT73), .ZN(n418) );
  NAND2_X1 U466 ( .A1(n366), .A2(n582), .ZN(n419) );
  XOR2_X1 U467 ( .A(KEYINPUT62), .B(n653), .Z(n654) );
  XNOR2_X1 U468 ( .A(n515), .B(n460), .ZN(n755) );
  XNOR2_X1 U469 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U470 ( .A(n770), .B(n347), .ZN(n496) );
  XNOR2_X1 U471 ( .A(n661), .B(n660), .ZN(n662) );
  OR2_X1 U472 ( .A1(n601), .A2(n442), .ZN(n538) );
  NAND2_X1 U473 ( .A1(n353), .A2(n384), .ZN(n373) );
  AND2_X1 U474 ( .A1(n379), .A2(n376), .ZN(n375) );
  XNOR2_X1 U475 ( .A(n573), .B(n572), .ZN(n617) );
  NAND2_X1 U476 ( .A1(n442), .A2(n575), .ZN(n571) );
  XOR2_X1 U477 ( .A(n598), .B(KEYINPUT107), .Z(n741) );
  NAND2_X1 U478 ( .A1(n346), .A2(n628), .ZN(n630) );
  INV_X1 U479 ( .A(KEYINPUT123), .ZN(n417) );
  NAND2_X1 U480 ( .A1(n370), .A2(n367), .ZN(n713) );
  NAND2_X1 U481 ( .A1(n369), .A2(n352), .ZN(n367) );
  NAND2_X1 U482 ( .A1(n371), .A2(KEYINPUT119), .ZN(n370) );
  INV_X1 U483 ( .A(n437), .ZN(n748) );
  AND2_X1 U484 ( .A1(n709), .A2(n704), .ZN(n344) );
  NOR2_X1 U485 ( .A1(n641), .A2(n356), .ZN(n345) );
  AND2_X1 U486 ( .A1(n362), .A2(n359), .ZN(n346) );
  XNOR2_X1 U487 ( .A(n497), .B(n441), .ZN(n596) );
  XOR2_X1 U488 ( .A(n489), .B(n488), .Z(n347) );
  AND2_X1 U489 ( .A1(n516), .A2(G217), .ZN(n348) );
  XOR2_X1 U490 ( .A(G107), .B(G110), .Z(n349) );
  OR2_X1 U491 ( .A1(n588), .A2(KEYINPUT19), .ZN(n350) );
  NOR2_X1 U492 ( .A1(G953), .A2(n707), .ZN(n351) );
  NOR2_X1 U493 ( .A1(n712), .A2(n368), .ZN(n352) );
  AND2_X1 U494 ( .A1(n381), .A2(n374), .ZN(n353) );
  INV_X1 U495 ( .A(n575), .ZN(n614) );
  XOR2_X1 U496 ( .A(KEYINPUT40), .B(KEYINPUT111), .Z(n354) );
  INV_X1 U497 ( .A(KEYINPUT34), .ZN(n401) );
  AND2_X1 U498 ( .A1(KEYINPUT66), .A2(KEYINPUT2), .ZN(n355) );
  AND2_X1 U499 ( .A1(n457), .A2(n355), .ZN(n356) );
  NAND2_X1 U500 ( .A1(n404), .A2(n403), .ZN(n613) );
  NAND2_X1 U501 ( .A1(n405), .A2(n407), .ZN(n404) );
  NAND2_X1 U502 ( .A1(n388), .A2(n389), .ZN(n357) );
  INV_X1 U503 ( .A(n686), .ZN(n359) );
  NAND2_X1 U504 ( .A1(n362), .A2(n361), .ZN(n360) );
  NOR2_X1 U505 ( .A1(n686), .A2(KEYINPUT109), .ZN(n361) );
  NAND2_X1 U506 ( .A1(n706), .A2(n705), .ZN(n369) );
  NAND2_X1 U507 ( .A1(n384), .A2(n381), .ZN(n610) );
  NOR2_X1 U508 ( .A1(n598), .A2(n354), .ZN(n374) );
  NAND2_X1 U509 ( .A1(n380), .A2(n354), .ZN(n379) );
  NOR2_X1 U510 ( .A1(n675), .A2(n387), .ZN(n382) );
  INV_X1 U511 ( .A(n608), .ZN(n383) );
  NAND2_X1 U512 ( .A1(n675), .A2(n387), .ZN(n385) );
  NAND2_X1 U513 ( .A1(n608), .A2(n387), .ZN(n386) );
  INV_X1 U514 ( .A(KEYINPUT39), .ZN(n387) );
  INV_X1 U515 ( .A(n402), .ZN(n388) );
  NAND2_X1 U516 ( .A1(n393), .A2(n390), .ZN(n638) );
  NAND2_X1 U517 ( .A1(n781), .A2(KEYINPUT44), .ZN(n391) );
  NAND2_X1 U518 ( .A1(n402), .A2(KEYINPUT44), .ZN(n392) );
  NAND2_X1 U519 ( .A1(n685), .A2(KEYINPUT34), .ZN(n394) );
  INV_X1 U520 ( .A(n629), .ZN(n400) );
  XNOR2_X2 U521 ( .A(n621), .B(KEYINPUT33), .ZN(n685) );
  XNOR2_X1 U522 ( .A(n618), .B(KEYINPUT80), .ZN(n402) );
  XNOR2_X2 U523 ( .A(n624), .B(KEYINPUT35), .ZN(n781) );
  NAND2_X1 U524 ( .A1(n619), .A2(n406), .ZN(n403) );
  INV_X1 U525 ( .A(n619), .ZN(n405) );
  NAND2_X1 U526 ( .A1(n453), .A2(n454), .ZN(n407) );
  AND2_X1 U527 ( .A1(n446), .A2(n612), .ZN(n445) );
  NAND2_X1 U528 ( .A1(n437), .A2(n603), .ZN(n609) );
  NAND2_X1 U529 ( .A1(n409), .A2(n676), .ZN(n408) );
  XNOR2_X1 U530 ( .A(n725), .B(n417), .ZN(G54) );
  XNOR2_X1 U531 ( .A(n410), .B(KEYINPUT105), .ZN(n616) );
  NAND2_X1 U532 ( .A1(n554), .A2(n555), .ZN(n659) );
  NAND2_X1 U533 ( .A1(n613), .A2(n687), .ZN(n410) );
  XNOR2_X1 U534 ( .A(n541), .B(n542), .ZN(n551) );
  NAND2_X1 U535 ( .A1(n754), .A2(G472), .ZN(n655) );
  NAND2_X2 U536 ( .A1(n424), .A2(n345), .ZN(n717) );
  NAND2_X1 U537 ( .A1(n561), .A2(KEYINPUT19), .ZN(n412) );
  OR2_X1 U538 ( .A1(n561), .A2(n350), .ZN(n413) );
  XNOR2_X2 U539 ( .A(n416), .B(n568), .ZN(n619) );
  NAND2_X1 U540 ( .A1(n594), .A2(n566), .ZN(n416) );
  INV_X1 U541 ( .A(n449), .ZN(n421) );
  AND2_X2 U542 ( .A1(n642), .A2(n457), .ZN(n423) );
  XNOR2_X2 U543 ( .A(n638), .B(KEYINPUT45), .ZN(n642) );
  NAND2_X1 U544 ( .A1(n456), .A2(n423), .ZN(n424) );
  INV_X1 U545 ( .A(n604), .ZN(n597) );
  INV_X1 U546 ( .A(n596), .ZN(n428) );
  NOR2_X1 U547 ( .A1(n751), .A2(G902), .ZN(n484) );
  XNOR2_X1 U548 ( .A(n430), .B(n429), .ZN(n751) );
  XNOR2_X1 U549 ( .A(n481), .B(n480), .ZN(n429) );
  XNOR2_X1 U550 ( .A(n482), .B(n431), .ZN(n430) );
  XNOR2_X1 U551 ( .A(n483), .B(n432), .ZN(n431) );
  NOR2_X1 U552 ( .A1(n687), .A2(n686), .ZN(n625) );
  XNOR2_X2 U553 ( .A(n576), .B(n443), .ZN(n687) );
  XNOR2_X2 U554 ( .A(n433), .B(G469), .ZN(n576) );
  NAND2_X1 U555 ( .A1(n434), .A2(n671), .ZN(n706) );
  NAND2_X1 U556 ( .A1(n642), .A2(n667), .ZN(n435) );
  NAND2_X1 U557 ( .A1(n604), .A2(n596), .ZN(n440) );
  NAND2_X1 U558 ( .A1(n754), .A2(G210), .ZN(n663) );
  AND2_X1 U559 ( .A1(n687), .A2(n614), .ZN(n634) );
  INV_X1 U560 ( .A(n687), .ZN(n442) );
  XNOR2_X1 U561 ( .A(n593), .B(KEYINPUT46), .ZN(n449) );
  NAND2_X1 U562 ( .A1(n450), .A2(KEYINPUT48), .ZN(n446) );
  NAND2_X1 U563 ( .A1(n449), .A2(KEYINPUT48), .ZN(n447) );
  XNOR2_X1 U564 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X2 U565 ( .A(G113), .B(KEYINPUT85), .ZN(n452) );
  NAND2_X1 U566 ( .A1(n459), .A2(KEYINPUT22), .ZN(n454) );
  INV_X1 U567 ( .A(n459), .ZN(n455) );
  INV_X1 U568 ( .A(n642), .ZN(n669) );
  BUF_X1 U569 ( .A(n659), .Z(n661) );
  XNOR2_X2 U570 ( .A(n483), .B(n470), .ZN(n543) );
  XOR2_X1 U571 ( .A(n517), .B(n348), .Z(n458) );
  AND2_X1 U572 ( .A1(n514), .A2(G221), .ZN(n460) );
  XNOR2_X1 U573 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U574 ( .A(n542), .B(n465), .ZN(n466) );
  INV_X1 U575 ( .A(KEYINPUT90), .ZN(n473) );
  AND2_X1 U576 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U577 ( .A(G104), .B(G101), .ZN(n461) );
  XNOR2_X1 U578 ( .A(n349), .B(n461), .ZN(n462) );
  XOR2_X1 U579 ( .A(KEYINPUT84), .B(n462), .Z(n542) );
  NAND2_X1 U580 ( .A1(G227), .A2(n773), .ZN(n464) );
  INV_X1 U581 ( .A(KEYINPUT74), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n466), .B(G140), .ZN(n474) );
  XNOR2_X2 U583 ( .A(G143), .B(KEYINPUT76), .ZN(n468) );
  INV_X1 U584 ( .A(G128), .ZN(n467) );
  XNOR2_X2 U585 ( .A(n468), .B(n467), .ZN(n483) );
  XNOR2_X1 U586 ( .A(n471), .B(G131), .ZN(n472) );
  INV_X1 U587 ( .A(G902), .ZN(n536) );
  XOR2_X1 U588 ( .A(G478), .B(KEYINPUT102), .Z(n475) );
  XNOR2_X1 U589 ( .A(KEYINPUT101), .B(n475), .ZN(n485) );
  XNOR2_X1 U590 ( .A(n477), .B(n476), .ZN(n481) );
  NAND2_X1 U591 ( .A1(G217), .A2(n514), .ZN(n482) );
  XNOR2_X1 U592 ( .A(n485), .B(n484), .ZN(n604) );
  XNOR2_X1 U593 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n498) );
  XNOR2_X1 U594 ( .A(n491), .B(n490), .ZN(n494) );
  XNOR2_X1 U595 ( .A(n492), .B(KEYINPUT72), .ZN(n523) );
  NAND2_X1 U596 ( .A1(G214), .A2(n523), .ZN(n493) );
  XOR2_X1 U597 ( .A(n494), .B(n493), .Z(n495) );
  XNOR2_X1 U598 ( .A(n496), .B(n495), .ZN(n647) );
  NOR2_X1 U599 ( .A1(G902), .A2(n647), .ZN(n497) );
  INV_X1 U600 ( .A(G475), .ZN(n644) );
  NAND2_X1 U601 ( .A1(n639), .A2(G234), .ZN(n500) );
  XNOR2_X1 U602 ( .A(n500), .B(KEYINPUT20), .ZN(n516) );
  AND2_X1 U603 ( .A1(n516), .A2(G221), .ZN(n501) );
  XNOR2_X1 U604 ( .A(n501), .B(KEYINPUT21), .ZN(n690) );
  INV_X1 U605 ( .A(n690), .ZN(n507) );
  XOR2_X1 U606 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n503) );
  XNOR2_X1 U607 ( .A(n503), .B(n502), .ZN(n504) );
  AND2_X1 U608 ( .A1(n504), .A2(G952), .ZN(n708) );
  AND2_X1 U609 ( .A1(n708), .A2(n773), .ZN(n704) );
  NAND2_X1 U610 ( .A1(G902), .A2(n504), .ZN(n563) );
  OR2_X1 U611 ( .A1(n773), .A2(n563), .ZN(n505) );
  NOR2_X1 U612 ( .A1(G900), .A2(n505), .ZN(n506) );
  NOR2_X1 U613 ( .A1(n704), .A2(n506), .ZN(n579) );
  NOR2_X1 U614 ( .A1(n507), .A2(n579), .ZN(n508) );
  XNOR2_X1 U615 ( .A(KEYINPUT70), .B(n508), .ZN(n519) );
  XNOR2_X1 U616 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U617 ( .A(n511), .B(KEYINPUT23), .Z(n513) );
  XNOR2_X1 U618 ( .A(n770), .B(KEYINPUT24), .ZN(n512) );
  XOR2_X1 U619 ( .A(KEYINPUT91), .B(KEYINPUT25), .Z(n517) );
  NAND2_X1 U620 ( .A1(n519), .A2(n575), .ZN(n584) );
  XOR2_X1 U621 ( .A(KEYINPUT3), .B(G119), .Z(n520) );
  XNOR2_X1 U622 ( .A(n522), .B(n521), .ZN(n525) );
  NAND2_X1 U623 ( .A1(G210), .A2(n523), .ZN(n524) );
  XNOR2_X1 U624 ( .A(n524), .B(n525), .ZN(n526) );
  XNOR2_X1 U625 ( .A(n540), .B(n526), .ZN(n527) );
  XNOR2_X1 U626 ( .A(n528), .B(n527), .ZN(n653) );
  NAND2_X1 U627 ( .A1(n653), .A2(n536), .ZN(n531) );
  INV_X1 U628 ( .A(KEYINPUT93), .ZN(n529) );
  XNOR2_X1 U629 ( .A(n529), .B(G472), .ZN(n530) );
  INV_X1 U630 ( .A(KEYINPUT6), .ZN(n532) );
  XNOR2_X1 U631 ( .A(n693), .B(n532), .ZN(n620) );
  INV_X1 U632 ( .A(n620), .ZN(n570) );
  NOR2_X1 U633 ( .A1(n584), .A2(n570), .ZN(n533) );
  XOR2_X1 U634 ( .A(KEYINPUT108), .B(n533), .Z(n534) );
  NAND2_X1 U635 ( .A1(n536), .A2(n535), .ZN(n556) );
  NAND2_X1 U636 ( .A1(n556), .A2(G214), .ZN(n537) );
  XNOR2_X1 U637 ( .A(n537), .B(KEYINPUT88), .ZN(n676) );
  XNOR2_X1 U638 ( .A(n538), .B(KEYINPUT43), .ZN(n560) );
  INV_X1 U639 ( .A(n543), .ZN(n550) );
  NAND2_X1 U640 ( .A1(n773), .A2(G224), .ZN(n544) );
  XNOR2_X1 U641 ( .A(n544), .B(KEYINPUT86), .ZN(n548) );
  XNOR2_X1 U642 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U643 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U644 ( .A(n550), .B(n549), .ZN(n552) );
  NAND2_X1 U645 ( .A1(n551), .A2(n552), .ZN(n555) );
  INV_X1 U646 ( .A(n551), .ZN(n759) );
  INV_X1 U647 ( .A(n552), .ZN(n553) );
  NAND2_X1 U648 ( .A1(n759), .A2(n553), .ZN(n554) );
  NAND2_X1 U649 ( .A1(n556), .A2(G210), .ZN(n558) );
  INV_X1 U650 ( .A(KEYINPUT87), .ZN(n557) );
  XNOR2_X1 U651 ( .A(n558), .B(n557), .ZN(n559) );
  AND2_X1 U652 ( .A1(n560), .A2(n605), .ZN(n611) );
  XOR2_X1 U653 ( .A(n611), .B(G140), .Z(G42) );
  XNOR2_X1 U654 ( .A(G119), .B(KEYINPUT127), .ZN(n574) );
  INV_X1 U655 ( .A(n676), .ZN(n588) );
  INV_X1 U656 ( .A(n704), .ZN(n565) );
  NOR2_X1 U657 ( .A1(G898), .A2(n773), .ZN(n562) );
  XNOR2_X1 U658 ( .A(KEYINPUT89), .B(n562), .ZN(n761) );
  OR2_X1 U659 ( .A1(n761), .A2(n563), .ZN(n564) );
  NAND2_X1 U660 ( .A1(n565), .A2(n564), .ZN(n566) );
  INV_X1 U661 ( .A(KEYINPUT67), .ZN(n567) );
  XNOR2_X1 U662 ( .A(n567), .B(KEYINPUT0), .ZN(n568) );
  INV_X1 U663 ( .A(KEYINPUT22), .ZN(n569) );
  NAND2_X1 U664 ( .A1(n613), .A2(n570), .ZN(n633) );
  NOR2_X1 U665 ( .A1(n633), .A2(n571), .ZN(n573) );
  XNOR2_X1 U666 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n572) );
  XOR2_X1 U667 ( .A(n574), .B(n617), .Z(G21) );
  INV_X1 U668 ( .A(n576), .ZN(n586) );
  XOR2_X1 U669 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n578) );
  NAND2_X1 U670 ( .A1(n693), .A2(n676), .ZN(n577) );
  XNOR2_X1 U671 ( .A(n578), .B(n577), .ZN(n581) );
  INV_X1 U672 ( .A(KEYINPUT38), .ZN(n583) );
  XNOR2_X1 U673 ( .A(n605), .B(n583), .ZN(n675) );
  INV_X1 U674 ( .A(n693), .ZN(n628) );
  NOR2_X1 U675 ( .A1(n584), .A2(n628), .ZN(n585) );
  XOR2_X1 U676 ( .A(KEYINPUT28), .B(n585), .Z(n587) );
  NOR2_X1 U677 ( .A1(n587), .A2(n586), .ZN(n595) );
  OR2_X1 U678 ( .A1(n675), .A2(n588), .ZN(n680) );
  OR2_X1 U679 ( .A1(n680), .A2(n679), .ZN(n590) );
  INV_X1 U680 ( .A(KEYINPUT41), .ZN(n589) );
  XNOR2_X1 U681 ( .A(n590), .B(n589), .ZN(n699) );
  INV_X1 U682 ( .A(n699), .ZN(n591) );
  NAND2_X1 U683 ( .A1(n595), .A2(n591), .ZN(n592) );
  XNOR2_X1 U684 ( .A(KEYINPUT42), .B(n592), .ZN(n782) );
  NAND2_X1 U685 ( .A1(n783), .A2(n782), .ZN(n593) );
  NAND2_X1 U686 ( .A1(n595), .A2(n343), .ZN(n738) );
  NAND2_X1 U687 ( .A1(n428), .A2(n597), .ZN(n744) );
  AND2_X1 U688 ( .A1(n744), .A2(n598), .ZN(n599) );
  XNOR2_X1 U689 ( .A(n599), .B(KEYINPUT104), .ZN(n681) );
  NOR2_X1 U690 ( .A1(n738), .A2(n681), .ZN(n600) );
  XNOR2_X1 U691 ( .A(n600), .B(KEYINPUT47), .ZN(n603) );
  NOR2_X1 U692 ( .A1(n601), .A2(n605), .ZN(n602) );
  NOR2_X1 U693 ( .A1(n428), .A2(n604), .ZN(n622) );
  INV_X1 U694 ( .A(n605), .ZN(n606) );
  NAND2_X1 U695 ( .A1(n622), .A2(n606), .ZN(n607) );
  NOR2_X1 U696 ( .A1(n608), .A2(n607), .ZN(n737) );
  NOR2_X1 U697 ( .A1(n610), .A2(n744), .ZN(n750) );
  NOR2_X1 U698 ( .A1(n750), .A2(n611), .ZN(n612) );
  NOR2_X1 U699 ( .A1(n614), .A2(n693), .ZN(n615) );
  NAND2_X1 U700 ( .A1(n714), .A2(n617), .ZN(n618) );
  XOR2_X1 U701 ( .A(n622), .B(KEYINPUT75), .Z(n623) );
  NAND2_X1 U702 ( .A1(n693), .A2(n625), .ZN(n697) );
  XNOR2_X1 U703 ( .A(KEYINPUT31), .B(KEYINPUT94), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n627), .B(n626), .ZN(n745) );
  OR2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n730) );
  NAND2_X1 U706 ( .A1(n745), .A2(n730), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT95), .ZN(n632) );
  NOR2_X1 U708 ( .A1(n632), .A2(n681), .ZN(n636) );
  INV_X1 U709 ( .A(n633), .ZN(n635) );
  AND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n726) );
  NOR2_X1 U711 ( .A1(n636), .A2(n726), .ZN(n637) );
  INV_X1 U712 ( .A(KEYINPUT2), .ZN(n643) );
  NOR2_X1 U713 ( .A1(n639), .A2(n643), .ZN(n640) );
  NOR2_X1 U714 ( .A1(n640), .A2(KEYINPUT66), .ZN(n641) );
  NOR2_X1 U715 ( .A1(n772), .A2(n643), .ZN(n668) );
  NAND2_X1 U716 ( .A1(n642), .A2(n668), .ZN(n715) );
  NAND2_X1 U717 ( .A1(n717), .A2(n715), .ZN(n645) );
  NOR2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n649) );
  XNOR2_X1 U719 ( .A(KEYINPUT82), .B(KEYINPUT59), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n649), .B(n648), .ZN(n651) );
  INV_X1 U722 ( .A(G952), .ZN(n650) );
  AND2_X1 U723 ( .A1(n650), .A2(G953), .ZN(n758) );
  NOR2_X1 U724 ( .A1(n651), .A2(n758), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U726 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X2 U727 ( .A1(n656), .A2(n758), .ZN(n658) );
  XNOR2_X1 U728 ( .A(KEYINPUT81), .B(KEYINPUT63), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n658), .B(n657), .ZN(G57) );
  XNOR2_X1 U730 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X2 U732 ( .A1(n664), .A2(n758), .ZN(n666) );
  XNOR2_X1 U733 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n665) );
  XNOR2_X1 U734 ( .A(n666), .B(n665), .ZN(G51) );
  INV_X1 U735 ( .A(KEYINPUT79), .ZN(n667) );
  XNOR2_X1 U736 ( .A(KEYINPUT2), .B(KEYINPUT77), .ZN(n672) );
  XNOR2_X1 U737 ( .A(n672), .B(KEYINPUT79), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n669), .A2(n670), .ZN(n671) );
  NAND2_X1 U739 ( .A1(n772), .A2(n672), .ZN(n705) );
  AND2_X1 U740 ( .A1(n705), .A2(n773), .ZN(n673) );
  NAND2_X1 U741 ( .A1(n706), .A2(n673), .ZN(n674) );
  OR2_X1 U742 ( .A1(n699), .A2(n685), .ZN(n707) );
  INV_X1 U743 ( .A(n675), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n683) );
  NOR2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n702) );
  NAND2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n689) );
  XNOR2_X1 U750 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n688) );
  XNOR2_X1 U751 ( .A(n689), .B(n688), .ZN(n695) );
  NOR2_X1 U752 ( .A1(n614), .A2(n690), .ZN(n691) );
  XOR2_X1 U753 ( .A(KEYINPUT49), .B(n691), .Z(n692) );
  NOR2_X1 U754 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U755 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U756 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U757 ( .A(KEYINPUT51), .B(n698), .ZN(n700) );
  NOR2_X1 U758 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U759 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U760 ( .A(n703), .B(KEYINPUT52), .Z(n709) );
  NAND2_X1 U761 ( .A1(n709), .A2(n708), .ZN(n711) );
  NOR2_X1 U762 ( .A1(G953), .A2(KEYINPUT119), .ZN(n710) );
  NAND2_X1 U763 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U764 ( .A(n713), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U765 ( .A(n714), .B(G110), .ZN(G12) );
  AND2_X1 U766 ( .A1(n715), .A2(G469), .ZN(n716) );
  NAND2_X1 U767 ( .A1(n717), .A2(n716), .ZN(n723) );
  XOR2_X1 U768 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n719) );
  XNOR2_X1 U769 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n718) );
  XNOR2_X1 U770 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U772 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U773 ( .A1(n724), .A2(n758), .ZN(n725) );
  XOR2_X1 U774 ( .A(G101), .B(n726), .Z(G3) );
  NOR2_X1 U775 ( .A1(n741), .A2(n730), .ZN(n728) );
  XNOR2_X1 U776 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n727) );
  XNOR2_X1 U777 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U778 ( .A(G104), .B(n729), .ZN(G6) );
  NOR2_X1 U779 ( .A1(n744), .A2(n730), .ZN(n732) );
  XNOR2_X1 U780 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X1 U782 ( .A(G107), .B(n733), .ZN(G9) );
  NOR2_X1 U783 ( .A1(n738), .A2(n744), .ZN(n735) );
  XNOR2_X1 U784 ( .A(KEYINPUT29), .B(KEYINPUT114), .ZN(n734) );
  XNOR2_X1 U785 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U786 ( .A(G128), .B(n736), .ZN(G30) );
  XOR2_X1 U787 ( .A(G143), .B(n737), .Z(G45) );
  NOR2_X1 U788 ( .A1(n741), .A2(n738), .ZN(n740) );
  XNOR2_X1 U789 ( .A(G146), .B(KEYINPUT115), .ZN(n739) );
  XNOR2_X1 U790 ( .A(n740), .B(n739), .ZN(G48) );
  NOR2_X1 U791 ( .A1(n745), .A2(n741), .ZN(n742) );
  XOR2_X1 U792 ( .A(KEYINPUT116), .B(n742), .Z(n743) );
  XNOR2_X1 U793 ( .A(G113), .B(n743), .ZN(G15) );
  NOR2_X1 U794 ( .A1(n745), .A2(n744), .ZN(n747) );
  XNOR2_X1 U795 ( .A(G116), .B(KEYINPUT117), .ZN(n746) );
  XNOR2_X1 U796 ( .A(n747), .B(n746), .ZN(G18) );
  XNOR2_X1 U797 ( .A(G125), .B(n748), .ZN(n749) );
  XNOR2_X1 U798 ( .A(n749), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U799 ( .A(G134), .B(n750), .Z(G36) );
  NAND2_X1 U800 ( .A1(n754), .A2(G478), .ZN(n752) );
  XNOR2_X1 U801 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U802 ( .A1(n758), .A2(n753), .ZN(G63) );
  NAND2_X1 U803 ( .A1(n754), .A2(G217), .ZN(n756) );
  XNOR2_X1 U804 ( .A(n756), .B(n755), .ZN(n757) );
  NOR2_X1 U805 ( .A1(n758), .A2(n757), .ZN(G66) );
  INV_X1 U806 ( .A(n759), .ZN(n760) );
  XNOR2_X1 U807 ( .A(n760), .B(KEYINPUT125), .ZN(n762) );
  NAND2_X1 U808 ( .A1(n762), .A2(n761), .ZN(n769) );
  NOR2_X1 U809 ( .A1(n669), .A2(G953), .ZN(n767) );
  NAND2_X1 U810 ( .A1(G953), .A2(G224), .ZN(n763) );
  XNOR2_X1 U811 ( .A(KEYINPUT61), .B(n763), .ZN(n764) );
  NAND2_X1 U812 ( .A1(n764), .A2(G898), .ZN(n765) );
  XOR2_X1 U813 ( .A(KEYINPUT124), .B(n765), .Z(n766) );
  NOR2_X1 U814 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U815 ( .A(n769), .B(n768), .ZN(G69) );
  XOR2_X1 U816 ( .A(n771), .B(n770), .Z(n775) );
  XNOR2_X1 U817 ( .A(n772), .B(n775), .ZN(n774) );
  NAND2_X1 U818 ( .A1(n774), .A2(n773), .ZN(n780) );
  XNOR2_X1 U819 ( .A(G227), .B(n775), .ZN(n776) );
  NAND2_X1 U820 ( .A1(n776), .A2(G900), .ZN(n777) );
  XNOR2_X1 U821 ( .A(KEYINPUT126), .B(n777), .ZN(n778) );
  NAND2_X1 U822 ( .A1(n778), .A2(G953), .ZN(n779) );
  NAND2_X1 U823 ( .A1(n780), .A2(n779), .ZN(G72) );
  XOR2_X1 U824 ( .A(n781), .B(G122), .Z(G24) );
  XNOR2_X1 U825 ( .A(G137), .B(n782), .ZN(G39) );
  XNOR2_X1 U826 ( .A(n783), .B(G131), .ZN(G33) );
endmodule

