//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT0), .B(G128), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  OR2_X1    g012(.A1(KEYINPUT65), .A2(G137), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT11), .A2(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT65), .A2(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT11), .A2(G134), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT11), .A2(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n206), .B1(new_n202), .B2(new_n205), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n198), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n199), .A2(new_n211), .A3(new_n201), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n206), .B1(G134), .B2(G137), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n190), .B(new_n192), .C1(KEYINPUT1), .C2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n191), .A2(G146), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n189), .A2(G143), .ZN(new_n219));
  OAI211_X1 g033(.A(G128), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n207), .A2(new_n214), .A3(new_n216), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n210), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G116), .ZN(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G113), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT2), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G113), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n231), .ZN(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n236), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n210), .A2(new_n238), .A3(new_n221), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n188), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n188), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(G237), .A2(G953), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G210), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT27), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G101), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n248), .A2(KEYINPUT29), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n243), .A2(KEYINPUT69), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT69), .B1(new_n243), .B2(new_n249), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n187), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n253));
  AND4_X1   g067(.A1(new_n207), .A2(new_n214), .A3(new_n216), .A4(new_n220), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n194), .B(new_n255), .C1(new_n195), .C2(new_n196), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  OR2_X1    g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n258), .B(new_n259), .C1(new_n218), .C2(new_n219), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n255), .B1(new_n260), .B2(new_n194), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n202), .A2(new_n205), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G131), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n207), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n254), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n253), .B1(new_n266), .B2(KEYINPUT30), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n210), .A2(KEYINPUT30), .A3(new_n221), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n197), .A2(KEYINPUT64), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n269), .B(new_n256), .C1(new_n208), .C2(new_n209), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n221), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(KEYINPUT66), .A3(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n267), .A2(new_n236), .A3(new_n268), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n239), .ZN(new_n275));
  INV_X1    g089(.A(new_n248), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT68), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n278));
  AOI211_X1 g092(.A(new_n278), .B(new_n248), .C1(new_n274), .C2(new_n239), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n238), .B1(new_n270), .B2(new_n221), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n210), .A2(new_n238), .A3(new_n221), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT28), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n281), .B1(new_n284), .B2(new_n241), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n239), .B1(new_n266), .B2(new_n238), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT67), .B1(new_n286), .B2(KEYINPUT28), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n285), .A2(new_n287), .A3(new_n276), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(KEYINPUT29), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n252), .B1(new_n280), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G472), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n276), .B1(new_n285), .B2(new_n287), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n283), .A2(new_n276), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n274), .A2(KEYINPUT31), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT31), .B1(new_n274), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n300));
  OAI22_X1  g114(.A1(new_n290), .A2(new_n291), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G214), .B1(G237), .B2(G902), .ZN(new_n302));
  OAI21_X1  g116(.A(G210), .B1(G237), .B2(G902), .ZN(new_n303));
  XNOR2_X1  g117(.A(G110), .B(G122), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G104), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT3), .B1(new_n306), .B2(G107), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n308));
  INV_X1    g122(.A(G107), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(G104), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(G107), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n307), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(G101), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n236), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(KEYINPUT74), .A3(G101), .ZN(new_n316));
  AOI21_X1  g130(.A(G101), .B1(new_n306), .B2(G107), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n307), .A2(new_n317), .A3(new_n310), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n316), .A2(KEYINPUT4), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n312), .A2(G101), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n315), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n225), .A2(G119), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT5), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n228), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT5), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n235), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n306), .A2(G107), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n309), .A2(G104), .ZN(new_n331));
  OAI21_X1  g145(.A(G101), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n318), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT78), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n332), .A2(new_n318), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n326), .A2(new_n327), .B1(new_n234), .B2(new_n233), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n305), .B1(new_n323), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n318), .A2(KEYINPUT4), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n322), .A2(new_n316), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n236), .A3(new_n314), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n343), .A2(new_n304), .A3(new_n334), .A4(new_n338), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n340), .A2(new_n344), .A3(new_n345), .A4(KEYINPUT6), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n340), .A2(new_n344), .A3(KEYINPUT6), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT6), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n348), .B(new_n305), .C1(new_n323), .C2(new_n339), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT79), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n346), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  AOI211_X1 g165(.A(KEYINPUT80), .B(G125), .C1(new_n220), .C2(new_n216), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n220), .A2(new_n216), .ZN(new_n353));
  INV_X1    g167(.A(G125), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n197), .B2(G125), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n352), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G224), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G953), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n358), .B(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n351), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n357), .A2(new_n355), .ZN(new_n365));
  OAI211_X1 g179(.A(KEYINPUT7), .B(new_n361), .C1(new_n365), .C2(new_n352), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(KEYINPUT7), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n358), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT81), .B1(new_n335), .B2(new_n336), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n329), .A2(new_n333), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n329), .A2(KEYINPUT81), .A3(new_n333), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n304), .B(KEYINPUT8), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n366), .A2(new_n368), .A3(new_n374), .A4(KEYINPUT82), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n375), .A2(new_n344), .ZN(new_n376));
  INV_X1    g190(.A(new_n373), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n369), .B2(new_n370), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n372), .A2(new_n378), .B1(new_n358), .B2(new_n367), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n366), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(G902), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n303), .B1(new_n364), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n340), .A2(new_n344), .A3(KEYINPUT6), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT79), .A3(new_n349), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n362), .B1(new_n386), .B2(new_n346), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n375), .A2(new_n344), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT82), .B1(new_n379), .B2(new_n366), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n187), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n303), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n387), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n302), .B1(new_n384), .B2(new_n392), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n314), .A2(new_n194), .A3(new_n260), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n342), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n265), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n220), .A2(new_n332), .A3(new_n318), .A4(new_n216), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT75), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT10), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT10), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n395), .A2(new_n396), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT76), .A2(KEYINPUT12), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n353), .A2(new_n333), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n397), .ZN(new_n406));
  NOR2_X1   g220(.A1(KEYINPUT76), .A2(KEYINPUT12), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(new_n264), .B2(new_n207), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n408), .A3(new_n404), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n403), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G110), .B(G140), .ZN(new_n413));
  INV_X1    g227(.A(G953), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n414), .A2(G227), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n400), .A2(new_n402), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n198), .A2(new_n314), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n319), .B2(new_n322), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n265), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n416), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n403), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(G902), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G469), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT77), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n421), .A2(new_n403), .A3(new_n422), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n406), .A2(new_n408), .A3(new_n404), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(new_n409), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n422), .B1(new_n429), .B2(new_n403), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n187), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT77), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(G469), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n412), .A2(new_n416), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n422), .B1(new_n421), .B2(new_n403), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n425), .B(new_n187), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n426), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT9), .B(G234), .ZN(new_n438));
  OAI21_X1  g252(.A(G221), .B1(new_n438), .B2(G902), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n393), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT22), .B(G137), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n414), .A2(G221), .A3(G234), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n354), .A2(KEYINPUT16), .A3(G140), .ZN(new_n446));
  XNOR2_X1  g260(.A(G125), .B(G140), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n446), .B1(new_n447), .B2(KEYINPUT16), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G146), .ZN(new_n449));
  INV_X1    g263(.A(G140), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G125), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n354), .A2(G140), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT73), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT73), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n189), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n449), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g272(.A(KEYINPUT71), .B(G110), .Z(new_n459));
  NAND3_X1  g273(.A1(new_n215), .A2(KEYINPUT23), .A3(G119), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n223), .A2(G128), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT23), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n223), .B2(G128), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n459), .A2(new_n460), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT72), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n215), .A2(G119), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT24), .B(G110), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n464), .A2(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n463), .A2(new_n461), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n470), .A2(KEYINPUT72), .A3(new_n460), .A4(new_n459), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n458), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n467), .A2(new_n468), .ZN(new_n473));
  INV_X1    g287(.A(new_n446), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT16), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n474), .A2(new_n475), .A3(G146), .ZN(new_n476));
  AOI21_X1  g290(.A(G146), .B1(new_n474), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n463), .A2(new_n460), .A3(new_n461), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n463), .A2(new_n460), .A3(KEYINPUT70), .A4(new_n461), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n481), .A2(G110), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n445), .B1(new_n472), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n464), .A2(new_n465), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n467), .A2(new_n468), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n471), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n458), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n481), .A2(G110), .A3(new_n482), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n491), .B(new_n473), .C1(new_n477), .C2(new_n476), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n444), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n485), .A2(new_n493), .A3(new_n187), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n485), .A2(new_n493), .A3(KEYINPUT25), .A4(new_n187), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G217), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(G234), .B2(new_n187), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n485), .A2(new_n493), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n500), .A2(G902), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n244), .A2(G143), .A3(G214), .ZN(new_n507));
  AOI21_X1  g321(.A(G143), .B1(new_n244), .B2(G214), .ZN(new_n508));
  OAI21_X1  g322(.A(G131), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n510));
  INV_X1    g324(.A(G237), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n414), .A3(G214), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n191), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n244), .A2(G143), .A3(G214), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n206), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n509), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n477), .ZN(new_n517));
  OAI211_X1 g331(.A(KEYINPUT17), .B(G131), .C1(new_n507), .C2(new_n508), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n449), .A4(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(KEYINPUT83), .A2(KEYINPUT18), .ZN(new_n520));
  OAI211_X1 g334(.A(G131), .B(new_n520), .C1(new_n507), .C2(new_n508), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(G131), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n514), .A3(new_n522), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n455), .A2(new_n189), .A3(new_n456), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n447), .A2(new_n189), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n521), .B(new_n523), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G113), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(new_n306), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n519), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT19), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n455), .A2(new_n530), .A3(new_n456), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT84), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n453), .A2(new_n532), .A3(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT84), .B1(new_n447), .B2(new_n530), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n531), .A2(new_n189), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n509), .A2(new_n515), .B1(new_n448), .B2(G146), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n528), .B1(new_n537), .B2(new_n526), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n529), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G475), .A2(G902), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT86), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n540), .B1(new_n541), .B2(KEYINPUT20), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n541), .B2(new_n540), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT85), .B1(new_n529), .B2(new_n538), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n519), .A2(new_n526), .A3(new_n528), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT85), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n521), .A2(new_n523), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n457), .B1(new_n189), .B2(new_n447), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n548), .A2(new_n549), .B1(new_n535), .B2(new_n536), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n546), .B(new_n547), .C1(new_n550), .C2(new_n528), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n545), .A2(new_n540), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n544), .B1(new_n552), .B2(KEYINPUT20), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n519), .A2(new_n526), .ZN(new_n554));
  INV_X1    g368(.A(new_n528), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n556), .B2(new_n546), .ZN(new_n557));
  INV_X1    g371(.A(G475), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G478), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n438), .A2(new_n499), .A3(G953), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G122), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G116), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(KEYINPUT87), .A2(G122), .ZN(new_n569));
  NAND2_X1  g383(.A1(KEYINPUT87), .A2(G122), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n309), .B(new_n568), .C1(new_n571), .C2(new_n225), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n225), .B1(new_n569), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT14), .B1(new_n566), .B2(G116), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT14), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n225), .A3(G122), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G107), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(G128), .B(G143), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n579), .A2(G134), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(G134), .ZN(new_n581));
  AND4_X1   g395(.A1(new_n572), .A2(new_n578), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(G107), .B1(new_n573), .B2(new_n567), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n215), .A2(G143), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n211), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n586), .A2(new_n579), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n579), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n572), .A2(new_n583), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n565), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n572), .A2(new_n578), .A3(new_n580), .A4(new_n581), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n572), .A2(new_n583), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n587), .A2(new_n588), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n591), .B(new_n564), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n563), .B1(new_n595), .B2(new_n187), .ZN(new_n596));
  AOI211_X1 g410(.A(G902), .B(new_n562), .C1(new_n590), .C2(new_n594), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n560), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n414), .A2(G952), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(G234), .B2(G237), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT21), .B(G898), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT88), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n187), .B(new_n414), .C1(G234), .C2(G237), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n301), .A2(new_n441), .A3(new_n506), .A4(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  NAND3_X1  g423(.A1(new_n364), .A2(new_n383), .A3(new_n303), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n391), .B1(new_n387), .B2(new_n390), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n606), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n302), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n595), .A2(new_n561), .A3(new_n187), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n561), .A2(new_n187), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n595), .A2(KEYINPUT33), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n590), .B2(new_n594), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n618), .B1(new_n622), .B2(G478), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n614), .A2(new_n560), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n296), .A2(new_n298), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n274), .A2(new_n293), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT31), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n274), .A2(KEYINPUT31), .A3(new_n293), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(G902), .B1(new_n631), .B2(new_n292), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n626), .B1(new_n632), .B2(new_n291), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n633), .A2(new_n440), .A3(new_n505), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n625), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT89), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT34), .B(G104), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  INV_X1    g452(.A(KEYINPUT20), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n552), .B(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n598), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n556), .A2(new_n546), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n187), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT90), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n645), .A3(G475), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT90), .B1(new_n557), .B2(new_n558), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n641), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n614), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n634), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  AOI21_X1  g467(.A(new_n291), .B1(new_n296), .B2(new_n187), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n298), .B2(new_n296), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n445), .A2(KEYINPUT36), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n492), .B2(new_n490), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n472), .A2(new_n484), .A3(new_n656), .ZN(new_n659));
  INV_X1    g473(.A(new_n503), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n498), .B2(new_n500), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n441), .A2(new_n607), .A3(new_n655), .A4(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n601), .B1(new_n605), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n641), .A2(new_n642), .A3(new_n648), .A4(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n662), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n301), .A2(new_n441), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  INV_X1    g487(.A(new_n440), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n668), .B(KEYINPUT39), .Z(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT40), .Z(new_n677));
  INV_X1    g491(.A(KEYINPUT92), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n612), .B(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n276), .B1(new_n274), .B2(new_n239), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n237), .A2(new_n239), .A3(new_n276), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n187), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n299), .B2(new_n300), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n560), .A2(new_n598), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n302), .A3(new_n662), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n680), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n677), .A2(new_n678), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n689), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n676), .B(KEYINPUT40), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT92), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n191), .ZN(G45));
  OAI211_X1 g509(.A(new_n623), .B(new_n669), .C1(new_n553), .C2(new_n559), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n662), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n301), .A2(new_n441), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NOR4_X1   g513(.A1(new_n277), .A2(new_n279), .A3(new_n288), .A4(KEYINPUT29), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n700), .B2(new_n252), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n626), .A2(KEYINPUT32), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n505), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n187), .B1(new_n434), .B2(new_n435), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n439), .A3(new_n436), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT93), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT93), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n710), .A3(new_n439), .A4(new_n436), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n625), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT94), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n715), .B(new_n717), .ZN(G15));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n650), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  NOR2_X1   g534(.A1(new_n393), .A2(new_n708), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n599), .A2(new_n606), .A3(new_n662), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n301), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  AND3_X1   g538(.A1(new_n709), .A2(new_n613), .A3(new_n711), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n612), .A2(new_n302), .A3(new_n687), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n298), .B(KEYINPUT95), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n276), .B1(new_n240), .B2(new_n242), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n728), .B1(new_n631), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n654), .A2(new_n730), .A3(new_n505), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n725), .A2(new_n726), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT96), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n566), .ZN(G24));
  NOR3_X1   g549(.A1(new_n654), .A2(new_n730), .A3(new_n662), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT97), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n696), .B(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n721), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  INV_X1    g554(.A(new_n302), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n612), .A2(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n301), .A2(new_n506), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n439), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n417), .A2(KEYINPUT98), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT98), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n430), .A2(new_n746), .ZN(new_n747));
  AND4_X1   g561(.A1(G469), .A2(new_n745), .A3(new_n747), .A4(new_n423), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n425), .A2(new_n187), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n436), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT99), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n427), .B1(new_n746), .B2(new_n430), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(G469), .A3(new_n745), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT99), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n436), .A4(new_n750), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n744), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n743), .A2(KEYINPUT42), .A3(new_n738), .A4(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n301), .A2(new_n506), .A3(new_n757), .A4(new_n742), .ZN(new_n760));
  INV_X1    g574(.A(new_n738), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n758), .A2(KEYINPUT100), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT100), .B1(new_n758), .B2(new_n762), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  INV_X1    g580(.A(new_n670), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n705), .A2(new_n767), .A3(new_n757), .A4(new_n742), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  AND3_X1   g583(.A1(new_n753), .A2(KEYINPUT45), .A3(new_n745), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT45), .B1(new_n417), .B2(new_n423), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n770), .A2(new_n425), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n749), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(KEYINPUT46), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n436), .B1(new_n773), .B2(KEYINPUT46), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n439), .B(new_n675), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n553), .A2(new_n559), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT101), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n553), .A2(KEYINPUT101), .A3(new_n559), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(KEYINPUT43), .A3(new_n779), .A4(new_n623), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n777), .B2(new_n624), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT102), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(KEYINPUT102), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n655), .A2(new_n662), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n776), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n784), .A2(KEYINPUT44), .A3(new_n785), .A4(new_n786), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT103), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n790), .A2(new_n791), .A3(new_n742), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n791), .B1(new_n790), .B2(new_n742), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  INV_X1    g609(.A(new_n301), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n506), .A2(new_n696), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n742), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n439), .B1(new_n774), .B2(new_n775), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT47), .B(new_n439), .C1(new_n774), .C2(new_n775), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(new_n450), .ZN(G42));
  NOR2_X1   g618(.A1(new_n440), .A2(new_n505), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n560), .A2(new_n623), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n598), .B2(new_n560), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n741), .B(new_n606), .C1(new_n610), .C2(new_n611), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n805), .A2(new_n655), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n723), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n705), .B(new_n712), .C1(new_n625), .C2(new_n650), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n608), .A4(new_n664), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n646), .A2(new_n598), .A3(new_n647), .A4(new_n669), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n640), .A2(new_n813), .A3(new_n662), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n440), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n301), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n738), .A2(new_n757), .A3(new_n736), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n742), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n768), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n812), .A2(new_n820), .A3(new_n734), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n758), .B2(new_n762), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n301), .B(new_n441), .C1(new_n671), .C2(new_n697), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n662), .A2(new_n669), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT105), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n726), .A2(new_n685), .A3(new_n757), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n825), .A2(KEYINPUT52), .A3(new_n739), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT106), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n825), .A2(new_n739), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT106), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT52), .A4(new_n829), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n825), .A2(new_n739), .A3(new_n829), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT107), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n836), .B1(new_n835), .B2(new_n837), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n831), .B(new_n834), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT108), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n835), .A2(new_n837), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT107), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n830), .B(new_n833), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT108), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n824), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n843), .A2(new_n830), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n765), .A2(new_n821), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n822), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n849), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n765), .A2(new_n821), .A3(new_n822), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n840), .A2(new_n841), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT108), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n760), .A2(new_n670), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n819), .B1(new_n816), .B2(new_n817), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n732), .B(KEYINPUT96), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n608), .A2(new_n664), .A3(new_n723), .A4(new_n809), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .A4(new_n811), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n865), .A2(new_n763), .A3(new_n764), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n822), .B1(new_n866), .B2(new_n851), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n854), .B1(new_n869), .B2(new_n850), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  INV_X1    g685(.A(new_n736), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n819), .A2(new_n708), .ZN(new_n873));
  INV_X1    g687(.A(new_n601), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n780), .B2(new_n782), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT112), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n873), .A2(KEYINPUT112), .A3(new_n875), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n872), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n506), .A2(new_n873), .A3(new_n601), .A4(new_n686), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(new_n560), .A3(new_n624), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n875), .A2(new_n731), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n708), .A2(new_n302), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n680), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(KEYINPUT110), .B2(KEYINPUT50), .ZN(new_n889));
  NOR2_X1   g703(.A1(KEYINPUT110), .A2(KEYINPUT50), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n885), .B2(new_n887), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n884), .A2(KEYINPUT113), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT113), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n881), .A2(new_n893), .A3(new_n883), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n871), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n883), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT113), .B1(new_n896), .B2(new_n880), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n889), .A2(new_n891), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n894), .A3(new_n871), .A4(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n707), .A2(new_n744), .A3(new_n436), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n801), .A2(new_n802), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n885), .A2(new_n819), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT115), .B1(new_n895), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n600), .B(KEYINPUT116), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n885), .A2(new_n393), .A3(new_n708), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n560), .A2(new_n624), .ZN(new_n909));
  AOI211_X1 g723(.A(new_n907), .B(new_n908), .C1(new_n909), .C2(new_n882), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n878), .A2(new_n879), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT48), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n912), .A3(new_n705), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n912), .B1(new_n911), .B2(new_n705), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n884), .B1(KEYINPUT111), .B2(new_n898), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n801), .A2(KEYINPUT109), .A3(new_n802), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n901), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT109), .B1(new_n801), .B2(new_n802), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n903), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n898), .A2(KEYINPUT111), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n917), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n916), .B1(new_n923), .B2(new_n900), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n897), .A2(new_n894), .A3(new_n898), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT114), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT115), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n926), .A2(new_n927), .A3(new_n899), .A4(new_n904), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n906), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  OAI22_X1  g743(.A1(new_n870), .A2(new_n929), .B1(G952), .B2(G953), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n623), .A2(new_n302), .A3(new_n439), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n707), .A2(new_n436), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n505), .B(new_n931), .C1(KEYINPUT49), .C2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n778), .A3(new_n779), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT104), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n680), .B(new_n686), .C1(KEYINPUT49), .C2(new_n932), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(G75));
  AOI21_X1  g751(.A(new_n187), .B1(new_n849), .B2(new_n853), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(G210), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n351), .B(new_n363), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT55), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n941), .A2(KEYINPUT56), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n414), .A2(G952), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT117), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT56), .B1(new_n939), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n938), .A2(KEYINPUT117), .A3(G210), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n946), .B1(new_n950), .B2(new_n941), .ZN(G51));
  XNOR2_X1  g765(.A(new_n749), .B(KEYINPUT57), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n821), .A2(new_n823), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n856), .B2(new_n857), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT53), .B1(new_n866), .B2(new_n851), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT54), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n850), .B1(new_n849), .B2(new_n853), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n435), .B2(new_n434), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n938), .A2(new_n772), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n944), .B1(new_n959), .B2(new_n960), .ZN(G54));
  NAND2_X1  g775(.A1(new_n545), .A2(new_n551), .ZN(new_n962));
  INV_X1    g776(.A(new_n938), .ZN(new_n963));
  NAND2_X1  g777(.A1(KEYINPUT58), .A2(G475), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n945), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n963), .A2(new_n962), .A3(new_n964), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(G60));
  INV_X1    g782(.A(new_n622), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n616), .B(KEYINPUT59), .Z(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n956), .B2(new_n957), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(KEYINPUT118), .A3(new_n945), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT118), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT54), .B1(new_n954), .B2(new_n955), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n971), .B1(new_n854), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n975), .B1(new_n977), .B2(new_n944), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n858), .A2(new_n850), .A3(new_n867), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n970), .B1(new_n979), .B2(new_n956), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n622), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n974), .A2(new_n978), .A3(new_n981), .ZN(G63));
  NAND2_X1  g796(.A1(G217), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT119), .Z(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT60), .Z(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n954), .B2(new_n955), .ZN(new_n986));
  INV_X1    g800(.A(new_n502), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n944), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n985), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n849), .B2(new_n853), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n658), .A2(new_n659), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT120), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n991), .B(new_n985), .C1(new_n954), .C2(new_n955), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT120), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n988), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT61), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g812(.A(KEYINPUT61), .B(new_n988), .C1(new_n992), .C2(new_n995), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(G66));
  AOI21_X1  g814(.A(new_n414), .B1(new_n603), .B2(G224), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n812), .A2(new_n734), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1001), .B1(new_n1003), .B2(new_n414), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n386), .B(new_n346), .C1(G898), .C2(new_n414), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1004), .B(new_n1005), .Z(G69));
  NAND3_X1  g820(.A1(new_n267), .A2(new_n268), .A3(new_n273), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G900), .A2(G953), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n705), .A2(new_n726), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n832), .B(new_n768), .C1(new_n776), .C2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n803), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n794), .A2(new_n1013), .A3(new_n765), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1009), .B(new_n1010), .C1(new_n1014), .C2(G953), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT124), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  INV_X1    g832(.A(new_n803), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n743), .A2(new_n674), .A3(new_n675), .A4(new_n807), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n794), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT62), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n690), .A2(new_n693), .A3(new_n1022), .A4(new_n832), .ZN(new_n1023));
  OR2_X1    g837(.A1(new_n1023), .A2(KEYINPUT121), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(KEYINPUT121), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n690), .A2(new_n693), .A3(new_n832), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT122), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(G953), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n1017), .B(new_n1018), .C1(new_n1031), .C2(new_n1009), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n414), .B1(G227), .B2(G900), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1033), .B(KEYINPUT123), .Z(new_n1035));
  OAI211_X1 g849(.A(new_n1015), .B(new_n1035), .C1(new_n1031), .C2(new_n1009), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1034), .A2(new_n1036), .ZN(G72));
  NAND2_X1  g851(.A1(G472), .A2(G902), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT63), .Z(new_n1039));
  XNOR2_X1  g853(.A(new_n1039), .B(KEYINPUT125), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1040), .B1(new_n1014), .B2(new_n1003), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n275), .A2(new_n248), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n944), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n280), .A2(new_n627), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(new_n1039), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1043), .B1(new_n869), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1021), .ZN(new_n1048));
  NAND4_X1  g862(.A1(new_n1030), .A2(new_n1002), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1049), .A2(new_n1040), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1050), .A2(new_n681), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1051), .A2(KEYINPUT126), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT126), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1050), .A2(new_n1053), .A3(new_n681), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1046), .B1(new_n1052), .B2(new_n1054), .ZN(G57));
endmodule


