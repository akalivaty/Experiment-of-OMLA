//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n434, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n568, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(new_n434));
  INV_X1    g009(.A(new_n434), .ZN(G218));
  INV_X1    g010(.A(G132), .ZN(G219));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(KEYINPUT70), .B(KEYINPUT3), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n472), .B1(new_n466), .B2(G2104), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n464), .B(new_n465), .C1(new_n471), .C2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  INV_X1    g050(.A(G101), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n469), .A2(new_n465), .A3(new_n470), .ZN(new_n477));
  OAI22_X1  g052(.A1(new_n474), .A2(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  XNOR2_X1  g056(.A(KEYINPUT3), .B(G2104), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G125), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  NAND2_X1  g063(.A1(new_n469), .A2(new_n470), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n473), .B1(new_n489), .B2(KEYINPUT3), .ZN(new_n490));
  INV_X1    g065(.A(new_n464), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(G124), .A3(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n474), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  OR2_X1    g070(.A1(G100), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR4_X1   g075(.A1(new_n483), .A2(KEYINPUT4), .A3(new_n500), .A4(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT74), .B1(new_n474), .B2(new_n500), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT3), .B1(new_n462), .B2(new_n463), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT70), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n507), .A2(G138), .A3(new_n465), .A4(new_n464), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(KEYINPUT74), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n502), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT73), .B(G114), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G2105), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n507), .A2(G126), .A3(G2105), .A4(new_n464), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(KEYINPUT72), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n492), .A2(new_n516), .A3(G126), .A4(G2105), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n510), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G164));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT5), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT75), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT6), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT6), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(KEYINPUT75), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n526), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  INV_X1    g108(.A(G50), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n529), .A2(G543), .A3(new_n531), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n526), .A2(G62), .ZN(new_n537));
  NAND2_X1  g112(.A1(G75), .A2(G543), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT76), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n528), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n536), .A2(new_n540), .ZN(G166));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT77), .Z(new_n543));
  INV_X1    g118(.A(new_n535), .ZN(new_n544));
  AOI22_X1  g119(.A1(KEYINPUT7), .A2(new_n543), .B1(new_n544), .B2(G51), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n545), .B1(KEYINPUT7), .B2(new_n543), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n547));
  INV_X1    g122(.A(G89), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n532), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G168));
  NAND2_X1  g125(.A1(new_n529), .A2(new_n531), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n523), .A2(new_n525), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(G90), .A2(new_n553), .B1(new_n544), .B2(G52), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT78), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n528), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  NAND2_X1  g134(.A1(new_n553), .A2(G81), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n544), .A2(G43), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n560), .B(new_n561), .C1(new_n528), .C2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT79), .ZN(G188));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OR3_X1    g147(.A1(new_n535), .A2(KEYINPUT9), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT9), .B1(new_n535), .B2(new_n572), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n552), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n573), .A2(new_n574), .B1(G651), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n553), .B(KEYINPUT80), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n579), .A2(KEYINPUT81), .A3(G91), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT81), .B1(new_n579), .B2(G91), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G168), .ZN(G286));
  INV_X1    g158(.A(G166), .ZN(G303));
  AND2_X1   g159(.A1(new_n579), .A2(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(new_n535), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n526), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G48), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n591), .A2(new_n528), .B1(new_n592), .B2(new_n535), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n579), .B2(G86), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT82), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n553), .A2(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n544), .A2(G47), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n597), .B(new_n598), .C1(new_n528), .C2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n579), .A2(G92), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT10), .Z(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT83), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n552), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(new_n544), .B2(G54), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G297));
  XNOR2_X1  g189(.A(G297), .B(KEYINPUT84), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n609), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n564), .ZN(new_n620));
  MUX2_X1   g195(.A(new_n619), .B(new_n620), .S(KEYINPUT85), .Z(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g197(.A1(new_n483), .A2(new_n477), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n494), .A2(G135), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n465), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n492), .A2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(G123), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n627), .B1(new_n628), .B2(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n626), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G1341), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT87), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G1348), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(new_n654), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n659), .A2(KEYINPUT17), .A3(new_n656), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n656), .B1(new_n659), .B2(KEYINPUT17), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n660), .A2(new_n661), .A3(new_n655), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n673), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  OAI221_X1 g252(.A(new_n674), .B1(new_n673), .B2(new_n671), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n677), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1991), .ZN(new_n680));
  INV_X1    g255(.A(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1986), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT88), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1981), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n595), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G6), .B2(new_n690), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(G16), .A2(G23), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n589), .B2(G16), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT33), .B(G1976), .Z(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n690), .A2(G22), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G166), .B2(new_n690), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n702), .A2(G1971), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(G1971), .ZN(new_n704));
  NOR4_X1   g279(.A1(new_n699), .A2(new_n700), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n694), .A2(new_n695), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT34), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n494), .A2(G131), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n465), .A2(G107), .ZN(new_n709));
  OAI21_X1  g284(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n710));
  INV_X1    g285(.A(G119), .ZN(new_n711));
  OAI221_X1 g286(.A(new_n708), .B1(new_n709), .B2(new_n710), .C1(new_n630), .C2(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G25), .B(new_n712), .S(G29), .Z(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT35), .B(G1991), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n690), .A2(G24), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G290), .B2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G1986), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT89), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n718), .B2(new_n719), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n707), .A2(new_n716), .A3(new_n720), .A4(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G32), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT94), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT26), .ZN(new_n731));
  INV_X1    g306(.A(G105), .ZN(new_n732));
  OAI22_X1  g307(.A1(new_n730), .A2(new_n731), .B1(new_n732), .B2(new_n477), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n731), .B2(new_n730), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n494), .A2(G141), .ZN(new_n735));
  INV_X1    g310(.A(G129), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n734), .B(new_n735), .C1(new_n736), .C2(new_n630), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT95), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(KEYINPUT95), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n728), .B1(new_n741), .B2(new_n727), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT96), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n742), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n727), .A2(G26), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT28), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n494), .A2(G140), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n465), .A2(G116), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G128), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n748), .B1(new_n749), .B2(new_n750), .C1(new_n630), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G29), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(KEYINPUT91), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(KEYINPUT91), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n747), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2067), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n727), .A2(G27), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G164), .B2(new_n727), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G2078), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n745), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n727), .A2(G33), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  INV_X1    g339(.A(G139), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n474), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT92), .Z(new_n767));
  AOI22_X1  g342(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n465), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT93), .Z(new_n770));
  OAI21_X1  g345(.A(new_n762), .B1(new_n770), .B2(new_n727), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2072), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n690), .A2(G4), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n609), .B2(new_n690), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT90), .B(G1348), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n774), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n690), .A2(G21), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G168), .B2(new_n690), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT97), .B(G1966), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n690), .A2(G19), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n564), .B2(new_n690), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1341), .ZN(new_n784));
  INV_X1    g359(.A(G28), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(KEYINPUT30), .ZN(new_n786));
  AOI21_X1  g361(.A(G29), .B1(new_n785), .B2(KEYINPUT30), .ZN(new_n787));
  OR2_X1    g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  NAND2_X1  g363(.A1(KEYINPUT31), .A2(G11), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n632), .B2(new_n727), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n781), .A2(new_n784), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G5), .A2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G171), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1961), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n777), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT24), .ZN(new_n798));
  INV_X1    g373(.A(G34), .ZN(new_n799));
  AOI21_X1  g374(.A(G29), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n798), .B2(new_n799), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G160), .B2(new_n727), .ZN(new_n802));
  INV_X1    g377(.A(G2084), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n727), .A2(G35), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT98), .Z(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G162), .B2(new_n727), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT29), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n804), .B1(G2090), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n690), .A2(G20), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT99), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT23), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n613), .B2(new_n690), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G1956), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n808), .A2(G2090), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n772), .A2(new_n797), .A3(new_n809), .A4(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n725), .A2(new_n726), .A3(new_n761), .A4(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  NAND2_X1  g394(.A1(new_n609), .A2(G559), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n553), .A2(G93), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n544), .A2(G55), .ZN(new_n822));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  INV_X1    g398(.A(G67), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n552), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G651), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n821), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n564), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n829), .B(new_n830), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n820), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n834));
  AOI21_X1  g409(.A(G860), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n827), .A2(G860), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT101), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(G145));
  XNOR2_X1  g415(.A(new_n740), .B(new_n752), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n520), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  INV_X1    g418(.A(new_n770), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n844), .B2(KEYINPUT102), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n842), .B(new_n845), .C1(new_n843), .C2(new_n844), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n842), .B2(new_n845), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n712), .B(new_n624), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n487), .B(new_n632), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n494), .A2(G142), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n465), .A2(G118), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  INV_X1    g428(.A(G130), .ZN(new_n854));
  OAI221_X1 g429(.A(new_n851), .B1(new_n852), .B2(new_n853), .C1(new_n630), .C2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G162), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n850), .B(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(G37), .B1(new_n849), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n849), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT40), .ZN(G395));
  OR3_X1    g435(.A1(new_n609), .A2(KEYINPUT104), .A3(G299), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT104), .B1(new_n609), .B2(G299), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n609), .A2(G299), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n618), .B(new_n831), .Z(new_n867));
  MUX2_X1   g442(.A(new_n864), .B(new_n866), .S(new_n867), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n595), .B(G166), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n589), .B(G290), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n872));
  OR3_X1    g447(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT42), .ZN(new_n873));
  INV_X1    g448(.A(new_n871), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n868), .B(new_n876), .ZN(new_n877));
  MUX2_X1   g452(.A(new_n827), .B(new_n877), .S(G868), .Z(G295));
  MUX2_X1   g453(.A(new_n827), .B(new_n877), .S(G868), .Z(G331));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n880));
  AOI21_X1  g455(.A(G168), .B1(G301), .B2(KEYINPUT107), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(KEYINPUT107), .B2(G301), .ZN(new_n882));
  OR3_X1    g457(.A1(G301), .A2(G286), .A3(KEYINPUT107), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(new_n831), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n831), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n885), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n888), .B1(new_n885), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n890), .A2(new_n864), .B1(new_n866), .B2(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(new_n874), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n889), .A2(new_n866), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n889), .A2(new_n866), .A3(KEYINPUT109), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n864), .B1(new_n892), .B2(new_n893), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n899), .A2(new_n874), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n896), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n880), .B1(new_n904), .B2(KEYINPUT43), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n903), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n900), .A2(new_n901), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n874), .B1(new_n907), .B2(new_n899), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n910));
  OAI21_X1  g485(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n906), .B2(new_n908), .ZN(new_n913));
  INV_X1    g488(.A(new_n910), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n896), .A2(new_n902), .A3(new_n903), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n912), .B1(new_n916), .B2(new_n880), .ZN(new_n917));
  AOI211_X1 g492(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n913), .C2(new_n915), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n911), .B1(new_n917), .B2(new_n918), .ZN(G397));
  INV_X1    g494(.A(G1384), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT4), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n508), .B2(KEYINPUT74), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT74), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n492), .A2(new_n923), .A3(G138), .A4(new_n465), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n501), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n920), .B1(new_n925), .B2(new_n518), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n480), .A2(G40), .A3(new_n486), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n712), .A2(new_n714), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n741), .A2(new_n681), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n740), .A2(G1996), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n752), .B(G2067), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n930), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(G2067), .B2(new_n752), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT124), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n930), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n939), .B2(new_n938), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n930), .A2(new_n681), .ZN(new_n942));
  NAND2_X1  g517(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n942), .B(new_n943), .Z(new_n944));
  OAI21_X1  g519(.A(new_n930), .B1(new_n740), .B2(new_n934), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n944), .B(new_n945), .C1(KEYINPUT125), .C2(KEYINPUT46), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT47), .Z(new_n947));
  OR3_X1    g522(.A1(new_n936), .A2(G1986), .A3(G290), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n712), .B(new_n715), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n935), .A2(new_n952), .ZN(new_n953));
  AOI211_X1 g528(.A(new_n950), .B(new_n951), .C1(new_n930), .C2(new_n953), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n941), .A2(new_n947), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT123), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n478), .A2(KEYINPUT71), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n478), .A2(KEYINPUT71), .ZN(new_n958));
  AND4_X1   g533(.A1(G40), .A2(new_n957), .A3(new_n486), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT112), .B1(new_n520), .B2(new_n920), .ZN(new_n960));
  OAI211_X1 g535(.A(KEYINPUT112), .B(new_n920), .C1(new_n925), .C2(new_n518), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1976), .ZN(new_n964));
  NOR2_X1   g539(.A1(G288), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(G8), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n926), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n929), .B1(new_n969), .B2(new_n961), .ZN(new_n970));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1981), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n594), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT114), .B(G86), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n553), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(G1981), .B1(new_n593), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n974), .A2(KEYINPUT49), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT49), .B1(new_n974), .B2(new_n977), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n967), .A2(KEYINPUT52), .B1(new_n972), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT52), .B1(G288), .B2(new_n964), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n963), .A2(new_n966), .A3(G8), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(G303), .A2(G8), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n984), .B(KEYINPUT55), .Z(new_n985));
  NAND3_X1  g560(.A1(new_n969), .A2(KEYINPUT50), .A3(new_n961), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n510), .B2(new_n519), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n929), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G2090), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n986), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1971), .ZN(new_n992));
  INV_X1    g567(.A(new_n928), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT45), .B(new_n920), .C1(new_n925), .C2(new_n518), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n959), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n992), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n971), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n981), .B(new_n983), .C1(new_n985), .C2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT50), .B1(new_n969), .B2(new_n961), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n959), .B1(new_n987), .B2(new_n988), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n999), .A2(new_n1000), .A3(G2090), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n959), .A2(new_n994), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1971), .B1(new_n1002), .B2(new_n928), .ZN(new_n1003));
  OAI211_X1 g578(.A(G8), .B(new_n985), .C1(new_n1001), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n988), .B1(new_n960), .B2(new_n962), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1000), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n990), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n971), .B1(new_n1009), .B2(new_n996), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(KEYINPUT113), .A3(new_n985), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n998), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G168), .A2(new_n971), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n969), .A2(new_n927), .A3(new_n961), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n1002), .ZN(new_n1019));
  INV_X1    g594(.A(G1966), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1007), .A2(new_n1008), .A3(new_n803), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(G8), .B(new_n1017), .C1(new_n1023), .C2(G286), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n999), .A2(new_n1000), .A3(G2084), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1966), .B1(new_n1018), .B2(new_n1002), .ZN(new_n1026));
  OAI21_X1  g601(.A(G8), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1014), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n1016), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1023), .A2(new_n1014), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1024), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n795), .B1(new_n999), .B2(new_n1000), .ZN(new_n1032));
  INV_X1    g607(.A(G2078), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n928), .A2(new_n1033), .A3(new_n959), .A4(new_n994), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(G2078), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1018), .A2(new_n1002), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1032), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G171), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1012), .A2(KEYINPUT62), .A3(new_n1031), .A4(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n963), .A2(new_n980), .A3(G8), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n970), .A2(new_n971), .A3(new_n965), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n983), .B(new_n1043), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1006), .A2(new_n1011), .A3(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1043), .A2(new_n964), .A3(new_n589), .ZN(new_n1049));
  INV_X1    g624(.A(new_n974), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n972), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1042), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n985), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n999), .A2(new_n1000), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1003), .B1(new_n1055), .B2(new_n990), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1054), .B1(new_n1056), .B2(new_n971), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1047), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1009), .A2(new_n996), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n985), .B1(new_n1060), .B2(G8), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT115), .B1(new_n1061), .B2(new_n1046), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1006), .A2(new_n1011), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1023), .A2(G8), .A3(G168), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT63), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n997), .A2(new_n985), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(new_n1046), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1065), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1064), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1063), .A2(new_n1068), .B1(new_n1072), .B2(new_n1066), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1053), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT113), .B1(new_n1010), .B2(new_n985), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1070), .B(new_n1041), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1024), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(KEYINPUT62), .B2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1032), .A2(new_n1038), .A3(G301), .A4(new_n1036), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n485), .A2(KEYINPUT120), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n465), .B1(new_n485), .B2(KEYINPUT120), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n480), .A2(G40), .A3(new_n1083), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1084), .A2(KEYINPUT121), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1037), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(new_n1084), .B2(KEYINPUT121), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1085), .A2(new_n1087), .A3(new_n994), .A4(new_n928), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n1036), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1032), .A2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT119), .B(new_n795), .C1(new_n999), .C2(new_n1000), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT54), .B(new_n1080), .C1(new_n1093), .C2(G301), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(new_n1064), .A3(new_n1070), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n776), .B1(new_n999), .B2(new_n1000), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n1097));
  INV_X1    g672(.A(G2067), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n970), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1096), .A2(new_n1097), .A3(new_n609), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n928), .A2(new_n681), .A3(new_n959), .A4(new_n994), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT58), .B(G1341), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1102), .B1(new_n970), .B2(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1104), .A2(KEYINPUT59), .A3(new_n564), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT59), .B1(new_n1104), .B2(new_n564), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1101), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n1108));
  XNOR2_X1  g683(.A(G299), .B(KEYINPUT57), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n986), .A2(new_n989), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT116), .B(G1956), .Z(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT56), .B(G2072), .Z(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AND4_X1   g690(.A1(new_n959), .A2(new_n928), .A3(new_n994), .A4(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1110), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1112), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n986), .B2(new_n989), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1120), .A2(new_n1109), .A3(new_n1116), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1108), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1113), .A2(new_n1110), .A3(new_n1117), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1109), .B1(new_n1120), .B2(new_n1116), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(KEYINPUT61), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n609), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1096), .A2(new_n1126), .A3(new_n1099), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT60), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1107), .A2(new_n1122), .A3(new_n1125), .A4(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1118), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1095), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1089), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(G301), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1040), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1135), .B1(new_n1093), .B2(G301), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1133), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1079), .B1(new_n1132), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1074), .B1(new_n1141), .B2(new_n1031), .ZN(new_n1142));
  XNOR2_X1  g717(.A(G290), .B(G1986), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n930), .B1(new_n953), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n956), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1094), .A2(new_n1064), .A3(new_n1070), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1122), .A2(new_n1147), .A3(new_n1100), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1129), .A2(new_n1125), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1131), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1150), .A3(new_n1140), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1078), .A2(KEYINPUT62), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1152), .A2(new_n1012), .A3(new_n1041), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1031), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1072), .A2(new_n1066), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1059), .A2(new_n1062), .A3(new_n1064), .A4(new_n1067), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(new_n1042), .A3(new_n1052), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n956), .B(new_n1144), .C1(new_n1154), .C2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n955), .B1(new_n1145), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT126), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1163), .B(new_n955), .C1(new_n1145), .C2(new_n1160), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g740(.A(G319), .ZN(new_n1167));
  NOR3_X1   g741(.A1(G401), .A2(new_n1167), .A3(G227), .ZN(new_n1168));
  NAND3_X1  g742(.A1(new_n687), .A2(new_n688), .A3(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g743(.A(new_n1169), .B(KEYINPUT127), .ZN(new_n1170));
  NAND3_X1  g744(.A1(new_n916), .A2(new_n859), .A3(new_n1170), .ZN(G225));
  INV_X1    g745(.A(G225), .ZN(G308));
endmodule


