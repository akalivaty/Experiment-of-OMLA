//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT76), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT76), .A2(G104), .ZN(new_n191));
  AOI21_X1  g005(.A(G107), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(G107), .A3(new_n191), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n196), .A3(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G101), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT76), .A2(G104), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT76), .A2(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n196), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT3), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT77), .B(G101), .Z(new_n204));
  NAND4_X1  g018(.A1(new_n203), .A2(new_n204), .A3(new_n195), .A4(new_n197), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(KEYINPUT4), .A3(new_n205), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT2), .B(G113), .Z(new_n207));
  XNOR2_X1  g021(.A(G116), .B(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G116), .ZN(new_n211));
  INV_X1    g025(.A(G116), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT2), .B(G113), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n209), .A2(KEYINPUT66), .A3(new_n216), .ZN(new_n217));
  OR3_X1    g031(.A1(new_n207), .A2(KEYINPUT66), .A3(new_n208), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n220), .B(G101), .C1(new_n194), .C2(new_n198), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n206), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n204), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n194), .A2(new_n198), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G101), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n196), .A2(G104), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n226), .B1(new_n202), .B2(KEYINPUT78), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT78), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(new_n196), .C1(new_n200), .C2(new_n201), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(G113), .B1(new_n211), .B2(KEYINPUT5), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n208), .A2(KEYINPUT5), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n233), .A2(new_n234), .B1(new_n208), .B2(new_n207), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n238));
  XNOR2_X1  g052(.A(G110), .B(G122), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n222), .A2(new_n236), .A3(new_n239), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT6), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n239), .B1(new_n222), .B2(new_n236), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n187), .B(new_n241), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n244), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n246), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n242), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G143), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(KEYINPUT1), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G128), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n250), .B(new_n252), .C1(KEYINPUT1), .C2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n250), .A2(new_n252), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT65), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G143), .B(G146), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT65), .A3(new_n259), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n262), .A2(new_n264), .B1(new_n253), .B2(new_n266), .ZN(new_n267));
  MUX2_X1   g081(.A(new_n258), .B(new_n267), .S(G125), .Z(new_n268));
  INV_X1    g082(.A(G224), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(G953), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n268), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n248), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G210), .B1(G237), .B2(G902), .ZN(new_n274));
  INV_X1    g088(.A(new_n231), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n235), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n239), .B(KEYINPUT8), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n232), .A2(KEYINPUT83), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n232), .A2(KEYINPUT83), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n234), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n280), .A2(new_n209), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n276), .B(new_n277), .C1(new_n275), .C2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT7), .B1(new_n269), .B2(G953), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n268), .B(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n284), .A3(new_n242), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n273), .A2(new_n274), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT84), .ZN(new_n290));
  INV_X1    g104(.A(new_n274), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n271), .B1(new_n245), .B2(new_n247), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(new_n287), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n273), .A2(KEYINPUT84), .A3(new_n274), .A4(new_n288), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT74), .ZN(new_n298));
  OAI21_X1  g112(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n299));
  XOR2_X1   g113(.A(new_n299), .B(KEYINPUT75), .Z(new_n300));
  NAND2_X1  g114(.A1(new_n255), .A2(new_n257), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n224), .B2(new_n230), .ZN(new_n302));
  INV_X1    g116(.A(new_n226), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(new_n192), .B2(new_n228), .ZN(new_n304));
  INV_X1    g118(.A(new_n229), .ZN(new_n305));
  OAI21_X1  g119(.A(G101), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(new_n258), .A3(new_n205), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT11), .ZN(new_n309));
  INV_X1    g123(.A(G134), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(G137), .ZN(new_n311));
  INV_X1    g125(.A(G137), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT11), .A3(G134), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(G137), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G131), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n311), .A2(new_n313), .A3(new_n317), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT12), .B1(new_n308), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT12), .ZN(new_n321));
  INV_X1    g135(.A(new_n319), .ZN(new_n322));
  AOI211_X1 g136(.A(new_n321), .B(new_n322), .C1(new_n302), .C2(new_n307), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT79), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n224), .A2(new_n230), .A3(new_n301), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n258), .B1(new_n306), .B2(new_n205), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n321), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n308), .A2(KEYINPUT12), .A3(new_n319), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT10), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n307), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n206), .A2(new_n267), .A3(new_n221), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n306), .A2(KEYINPUT10), .A3(new_n258), .A4(new_n205), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n322), .A4(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G140), .ZN(new_n337));
  INV_X1    g151(.A(G227), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(G953), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n337), .B(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n324), .A2(new_n331), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n319), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n336), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n340), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G469), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT70), .B(G902), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n336), .B1(new_n320), .B2(new_n323), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n340), .A2(new_n352), .B1(new_n342), .B2(new_n345), .ZN(new_n353));
  OAI21_X1  g167(.A(G469), .B1(new_n353), .B2(G902), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n300), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G125), .B(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT71), .ZN(new_n357));
  INV_X1    g171(.A(G140), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n358), .A2(KEYINPUT71), .A3(G125), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(KEYINPUT16), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT16), .B1(new_n358), .B2(G125), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G146), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n249), .A3(new_n363), .ZN(new_n366));
  NOR2_X1   g180(.A1(G237), .A2(G953), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G214), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n251), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(G143), .A3(G214), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(KEYINPUT17), .A3(G131), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(G131), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT17), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n369), .A2(new_n317), .A3(new_n370), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n365), .A2(new_n366), .A3(new_n372), .A4(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G113), .B(G122), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(new_n189), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT18), .A2(G131), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n371), .B(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT73), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n356), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n356), .A2(new_n382), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n249), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n359), .B1(new_n356), .B2(KEYINPUT71), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G146), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n377), .A2(new_n379), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n379), .B1(new_n377), .B2(new_n389), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n286), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G475), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n377), .A2(new_n379), .A3(new_n389), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n364), .A2(G146), .B1(new_n373), .B2(new_n375), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n386), .A2(KEYINPUT19), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n383), .A2(new_n384), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n249), .B(new_n396), .C1(new_n397), .C2(KEYINPUT19), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n395), .A2(new_n398), .B1(new_n381), .B2(new_n388), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n394), .B1(new_n379), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT20), .ZN(new_n401));
  NOR2_X1   g215(.A1(G475), .A2(G902), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n400), .B2(new_n402), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n393), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G478), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(KEYINPUT15), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(KEYINPUT15), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n350), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT13), .B1(new_n256), .B2(G143), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(new_n310), .ZN(new_n414));
  XNOR2_X1  g228(.A(G128), .B(G143), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G122), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G116), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n212), .A2(G122), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT85), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT85), .ZN(new_n422));
  AOI21_X1  g236(.A(G107), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n422), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n424), .A2(new_n420), .A3(new_n196), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n416), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n196), .B1(new_n424), .B2(new_n420), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n415), .B(new_n310), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n417), .A2(G116), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n196), .B1(new_n429), .B2(KEYINPUT14), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT14), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n418), .A2(new_n419), .A3(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n431), .B1(new_n430), .B2(new_n433), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n427), .B(new_n428), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n426), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G217), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n298), .A2(new_n438), .A3(G953), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n426), .A2(new_n439), .A3(new_n436), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n412), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT89), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n411), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(KEYINPUT87), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n426), .A2(new_n439), .A3(new_n436), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n439), .B1(new_n426), .B2(new_n436), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n350), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n411), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n443), .B2(KEYINPUT89), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n445), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G953), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G952), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(G234), .B2(G237), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n456), .B(new_n350), .C1(G234), .C2(G237), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(G898), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n405), .A2(new_n455), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n355), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G214), .B1(G237), .B2(G902), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT80), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT81), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n296), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n438), .B1(new_n350), .B2(G234), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT22), .B(G137), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n456), .A2(G221), .A3(G234), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT23), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n210), .B2(G128), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n256), .A2(KEYINPUT23), .A3(G119), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n473), .B(new_n474), .C1(G119), .C2(new_n256), .ZN(new_n475));
  XNOR2_X1  g289(.A(G119), .B(G128), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT24), .B(G110), .Z(new_n477));
  AOI22_X1  g291(.A1(new_n475), .A2(G110), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI211_X1 g292(.A(G146), .B(new_n362), .C1(new_n386), .C2(KEYINPUT16), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n249), .B1(new_n361), .B2(new_n363), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT72), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT72), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n483), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI22_X1  g299(.A1(new_n475), .A2(G110), .B1(new_n476), .B2(new_n477), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n385), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n480), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n471), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n471), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n488), .B(new_n491), .C1(new_n482), .C2(new_n484), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT25), .B1(new_n493), .B2(new_n350), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n495));
  NOR4_X1   g309(.A1(new_n490), .A2(new_n492), .A3(new_n495), .A4(new_n412), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n468), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n468), .A2(G902), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n267), .A2(new_n319), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n217), .A2(new_n218), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n310), .A2(G137), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n312), .A2(G134), .ZN(new_n504));
  OAI21_X1  g318(.A(G131), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n255), .A2(new_n318), .A3(new_n505), .A4(new_n257), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n501), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n502), .B1(new_n501), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT28), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XOR2_X1   g323(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n510));
  NAND2_X1  g324(.A1(new_n367), .A2(G210), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT26), .B(G101), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n318), .A2(new_n505), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n267), .A2(new_n319), .B1(new_n258), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n502), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT28), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n509), .A2(KEYINPUT29), .A3(new_n514), .A4(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT69), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT28), .B1(new_n516), .B2(new_n502), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n253), .A2(new_n266), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT65), .B1(new_n263), .B2(new_n259), .ZN(new_n524));
  AND4_X1   g338(.A1(KEYINPUT65), .A2(new_n250), .A3(new_n252), .A4(new_n259), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n506), .B1(new_n322), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n219), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n517), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n522), .B1(new_n529), .B2(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n514), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT29), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n516), .B2(KEYINPUT64), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT64), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n527), .A2(new_n535), .A3(KEYINPUT30), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n502), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(new_n507), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n531), .B(new_n532), .C1(new_n538), .C2(new_n514), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n521), .A2(new_n539), .A3(new_n350), .ZN(new_n540));
  NOR2_X1   g354(.A1(G472), .A2(G902), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n516), .A2(KEYINPUT64), .A3(new_n533), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT30), .B1(new_n527), .B2(new_n535), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n219), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n517), .A3(new_n514), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n514), .B1(new_n509), .B2(new_n519), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n546), .B1(KEYINPUT31), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT31), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n545), .A2(new_n549), .A3(new_n517), .A4(new_n514), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n542), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n540), .A2(G472), .B1(new_n551), .B2(KEYINPUT32), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n509), .A2(new_n519), .ZN(new_n553));
  INV_X1    g367(.A(new_n514), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT31), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n537), .A2(new_n507), .A3(new_n554), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n550), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n541), .ZN(new_n558));
  XOR2_X1   g372(.A(KEYINPUT68), .B(KEYINPUT32), .Z(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n500), .B1(new_n552), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n467), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(new_n223), .ZN(G3));
  INV_X1    g377(.A(new_n355), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n557), .A2(new_n350), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n551), .B1(G472), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n564), .A2(new_n567), .A3(new_n500), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT91), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT90), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n447), .B2(new_n448), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT33), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n570), .B(KEYINPUT33), .C1(new_n447), .C2(new_n448), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n350), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G478), .ZN(new_n577));
  AOI21_X1  g391(.A(G478), .B1(new_n446), .B2(new_n451), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n569), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n406), .B1(new_n575), .B2(new_n350), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n581), .A2(KEYINPUT91), .A3(new_n578), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n405), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AOI211_X1 g398(.A(new_n465), .B(new_n461), .C1(new_n289), .C2(new_n293), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n568), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT92), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT34), .B(G104), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G6));
  NAND2_X1  g403(.A1(new_n289), .A2(new_n293), .ZN(new_n590));
  INV_X1    g404(.A(new_n465), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT93), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n403), .B2(new_n404), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n395), .A2(new_n398), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n379), .B1(new_n594), .B2(new_n389), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n390), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n402), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT20), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(KEYINPUT93), .A3(new_n599), .ZN(new_n600));
  AND4_X1   g414(.A1(new_n393), .A2(new_n593), .A3(new_n455), .A4(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n461), .ZN(new_n602));
  AND4_X1   g416(.A1(new_n590), .A2(new_n591), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n568), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G107), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  NAND2_X1  g420(.A1(new_n485), .A2(new_n489), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n491), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n485), .A2(new_n489), .A3(new_n471), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n350), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n495), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n493), .A2(KEYINPUT25), .A3(new_n350), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n491), .A2(KEYINPUT36), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n607), .B(new_n614), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n613), .A2(new_n468), .B1(new_n498), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n567), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n467), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT37), .B(G110), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT94), .B(KEYINPUT95), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G12));
  AOI21_X1  g436(.A(new_n616), .B1(new_n552), .B2(new_n560), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n465), .B1(new_n289), .B2(new_n293), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n355), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n593), .A2(new_n455), .A3(new_n600), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT96), .B(G900), .Z(new_n627));
  NAND2_X1  g441(.A1(new_n459), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n458), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n393), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n625), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n256), .ZN(G30));
  XNOR2_X1  g449(.A(new_n630), .B(KEYINPUT39), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n355), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT97), .Z(new_n638));
  OR2_X1    g452(.A1(new_n638), .A2(KEYINPUT40), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(KEYINPUT40), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n296), .B(KEYINPUT38), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n551), .A2(KEYINPUT32), .ZN(new_n642));
  INV_X1    g456(.A(new_n538), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n514), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n286), .B1(new_n529), .B2(new_n514), .ZN(new_n646));
  OAI21_X1  g460(.A(G472), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n560), .A2(new_n642), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n405), .A2(new_n455), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n616), .A2(new_n591), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n641), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n639), .A2(new_n640), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n251), .ZN(G45));
  OAI211_X1 g467(.A(new_n405), .B(new_n630), .C1(new_n580), .C2(new_n582), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n623), .A2(new_n655), .A3(new_n355), .A4(new_n624), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(KEYINPUT98), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(KEYINPUT98), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G146), .ZN(G48));
  NAND2_X1  g474(.A1(new_n348), .A2(new_n350), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G469), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n351), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n300), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n561), .A2(new_n664), .A3(new_n584), .A4(new_n585), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT41), .B(G113), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT99), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n665), .B(new_n667), .ZN(G15));
  NAND3_X1  g482(.A1(new_n603), .A2(new_n561), .A3(new_n664), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G116), .ZN(G18));
  INV_X1    g484(.A(new_n300), .ZN(new_n671));
  AND4_X1   g485(.A1(new_n462), .A2(new_n662), .A3(new_n671), .A4(new_n351), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n623), .A2(KEYINPUT100), .A3(new_n672), .A4(new_n624), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n531), .A2(new_n532), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n514), .B1(new_n545), .B2(new_n517), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n350), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT69), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n520), .B(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n560), .A3(new_n642), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n615), .A2(new_n498), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n497), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n681), .A2(new_n624), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n462), .A2(new_n662), .A3(new_n671), .A4(new_n351), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n674), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n673), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n210), .ZN(G21));
  AND2_X1   g502(.A1(new_n624), .A2(new_n649), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n565), .A2(G472), .ZN(new_n690));
  AOI211_X1 g504(.A(KEYINPUT101), .B(new_n542), .C1(new_n548), .C2(new_n550), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n557), .B2(new_n541), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n690), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n500), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n689), .A2(new_n695), .A3(new_n664), .A4(new_n602), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G122), .ZN(G24));
  NOR3_X1   g511(.A1(new_n654), .A2(new_n694), .A3(new_n616), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n664), .A2(new_n624), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(G125), .Z(G27));
  AOI21_X1  g516(.A(new_n465), .B1(new_n294), .B2(new_n295), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n703), .A2(new_n655), .ZN(new_n704));
  OR3_X1    g518(.A1(new_n551), .A2(KEYINPUT104), .A3(KEYINPUT32), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT104), .B1(new_n551), .B2(KEYINPUT32), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n552), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n708));
  INV_X1    g522(.A(new_n500), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n708), .B1(new_n707), .B2(new_n709), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n704), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI211_X1 g526(.A(G469), .B(new_n412), .C1(new_n343), .C2(new_n347), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n345), .A2(new_n336), .A3(new_n341), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n330), .A2(new_n328), .B1(new_n715), .B2(new_n322), .ZN(new_n716));
  OAI211_X1 g530(.A(G469), .B(new_n714), .C1(new_n716), .C2(new_n341), .ZN(new_n717));
  NAND2_X1  g531(.A1(G469), .A2(G902), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT102), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n351), .A2(new_n354), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n671), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT103), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n720), .A2(new_n725), .A3(new_n722), .A4(new_n671), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT42), .B1(new_n712), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n724), .A2(new_n561), .A3(new_n726), .A4(new_n703), .ZN(new_n729));
  OR3_X1    g543(.A1(new_n729), .A2(KEYINPUT42), .A3(new_n654), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  AND3_X1   g546(.A1(new_n724), .A2(new_n726), .A3(new_n703), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(KEYINPUT106), .A3(new_n561), .A4(new_n632), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n735), .B1(new_n729), .B2(new_n633), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  OAI21_X1  g552(.A(G469), .B1(new_n353), .B2(KEYINPUT45), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n352), .A2(new_n340), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(KEYINPUT45), .A3(new_n714), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n718), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n744), .B(KEYINPUT107), .Z(new_n745));
  OR2_X1    g559(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n713), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n745), .B(new_n748), .C1(new_n747), .C2(new_n746), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(new_n671), .ZN(new_n750));
  INV_X1    g564(.A(new_n582), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT91), .B1(new_n581), .B2(new_n578), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n405), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n755), .B(KEYINPUT43), .Z(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n567), .A3(new_n683), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n703), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n750), .A2(new_n759), .A3(new_n636), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  XOR2_X1   g577(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n764));
  OR2_X1    g578(.A1(new_n750), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n750), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n709), .A2(new_n681), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n765), .A2(new_n704), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n771));
  OAI22_X1  g585(.A1(new_n699), .A2(new_n700), .B1(new_n625), .B2(new_n633), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n657), .B2(new_n658), .ZN(new_n773));
  INV_X1    g587(.A(new_n689), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n616), .A2(new_n630), .ZN(new_n775));
  OR4_X1    g589(.A1(new_n648), .A2(new_n774), .A3(new_n723), .A4(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(KEYINPUT52), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(new_n773), .B2(new_n776), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n771), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n779), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(KEYINPUT114), .A3(new_n777), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n696), .A2(new_n669), .A3(new_n665), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n687), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n296), .A2(new_n466), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n754), .A2(new_n455), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n461), .B1(new_n583), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n568), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n562), .A2(new_n618), .A3(new_n789), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n728), .A2(new_n785), .A3(new_n730), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n698), .A2(new_n724), .A3(new_n726), .A4(new_n703), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n455), .A2(new_n631), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n355), .A2(new_n600), .A3(new_n593), .A4(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(new_n623), .A3(new_n703), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n792), .B1(new_n737), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g613(.A(KEYINPUT112), .B(new_n797), .C1(new_n734), .C2(new_n736), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n791), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n791), .B(KEYINPUT113), .C1(new_n799), .C2(new_n800), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n783), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(KEYINPUT115), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n781), .A2(new_n777), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n803), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT115), .B1(new_n805), .B2(new_n806), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT54), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n809), .A2(new_n806), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT116), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n809), .A2(new_n815), .A3(new_n806), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n731), .A2(KEYINPUT53), .A3(new_n785), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n799), .A2(new_n800), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n790), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n821), .B1(new_n820), .B2(new_n790), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n783), .B(new_n819), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n817), .A2(new_n818), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n812), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n694), .A2(new_n500), .A3(new_n629), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n756), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n700), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n703), .A2(new_n458), .A3(new_n664), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n648), .A2(new_n709), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n457), .B(new_n830), .C1(new_n584), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n756), .A2(new_n831), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n710), .A2(new_n711), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n834), .B1(KEYINPUT48), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(KEYINPUT48), .B2(new_n837), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n641), .A2(new_n465), .A3(new_n664), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(KEYINPUT119), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(KEYINPUT119), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n756), .A3(new_n843), .A4(new_n828), .ZN(new_n844));
  XOR2_X1   g658(.A(KEYINPUT120), .B(KEYINPUT50), .Z(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n835), .A2(new_n616), .A3(new_n694), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n753), .A2(new_n405), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n847), .B1(new_n833), .B2(new_n848), .ZN(new_n849));
  OR2_X1    g663(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n846), .B(new_n849), .C1(new_n850), .C2(new_n844), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n765), .A2(new_n767), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n663), .B(KEYINPUT110), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n671), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n829), .A2(new_n760), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n851), .A2(KEYINPUT121), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(KEYINPUT51), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n851), .A2(KEYINPUT121), .ZN(new_n860));
  OAI221_X1 g674(.A(new_n839), .B1(KEYINPUT51), .B2(new_n856), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n827), .A2(new_n861), .B1(G952), .B2(G953), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n853), .B(KEYINPUT49), .Z(new_n863));
  NOR3_X1   g677(.A1(new_n755), .A2(new_n466), .A3(new_n300), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n641), .A3(new_n832), .A4(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT111), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n862), .A2(new_n866), .ZN(G75));
  NOR2_X1   g681(.A1(new_n456), .A2(G952), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n809), .A2(new_n815), .A3(new_n806), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n815), .B1(new_n809), .B2(new_n806), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n825), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(new_n412), .A3(new_n291), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n248), .A2(new_n272), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n292), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT55), .Z(new_n878));
  OAI21_X1  g692(.A(new_n869), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n350), .B1(new_n817), .B2(new_n825), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n880), .B2(new_n291), .ZN(new_n881));
  INV_X1    g695(.A(new_n878), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT122), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n884), .A3(new_n878), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n879), .B1(new_n883), .B2(new_n885), .ZN(G51));
  INV_X1    g700(.A(new_n818), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n872), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n888), .A2(new_n826), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n718), .B(KEYINPUT57), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n348), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n739), .A2(new_n741), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n880), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n868), .B1(new_n891), .B2(new_n893), .ZN(G54));
  NAND4_X1  g708(.A1(new_n872), .A2(KEYINPUT58), .A3(G475), .A4(new_n412), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n895), .A2(KEYINPUT123), .A3(new_n596), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n869), .B1(new_n895), .B2(new_n596), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT123), .B1(new_n895), .B2(new_n596), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(G60));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT59), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n575), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n869), .B1(new_n889), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n575), .B1(new_n827), .B2(new_n902), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(G63));
  NAND2_X1  g720(.A1(G217), .A2(G902), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT60), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n872), .A2(new_n615), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n817), .B2(new_n825), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n910), .B(new_n869), .C1(new_n911), .C2(new_n493), .ZN(new_n912));
  OAI211_X1 g726(.A(KEYINPUT124), .B(new_n869), .C1(new_n911), .C2(new_n493), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n872), .A2(new_n909), .ZN(new_n916));
  INV_X1    g730(.A(new_n493), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n868), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n918), .B(new_n910), .C1(KEYINPUT124), .C2(KEYINPUT61), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n919), .ZN(G66));
  INV_X1    g734(.A(new_n460), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n456), .B1(new_n921), .B2(G224), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n785), .A2(new_n790), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n923), .B2(new_n456), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n245), .B(new_n247), .C1(G898), .C2(new_n456), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n924), .B(new_n925), .Z(G69));
  NOR2_X1   g740(.A1(new_n543), .A2(new_n544), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n396), .B1(new_n397), .B2(KEYINPUT19), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n927), .B(new_n928), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(G900), .B(G953), .C1(new_n930), .C2(G227), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(G227), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n836), .A2(new_n774), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n750), .A2(new_n636), .A3(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n762), .A2(new_n773), .A3(new_n934), .ZN(new_n935));
  AND4_X1   g749(.A1(new_n731), .A2(new_n935), .A3(new_n769), .A4(new_n737), .ZN(new_n936));
  AOI21_X1  g750(.A(G953), .B1(new_n936), .B2(new_n930), .ZN(new_n937));
  INV_X1    g751(.A(new_n652), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n773), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT125), .ZN(new_n941));
  INV_X1    g755(.A(new_n561), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n583), .A2(new_n787), .ZN(new_n943));
  OR4_X1    g757(.A1(new_n942), .A2(new_n638), .A3(new_n760), .A4(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n762), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n769), .B(new_n945), .C1(KEYINPUT62), .C2(new_n939), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n929), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n932), .B1(new_n937), .B2(new_n947), .ZN(G72));
  NOR2_X1   g762(.A1(new_n676), .A2(new_n556), .ZN(new_n949));
  NAND2_X1  g763(.A1(G472), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT63), .Z(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n868), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n941), .A2(new_n946), .A3(new_n644), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n643), .A2(new_n514), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n936), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n953), .B1(new_n956), .B2(new_n923), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n949), .A2(new_n952), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT126), .Z(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n810), .B2(new_n811), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(G57));
endmodule


