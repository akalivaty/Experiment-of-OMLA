//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT67), .B(G120gat), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT68), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(G120gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n208), .B(G113gat), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n206), .A2(new_n207), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n214));
  XNOR2_X1  g013(.A(G127gat), .B(G134gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n217));
  INV_X1    g016(.A(G134gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G127gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(G113gat), .B(G120gat), .ZN(new_n220));
  OAI221_X1 g019(.A(new_n217), .B1(KEYINPUT66), .B2(new_n219), .C1(KEYINPUT1), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G155gat), .ZN(new_n223));
  INV_X1    g022(.A(G162gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(G141gat), .B(G148gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n225), .B(new_n226), .C1(new_n227), .C2(KEYINPUT2), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT73), .ZN(new_n229));
  INV_X1    g028(.A(G148gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G141gat), .ZN(new_n231));
  INV_X1    g030(.A(G141gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G148gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT2), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT73), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n236), .A2(new_n237), .A3(new_n225), .A4(new_n226), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT74), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n227), .A2(KEYINPUT74), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n226), .B1(new_n225), .B2(KEYINPUT2), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n229), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n222), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n229), .A2(new_n238), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n246), .A2(new_n243), .B1(new_n216), .B2(new_n221), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n203), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT75), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT5), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n222), .A2(new_n244), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n229), .A2(new_n238), .A3(new_n243), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(new_n221), .A3(new_n216), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n202), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT5), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT75), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n221), .A4(new_n216), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n229), .A2(new_n238), .A3(new_n243), .A4(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n222), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n258), .A2(new_n259), .A3(new_n202), .A4(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n250), .A2(new_n256), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n258), .A2(new_n259), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT76), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n263), .A2(new_n255), .A3(new_n202), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n258), .A2(KEYINPUT76), .A3(new_n259), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G1gat), .B(G29gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(G85gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT0), .B(G57gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n265), .A2(new_n271), .A3(new_n276), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n272), .A2(KEYINPUT6), .A3(new_n277), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  AND2_X1   g083(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n287), .A2(KEYINPUT28), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT26), .ZN(new_n292));
  INV_X1    g091(.A(G169gat), .ZN(new_n293));
  INV_X1    g092(.A(G176gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT26), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n292), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n287), .A2(KEYINPUT28), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n288), .A2(new_n289), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n289), .A2(KEYINPUT24), .ZN(new_n303));
  NOR2_X1   g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI22_X1  g104(.A1(new_n290), .A2(KEYINPUT23), .B1(new_n289), .B2(KEYINPUT24), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n305), .A2(new_n306), .A3(new_n295), .ZN(new_n307));
  AND2_X1   g106(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n309));
  OAI211_X1 g108(.A(KEYINPUT23), .B(new_n294), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n302), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n291), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G183gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n284), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(KEYINPUT24), .A3(new_n289), .ZN(new_n316));
  OR2_X1    g115(.A1(new_n289), .A2(KEYINPUT24), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n313), .A2(new_n316), .A3(new_n296), .A4(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT25), .B1(new_n291), .B2(new_n312), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n301), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n222), .ZN(new_n322));
  NAND2_X1  g121(.A1(G227gat), .A2(G233gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n302), .ZN(new_n324));
  INV_X1    g123(.A(new_n310), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n324), .B1(new_n318), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n319), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n307), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n329), .A2(new_n221), .A3(new_n216), .A4(new_n301), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n322), .A2(new_n323), .A3(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n331), .B(KEYINPUT34), .Z(new_n332));
  XNOR2_X1  g131(.A(G15gat), .B(G43gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(G71gat), .ZN(new_n334));
  INV_X1    g133(.A(G99gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n323), .B1(new_n322), .B2(new_n330), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(KEYINPUT33), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT32), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n322), .A2(new_n330), .ZN(new_n342));
  INV_X1    g141(.A(new_n323), .ZN(new_n343));
  AOI221_X4 g142(.A(new_n339), .B1(KEYINPUT33), .B2(new_n336), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n332), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n321), .A2(new_n222), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n329), .A2(new_n301), .B1(new_n216), .B2(new_n221), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT32), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT33), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n351), .A3(new_n336), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n331), .B(KEYINPUT34), .ZN(new_n353));
  INV_X1    g152(.A(new_n336), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n348), .B(KEYINPUT32), .C1(new_n350), .C2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n345), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G197gat), .B(G204gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT22), .ZN(new_n359));
  INV_X1    g158(.A(G211gat), .ZN(new_n360));
  INV_X1    g159(.A(G218gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G211gat), .B(G218gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n358), .A3(new_n362), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n261), .B1(new_n368), .B2(KEYINPUT78), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n367), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n370), .A2(KEYINPUT78), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n244), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n370), .B(KEYINPUT70), .Z(new_n376));
  NAND2_X1  g175(.A1(new_n262), .A2(new_n371), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(KEYINPUT79), .B(new_n244), .C1(new_n369), .C2(new_n372), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G228gat), .ZN(new_n381));
  INV_X1    g180(.A(G233gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n377), .A2(new_n367), .A3(new_n366), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n244), .B1(KEYINPUT3), .B2(new_n368), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n385), .B(new_n386), .C1(new_n381), .C2(new_n382), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389));
  INV_X1    g188(.A(G22gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(KEYINPUT31), .B(G50gat), .Z(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n384), .A2(new_n387), .A3(new_n393), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n357), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n399), .B(KEYINPUT71), .Z(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n321), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n329), .B2(new_n301), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(new_n401), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n376), .ZN(new_n405));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n402), .B(new_n370), .C1(new_n403), .C2(new_n401), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT72), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n405), .A2(KEYINPUT72), .A3(new_n409), .A4(new_n410), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n411), .A2(new_n415), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n405), .A2(new_n410), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n408), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n283), .A2(new_n398), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT35), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n281), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n278), .A2(KEYINPUT77), .A3(new_n279), .A4(new_n280), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n282), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n421), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT69), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n341), .B2(new_n344), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n353), .B1(new_n352), .B2(new_n355), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n353), .A2(new_n432), .B1(new_n433), .B2(new_n431), .ZN(new_n434));
  INV_X1    g233(.A(new_n397), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n430), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT69), .B1(new_n352), .B2(new_n355), .ZN(new_n437));
  OAI22_X1  g236(.A1(new_n345), .A2(KEYINPUT69), .B1(new_n437), .B2(new_n332), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n397), .A3(KEYINPUT82), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(KEYINPUT35), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n424), .B1(new_n429), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n357), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n442), .A2(KEYINPUT36), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n434), .A2(KEYINPUT36), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n445), .B1(new_n429), .B2(new_n435), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n405), .A2(new_n447), .A3(new_n410), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n404), .A2(new_n370), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n402), .B(new_n376), .C1(new_n403), .C2(new_n401), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(KEYINPUT37), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT38), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n448), .A2(new_n451), .A3(new_n452), .A4(new_n408), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n453), .A2(new_n413), .A3(new_n414), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n281), .A2(new_n454), .A3(new_n282), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT81), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n408), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n447), .B1(new_n405), .B2(new_n410), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT38), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n281), .A2(new_n454), .A3(new_n460), .A4(new_n282), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n456), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n268), .A2(new_n263), .A3(new_n270), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT39), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n203), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n276), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n251), .A2(new_n253), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT39), .B1(new_n468), .B2(new_n203), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT80), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT80), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(KEYINPUT39), .C1(new_n468), .C2(new_n203), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n203), .B2(new_n464), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n463), .B1(new_n467), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n464), .A2(new_n203), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(new_n470), .A3(new_n472), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n477), .A2(KEYINPUT40), .A3(new_n276), .A4(new_n466), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n475), .A2(new_n478), .A3(new_n420), .A4(new_n278), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n397), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n441), .B1(new_n446), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G15gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n390), .ZN(new_n483));
  NAND2_X1  g282(.A1(G15gat), .A2(G22gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G1gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT16), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n483), .A2(new_n486), .A3(new_n484), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT89), .B(G8gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(KEYINPUT87), .A3(new_n489), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n489), .A2(KEYINPUT87), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(G8gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT88), .A4(G8gat), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n492), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT21), .ZN(new_n500));
  NAND2_X1  g299(.A1(KEYINPUT91), .A2(G57gat), .ZN(new_n501));
  INV_X1    g300(.A(G64gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G71gat), .A2(G78gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(G71gat), .A2(G78gat), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n505), .B1(KEYINPUT9), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT92), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n501), .B(G64gat), .ZN(new_n509));
  INV_X1    g308(.A(new_n506), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT9), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n504), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n511), .B1(G57gat), .B2(G64gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(G57gat), .B2(G64gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n505), .A2(new_n506), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n499), .B1(new_n500), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(new_n314), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n508), .A2(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(KEYINPUT21), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n521), .B(G183gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n524), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G231gat), .A2(G233gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n526), .A2(new_n528), .A3(G231gat), .A4(G233gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G127gat), .B(G155gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G211gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n537));
  INV_X1    g336(.A(new_n535), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n531), .A2(new_n538), .A3(new_n532), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n537), .B1(new_n536), .B2(new_n539), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543));
  INV_X1    g342(.A(G85gat), .ZN(new_n544));
  INV_X1    g343(.A(G92gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(KEYINPUT8), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(KEYINPUT93), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G99gat), .B(G106gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n551), .A2(KEYINPUT95), .A3(new_n553), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n546), .A2(new_n552), .A3(new_n549), .A4(new_n550), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(KEYINPUT96), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n556), .A2(new_n557), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n559), .B(KEYINPUT94), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n562), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G43gat), .B(G50gat), .Z(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT85), .ZN(new_n570));
  XNOR2_X1  g369(.A(G43gat), .B(G50gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT85), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(KEYINPUT15), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G29gat), .A2(G36gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n577));
  OR3_X1    g376(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n569), .A2(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n574), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT86), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n581), .A3(new_n577), .ZN(new_n582));
  OAI211_X1 g381(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n582), .A2(new_n583), .A3(new_n575), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n580), .B1(new_n574), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n574), .A2(new_n575), .A3(new_n579), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n584), .A2(new_n574), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n562), .A2(new_n567), .A3(new_n563), .A4(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n586), .A2(new_n587), .A3(new_n591), .A4(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n595), .A2(KEYINPUT97), .A3(new_n596), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n599), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n600), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n481), .A2(new_n542), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT96), .B1(new_n558), .B2(new_n561), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n565), .A2(new_n566), .A3(new_n564), .ZN(new_n611));
  OAI211_X1 g410(.A(KEYINPUT10), .B(new_n523), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n520), .B1(new_n565), .B2(new_n566), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n551), .A2(KEYINPUT98), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n546), .A2(new_n616), .A3(new_n549), .A4(new_n550), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n553), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n561), .A2(new_n523), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n612), .A2(KEYINPUT99), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622));
  INV_X1    g421(.A(new_n620), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n523), .A2(KEYINPUT10), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n624), .B1(new_n562), .B2(new_n567), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n622), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n621), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n613), .B2(new_n619), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  INV_X1    g430(.A(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT100), .B(G176gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n628), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n627), .B(KEYINPUT101), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n639), .B1(new_n612), .B2(new_n620), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n635), .B1(new_n640), .B2(new_n629), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT102), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n637), .A2(new_n644), .A3(new_n641), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G229gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT90), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n563), .B1(new_n499), .B2(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n649), .A2(new_n590), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT90), .B1(new_n590), .B2(KEYINPUT17), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n651), .A2(new_n499), .ZN(new_n652));
  OAI211_X1 g451(.A(KEYINPUT18), .B(new_n647), .C1(new_n650), .C2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT18), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n649), .A2(new_n590), .B1(new_n651), .B2(new_n499), .ZN(new_n655));
  INV_X1    g454(.A(new_n647), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n499), .B(new_n590), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n647), .B(KEYINPUT13), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n653), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G169gat), .B(G197gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G113gat), .B(G141gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n653), .A2(new_n657), .A3(new_n668), .A4(new_n660), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n646), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n609), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n428), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n486), .ZN(G1324gat));
  NOR2_X1   g476(.A1(new_n675), .A2(new_n421), .ZN(new_n678));
  NAND2_X1  g477(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n679));
  OR2_X1    g478(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  INV_X1    g483(.A(G8gat), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n683), .B(new_n684), .C1(new_n685), .C2(new_n678), .ZN(G1325gat));
  INV_X1    g485(.A(new_n445), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n675), .A2(new_n482), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n675), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n357), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n482), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n397), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n480), .A2(new_n446), .ZN(new_n695));
  INV_X1    g494(.A(new_n441), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n607), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n540), .A2(new_n541), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(new_n673), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(G29gat), .A3(new_n428), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT45), .Z(new_n702));
  NAND2_X1  g501(.A1(new_n697), .A2(KEYINPUT44), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n481), .B2(new_n607), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n699), .B(KEYINPUT103), .Z(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n428), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n702), .A2(new_n709), .ZN(G1328gat));
  NOR3_X1   g509(.A1(new_n700), .A2(G36gat), .A3(new_n421), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT46), .ZN(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n708), .B2(new_n421), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1329gat));
  OAI21_X1  g513(.A(G43gat), .B1(new_n708), .B2(new_n687), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n700), .A2(G43gat), .A3(new_n442), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n715), .B2(new_n717), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(G1330gat));
  NAND2_X1  g519(.A1(new_n435), .A2(G50gat), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n700), .A2(new_n397), .ZN(new_n722));
  OAI22_X1  g521(.A1(new_n708), .A2(new_n721), .B1(G50gat), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g523(.A1(new_n646), .A2(new_n672), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n609), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n428), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g529(.A(new_n420), .B(KEYINPUT104), .Z(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  AND2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n733), .B2(new_n734), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n726), .B2(new_n442), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n726), .A2(new_n738), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n740), .A2(KEYINPUT105), .A3(new_n445), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT105), .B1(new_n740), .B2(new_n445), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n739), .B(new_n744), .C1(new_n741), .C2(new_n742), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1334gat));
  NOR2_X1   g547(.A1(new_n726), .A2(new_n397), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT107), .B(G78gat), .Z(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1335gat));
  NOR3_X1   g550(.A1(new_n428), .A2(G85gat), .A3(new_n646), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n672), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n540), .B2(new_n541), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT51), .B1(new_n697), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n481), .A2(new_n758), .A3(new_n607), .A4(new_n755), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT109), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n695), .A2(new_n696), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n608), .A3(new_n756), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n758), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n697), .A2(KEYINPUT51), .A3(new_n756), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n767), .A2(KEYINPUT108), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n770), .A3(new_n762), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n753), .B1(new_n764), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n646), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n703), .A2(new_n705), .A3(new_n773), .A4(new_n756), .ZN(new_n774));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774), .B2(new_n428), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT110), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n769), .A2(new_n770), .A3(new_n762), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n770), .B1(new_n769), .B2(new_n762), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n752), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n780), .A2(new_n781), .A3(new_n775), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n777), .A2(new_n782), .ZN(G1336gat));
  NOR3_X1   g582(.A1(new_n732), .A2(new_n646), .A3(G92gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n762), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  OAI21_X1  g585(.A(G92gat), .B1(new_n774), .B2(new_n732), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(KEYINPUT111), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(KEYINPUT111), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n774), .A2(new_n421), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n767), .A2(new_n768), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n791), .A2(G92gat), .B1(new_n792), .B2(new_n784), .ZN(new_n793));
  OAI22_X1  g592(.A1(new_n789), .A2(new_n790), .B1(new_n786), .B2(new_n793), .ZN(G1337gat));
  NOR3_X1   g593(.A1(new_n646), .A2(G99gat), .A3(new_n442), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT112), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n778), .B2(new_n779), .ZN(new_n797));
  OAI21_X1  g596(.A(G99gat), .B1(new_n774), .B2(new_n687), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1338gat));
  NOR3_X1   g598(.A1(new_n646), .A2(G106gat), .A3(new_n397), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n769), .A2(new_n762), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  OAI21_X1  g601(.A(G106gat), .B1(new_n774), .B2(new_n397), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n792), .A2(new_n800), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n806), .B2(new_n802), .ZN(G1339gat));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n636), .B1(new_n640), .B2(new_n808), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n621), .A2(new_n626), .A3(new_n627), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n612), .A2(new_n620), .A3(new_n639), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT54), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n809), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(KEYINPUT55), .B(new_n809), .C1(new_n810), .C2(new_n812), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n815), .A2(new_n816), .A3(new_n637), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n655), .A2(new_n656), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n658), .A2(new_n659), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n666), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n671), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n608), .A2(new_n817), .A3(KEYINPUT113), .A4(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n605), .A3(new_n606), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n815), .A2(new_n816), .A3(new_n637), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n672), .A2(new_n815), .A3(new_n816), .A4(new_n637), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n643), .A2(new_n821), .A3(new_n645), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n608), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n542), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n698), .A2(new_n646), .A3(new_n754), .A4(new_n607), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n439), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT82), .B1(new_n438), .B2(new_n397), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(new_n728), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n731), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n205), .A3(new_n672), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n831), .A2(new_n832), .ZN(new_n843));
  INV_X1    g642(.A(new_n398), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n731), .A2(new_n428), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n672), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT114), .B1(new_n848), .B2(G113gat), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n848), .A2(KEYINPUT114), .A3(G113gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n842), .B1(new_n849), .B2(new_n850), .ZN(G1340gat));
  OAI211_X1 g650(.A(new_n841), .B(new_n773), .C1(new_n210), .C2(new_n211), .ZN(new_n852));
  INV_X1    g651(.A(new_n847), .ZN(new_n853));
  OAI21_X1  g652(.A(G120gat), .B1(new_n853), .B2(new_n646), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1341gat));
  NAND2_X1  g654(.A1(new_n841), .A2(new_n698), .ZN(new_n856));
  INV_X1    g655(.A(G127gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n847), .A2(G127gat), .A3(new_n698), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT116), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n847), .A2(new_n861), .A3(G127gat), .A4(new_n698), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n858), .A2(KEYINPUT117), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866));
  AOI21_X1  g665(.A(G127gat), .B1(new_n841), .B2(new_n698), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n863), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n868), .ZN(G1342gat));
  NAND2_X1  g668(.A1(new_n839), .A2(new_n840), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n607), .A2(new_n420), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n218), .A3(new_n871), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n853), .B2(new_n607), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  NOR2_X1   g675(.A1(new_n846), .A2(new_n445), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n828), .A2(new_n879), .A3(new_n829), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n828), .B2(new_n829), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n880), .A2(new_n881), .A3(new_n608), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n542), .B1(new_n882), .B2(new_n827), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT119), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n885), .B(new_n542), .C1(new_n882), .C2(new_n827), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n832), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(KEYINPUT57), .A3(new_n435), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n833), .A2(new_n435), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n878), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n232), .B1(new_n892), .B2(new_n672), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n843), .A2(new_n428), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n445), .A2(new_n397), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n731), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n232), .A3(new_n672), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT58), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n754), .B(new_n878), .C1(new_n888), .C2(new_n891), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n901), .B(new_n898), .C1(new_n902), .C2(new_n232), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(G1344gat));
  AOI211_X1 g703(.A(KEYINPUT59), .B(new_n230), .C1(new_n892), .C2(new_n773), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n824), .A2(new_n825), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n542), .B1(new_n882), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n832), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(KEYINPUT122), .A3(new_n832), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n911), .A2(new_n890), .A3(new_n435), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n889), .A2(KEYINPUT57), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n877), .B(KEYINPUT121), .Z(new_n915));
  NAND4_X1  g714(.A1(new_n913), .A2(new_n914), .A3(new_n773), .A4(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n906), .B1(new_n916), .B2(G148gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n897), .A2(new_n230), .A3(new_n773), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n905), .A2(new_n917), .B1(new_n920), .B2(new_n921), .ZN(G1345gat));
  AOI21_X1  g721(.A(G155gat), .B1(new_n897), .B2(new_n698), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n542), .A2(new_n223), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n892), .B2(new_n924), .ZN(G1346gat));
  NAND2_X1  g724(.A1(new_n888), .A2(new_n891), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n608), .A3(new_n877), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n892), .A2(KEYINPUT123), .A3(new_n608), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(G162gat), .A3(new_n930), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n894), .A2(new_n224), .A3(new_n871), .A4(new_n895), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1347gat));
  NAND2_X1  g732(.A1(new_n428), .A2(new_n420), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT125), .Z(new_n935));
  NAND3_X1  g734(.A1(new_n833), .A2(new_n398), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(G169gat), .B1(new_n936), .B2(new_n754), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n843), .A2(new_n732), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n428), .A3(new_n836), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT124), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n938), .A2(new_n941), .A3(new_n428), .A4(new_n836), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n672), .B1(new_n309), .B2(new_n308), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n937), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n947), .B(new_n937), .C1(new_n943), .C2(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1348gat));
  NOR3_X1   g748(.A1(new_n936), .A2(new_n294), .A3(new_n646), .ZN(new_n950));
  INV_X1    g749(.A(new_n943), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n773), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n952), .B2(new_n294), .ZN(G1349gat));
  OAI21_X1  g752(.A(G183gat), .B1(new_n936), .B2(new_n542), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n698), .B1(new_n286), .B2(new_n285), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n939), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g756(.A1(new_n951), .A2(new_n284), .A3(new_n608), .ZN(new_n958));
  OAI21_X1  g757(.A(G190gat), .B1(new_n936), .B2(new_n607), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(KEYINPUT61), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n959), .A2(KEYINPUT61), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G1351gat));
  AND3_X1   g761(.A1(new_n938), .A2(new_n428), .A3(new_n895), .ZN(new_n963));
  INV_X1    g762(.A(G197gat), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(new_n964), .A3(new_n672), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n913), .A2(new_n914), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n935), .A2(new_n687), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n966), .A2(new_n672), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n965), .B1(new_n968), .B2(new_n964), .ZN(G1352gat));
  NAND3_X1  g768(.A1(new_n963), .A2(new_n632), .A3(new_n773), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n966), .A2(new_n773), .A3(new_n967), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n971), .B(new_n972), .C1(new_n973), .C2(new_n632), .ZN(G1353gat));
  NAND3_X1  g773(.A1(new_n963), .A2(new_n360), .A3(new_n698), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n913), .A2(new_n914), .A3(new_n698), .A4(new_n967), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n361), .A3(new_n608), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n966), .A2(new_n608), .A3(new_n967), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n981), .B2(new_n361), .ZN(G1355gat));
endmodule


