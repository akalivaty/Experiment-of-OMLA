

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758;

  AND2_X1 U369 ( .A1(n657), .A2(n608), .ZN(n612) );
  INV_X1 U370 ( .A(KEYINPUT40), .ZN(n349) );
  NOR2_X1 U371 ( .A1(n567), .A2(n376), .ZN(n569) );
  AND2_X1 U372 ( .A1(n418), .A2(n395), .ZN(n565) );
  OR2_X1 U373 ( .A1(n720), .A2(G902), .ZN(n388) );
  XNOR2_X1 U374 ( .A(n470), .B(G107), .ZN(n484) );
  XNOR2_X1 U375 ( .A(n452), .B(G113), .ZN(n483) );
  INV_X1 U376 ( .A(G116), .ZN(n470) );
  INV_X1 U377 ( .A(KEYINPUT68), .ZN(n397) );
  NAND2_X1 U378 ( .A1(n535), .A2(n513), .ZN(n514) );
  XNOR2_X2 U379 ( .A(n400), .B(n512), .ZN(n535) );
  AND2_X2 U380 ( .A1(n368), .A2(n365), .ZN(n364) );
  NAND2_X2 U381 ( .A1(n364), .A2(n362), .ZN(n370) );
  XNOR2_X2 U382 ( .A(n350), .B(n349), .ZN(n754) );
  NAND2_X1 U383 ( .A1(n602), .A2(n650), .ZN(n350) );
  INV_X1 U384 ( .A(n575), .ZN(n650) );
  AND2_X4 U385 ( .A1(n612), .A2(n611), .ZN(n714) );
  INV_X2 U386 ( .A(KEYINPUT66), .ZN(n432) );
  NOR2_X2 U387 ( .A1(n515), .A2(n517), .ZN(n516) );
  NOR2_X1 U388 ( .A1(n650), .A2(n652), .ZN(n542) );
  XOR2_X1 U389 ( .A(G472), .B(n521), .Z(n682) );
  INV_X2 U390 ( .A(G953), .ZN(n743) );
  NOR2_X1 U391 ( .A1(n533), .A2(n750), .ZN(n534) );
  NAND2_X1 U392 ( .A1(n407), .A2(n404), .ZN(n633) );
  NAND2_X1 U393 ( .A1(n391), .A2(n356), .ZN(n646) );
  NOR2_X1 U394 ( .A1(n556), .A2(n450), .ZN(n451) );
  AND2_X1 U395 ( .A1(n371), .A2(n359), .ZN(n374) );
  XNOR2_X1 U396 ( .A(n521), .B(n520), .ZN(n566) );
  XNOR2_X1 U397 ( .A(n401), .B(KEYINPUT19), .ZN(n582) );
  XNOR2_X1 U398 ( .A(n402), .B(n487), .ZN(n726) );
  XNOR2_X1 U399 ( .A(n483), .B(n484), .ZN(n402) );
  XNOR2_X1 U400 ( .A(KEYINPUT3), .B(G119), .ZN(n486) );
  XNOR2_X1 U401 ( .A(KEYINPUT70), .B(KEYINPUT16), .ZN(n485) );
  INV_X1 U402 ( .A(n607), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n551), .B(n550), .ZN(n729) );
  NAND2_X1 U404 ( .A1(n374), .A2(n372), .ZN(n376) );
  OR2_X1 U405 ( .A1(n610), .A2(KEYINPUT2), .ZN(n611) );
  OR2_X2 U406 ( .A1(n754), .A2(n386), .ZN(n385) );
  XNOR2_X1 U407 ( .A(n422), .B(G125), .ZN(n492) );
  INV_X1 U408 ( .A(G146), .ZN(n422) );
  INV_X1 U409 ( .A(n522), .ZN(n411) );
  XNOR2_X1 U410 ( .A(n464), .B(n438), .ZN(n739) );
  XNOR2_X1 U411 ( .A(n591), .B(KEYINPUT81), .ZN(n387) );
  NAND2_X1 U412 ( .A1(n380), .A2(n384), .ZN(n382) );
  AND2_X1 U413 ( .A1(n366), .A2(n751), .ZN(n365) );
  NAND2_X1 U414 ( .A1(n367), .A2(KEYINPUT48), .ZN(n366) );
  INV_X1 U415 ( .A(n387), .ZN(n367) );
  INV_X1 U416 ( .A(n633), .ZN(n360) );
  XOR2_X1 U417 ( .A(G137), .B(G140), .Z(n438) );
  INV_X1 U418 ( .A(G107), .ZN(n436) );
  INV_X1 U419 ( .A(KEYINPUT30), .ZN(n375) );
  OR2_X1 U420 ( .A1(n566), .A2(n354), .ZN(n372) );
  INV_X1 U421 ( .A(n665), .ZN(n373) );
  XNOR2_X1 U422 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U423 ( .A(n423), .B(n415), .ZN(n414) );
  XNOR2_X1 U424 ( .A(G128), .B(G119), .ZN(n423) );
  XNOR2_X1 U425 ( .A(n416), .B(KEYINPUT24), .ZN(n415) );
  INV_X1 U426 ( .A(KEYINPUT92), .ZN(n416) );
  XNOR2_X1 U427 ( .A(n421), .B(n492), .ZN(n464) );
  NAND2_X1 U428 ( .A1(n390), .A2(KEYINPUT78), .ZN(n389) );
  INV_X1 U429 ( .A(n583), .ZN(n390) );
  NAND2_X1 U430 ( .A1(n584), .A2(n394), .ZN(n393) );
  NAND2_X1 U431 ( .A1(n517), .A2(KEYINPUT101), .ZN(n410) );
  NAND2_X1 U432 ( .A1(n409), .A2(KEYINPUT101), .ZN(n408) );
  OR2_X2 U433 ( .A1(n708), .A2(G902), .ZN(n420) );
  XOR2_X1 U434 ( .A(KEYINPUT5), .B(G137), .Z(n446) );
  XNOR2_X1 U435 ( .A(G116), .B(G113), .ZN(n445) );
  XNOR2_X1 U436 ( .A(n370), .B(KEYINPUT85), .ZN(n609) );
  XNOR2_X1 U437 ( .A(n525), .B(KEYINPUT72), .ZN(n399) );
  AND2_X1 U438 ( .A1(n685), .A2(n524), .ZN(n525) );
  NAND2_X1 U439 ( .A1(n558), .A2(n355), .ZN(n419) );
  XNOR2_X1 U440 ( .A(n519), .B(n518), .ZN(n520) );
  AND2_X1 U441 ( .A1(n677), .A2(n355), .ZN(n557) );
  BUF_X1 U442 ( .A(n658), .Z(n742) );
  NAND2_X1 U443 ( .A1(n435), .A2(n434), .ZN(n379) );
  XOR2_X1 U444 ( .A(G140), .B(KEYINPUT12), .Z(n456) );
  INV_X1 U445 ( .A(G122), .ZN(n452) );
  XNOR2_X1 U446 ( .A(n440), .B(n488), .ZN(n441) );
  XNOR2_X1 U447 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U448 ( .A(n437), .B(n436), .ZN(n439) );
  NAND2_X1 U449 ( .A1(n582), .A2(n510), .ZN(n400) );
  XNOR2_X1 U450 ( .A(n426), .B(n413), .ZN(n412) );
  XNOR2_X1 U451 ( .A(n424), .B(n414), .ZN(n413) );
  XNOR2_X1 U452 ( .A(n498), .B(n497), .ZN(n615) );
  XNOR2_X1 U453 ( .A(n726), .B(n488), .ZN(n498) );
  XNOR2_X1 U454 ( .A(n532), .B(KEYINPUT35), .ZN(n750) );
  AND2_X1 U455 ( .A1(n393), .A2(n392), .ZN(n391) );
  NAND2_X1 U456 ( .A1(n583), .A2(n394), .ZN(n392) );
  NAND2_X1 U457 ( .A1(n406), .A2(n405), .ZN(n404) );
  AND2_X1 U458 ( .A1(n410), .A2(n408), .ZN(n407) );
  NOR2_X1 U459 ( .A1(n684), .A2(n352), .ZN(n405) );
  OR2_X1 U460 ( .A1(n411), .A2(KEYINPUT101), .ZN(n352) );
  XOR2_X1 U461 ( .A(KEYINPUT69), .B(G469), .Z(n353) );
  OR2_X1 U462 ( .A1(n373), .A2(KEYINPUT30), .ZN(n354) );
  OR2_X1 U463 ( .A1(n555), .A2(n554), .ZN(n355) );
  OR2_X1 U464 ( .A1(n584), .A2(n389), .ZN(n356) );
  AND2_X1 U465 ( .A1(n595), .A2(n656), .ZN(n357) );
  AND2_X1 U466 ( .A1(n406), .A2(n403), .ZN(n358) );
  OR2_X1 U467 ( .A1(n665), .A2(n375), .ZN(n359) );
  INV_X1 U468 ( .A(KEYINPUT78), .ZN(n394) );
  XNOR2_X1 U469 ( .A(n412), .B(n739), .ZN(n720) );
  INV_X1 U470 ( .A(KEYINPUT48), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n396), .B(n441), .ZN(n708) );
  NAND2_X1 U472 ( .A1(n361), .A2(n360), .ZN(n523) );
  INV_X1 U473 ( .A(n753), .ZN(n361) );
  NAND2_X1 U474 ( .A1(n363), .A2(KEYINPUT48), .ZN(n362) );
  INV_X1 U475 ( .A(n381), .ZN(n363) );
  NAND2_X1 U476 ( .A1(n381), .A2(n369), .ZN(n368) );
  AND2_X1 U477 ( .A1(n387), .A2(n417), .ZN(n369) );
  NAND2_X1 U478 ( .A1(n566), .A2(KEYINPUT30), .ZN(n371) );
  XNOR2_X2 U479 ( .A(n741), .B(G146), .ZN(n396) );
  XNOR2_X2 U480 ( .A(n476), .B(n377), .ZN(n741) );
  XNOR2_X2 U481 ( .A(n453), .B(n494), .ZN(n377) );
  NAND2_X1 U482 ( .A1(n379), .A2(n378), .ZN(n476) );
  NAND2_X1 U483 ( .A1(n493), .A2(G134), .ZN(n378) );
  NAND2_X1 U484 ( .A1(n754), .A2(KEYINPUT46), .ZN(n380) );
  NOR2_X2 U485 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U486 ( .A1(n357), .A2(n385), .ZN(n383) );
  NAND2_X1 U487 ( .A1(n758), .A2(KEYINPUT46), .ZN(n384) );
  OR2_X1 U488 ( .A1(n758), .A2(KEYINPUT46), .ZN(n386) );
  INV_X1 U489 ( .A(n677), .ZN(n556) );
  XNOR2_X2 U490 ( .A(n388), .B(n431), .ZN(n677) );
  NAND2_X1 U491 ( .A1(n646), .A2(n592), .ZN(n585) );
  NAND2_X1 U492 ( .A1(n560), .A2(n395), .ZN(n584) );
  NAND2_X1 U493 ( .A1(n685), .A2(n395), .ZN(n564) );
  XNOR2_X1 U494 ( .A(n395), .B(KEYINPUT1), .ZN(n524) );
  XNOR2_X2 U495 ( .A(n420), .B(n353), .ZN(n395) );
  XNOR2_X1 U496 ( .A(n396), .B(n449), .ZN(n627) );
  XNOR2_X2 U497 ( .A(n397), .B(G131), .ZN(n453) );
  NAND2_X1 U498 ( .A1(n399), .A2(n398), .ZN(n526) );
  INV_X1 U499 ( .A(n574), .ZN(n398) );
  AND2_X1 U500 ( .A1(n399), .A2(n682), .ZN(n690) );
  XNOR2_X2 U501 ( .A(n542), .B(KEYINPUT99), .ZN(n592) );
  XNOR2_X2 U502 ( .A(n432), .B(KEYINPUT4), .ZN(n494) );
  NAND2_X1 U503 ( .A1(n599), .A2(n665), .ZN(n401) );
  INV_X1 U504 ( .A(n684), .ZN(n403) );
  INV_X1 U505 ( .A(n517), .ZN(n406) );
  OR2_X1 U506 ( .A1(n684), .A2(n411), .ZN(n409) );
  XNOR2_X2 U507 ( .A(n514), .B(KEYINPUT22), .ZN(n517) );
  NOR2_X1 U508 ( .A1(n677), .A2(n419), .ZN(n418) );
  NOR2_X1 U509 ( .A1(n677), .A2(n676), .ZN(n685) );
  NAND2_X1 U510 ( .A1(n607), .A2(n606), .ZN(n657) );
  XOR2_X1 U511 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n421) );
  INV_X1 U512 ( .A(G472), .ZN(n518) );
  XNOR2_X1 U513 ( .A(n448), .B(n447), .ZN(n449) );
  INV_X1 U514 ( .A(KEYINPUT74), .ZN(n568) );
  BUF_X1 U515 ( .A(n524), .Z(n684) );
  INV_X1 U516 ( .A(KEYINPUT63), .ZN(n631) );
  INV_X1 U517 ( .A(KEYINPUT123), .ZN(n624) );
  XOR2_X1 U518 ( .A(KEYINPUT23), .B(G110), .Z(n424) );
  NAND2_X1 U519 ( .A1(G234), .A2(n743), .ZN(n425) );
  XOR2_X1 U520 ( .A(KEYINPUT8), .B(n425), .Z(n471) );
  NAND2_X1 U521 ( .A1(n471), .A2(G221), .ZN(n426) );
  INV_X1 U522 ( .A(KEYINPUT15), .ZN(n427) );
  XNOR2_X1 U523 ( .A(n427), .B(G902), .ZN(n608) );
  INV_X1 U524 ( .A(n608), .ZN(n499) );
  NAND2_X1 U525 ( .A1(G234), .A2(n499), .ZN(n428) );
  XNOR2_X1 U526 ( .A(KEYINPUT20), .B(n428), .ZN(n479) );
  NAND2_X1 U527 ( .A1(G217), .A2(n479), .ZN(n430) );
  XOR2_X1 U528 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n429) );
  INV_X2 U529 ( .A(G143), .ZN(n433) );
  XNOR2_X2 U530 ( .A(n433), .B(G128), .ZN(n493) );
  INV_X1 U531 ( .A(n493), .ZN(n435) );
  INV_X1 U532 ( .A(G134), .ZN(n434) );
  NAND2_X1 U533 ( .A1(G227), .A2(n743), .ZN(n437) );
  XOR2_X1 U534 ( .A(KEYINPUT65), .B(G101), .Z(n443) );
  XNOR2_X1 U535 ( .A(G110), .B(G104), .ZN(n724) );
  XNOR2_X1 U536 ( .A(n443), .B(n724), .ZN(n488) );
  NOR2_X2 U537 ( .A1(G953), .A2(G237), .ZN(n454) );
  NAND2_X1 U538 ( .A1(n454), .A2(G210), .ZN(n442) );
  XOR2_X1 U539 ( .A(n486), .B(n442), .Z(n444) );
  XNOR2_X1 U540 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U541 ( .A(n446), .B(n445), .Z(n447) );
  NOR2_X2 U542 ( .A1(G902), .A2(n627), .ZN(n521) );
  XNOR2_X1 U543 ( .A(n682), .B(KEYINPUT6), .ZN(n574) );
  NAND2_X1 U544 ( .A1(n684), .A2(n574), .ZN(n450) );
  XNOR2_X1 U545 ( .A(n451), .B(KEYINPUT77), .ZN(n515) );
  XNOR2_X1 U546 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n466) );
  XNOR2_X1 U547 ( .A(n453), .B(n483), .ZN(n462) );
  NAND2_X1 U548 ( .A1(n454), .A2(G214), .ZN(n455) );
  XNOR2_X1 U549 ( .A(n456), .B(n455), .ZN(n460) );
  XOR2_X1 U550 ( .A(KEYINPUT11), .B(KEYINPUT95), .Z(n458) );
  XNOR2_X1 U551 ( .A(G143), .B(G104), .ZN(n457) );
  XNOR2_X1 U552 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U553 ( .A(n460), .B(n459), .Z(n461) );
  XNOR2_X1 U554 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U555 ( .A(n464), .B(n463), .ZN(n715) );
  NOR2_X1 U556 ( .A1(G902), .A2(n715), .ZN(n465) );
  XNOR2_X1 U557 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U558 ( .A(G475), .B(n467), .ZN(n540) );
  INV_X1 U559 ( .A(n540), .ZN(n529) );
  XOR2_X1 U560 ( .A(KEYINPUT97), .B(KEYINPUT9), .Z(n469) );
  XNOR2_X1 U561 ( .A(G122), .B(KEYINPUT98), .ZN(n468) );
  XNOR2_X1 U562 ( .A(n469), .B(n468), .ZN(n475) );
  XOR2_X1 U563 ( .A(n484), .B(KEYINPUT7), .Z(n473) );
  NAND2_X1 U564 ( .A1(G217), .A2(n471), .ZN(n472) );
  XNOR2_X1 U565 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U566 ( .A(n475), .B(n474), .ZN(n477) );
  XOR2_X1 U567 ( .A(n477), .B(n476), .Z(n621) );
  NOR2_X1 U568 ( .A1(n621), .A2(G902), .ZN(n478) );
  XNOR2_X1 U569 ( .A(G478), .B(n478), .ZN(n541) );
  NAND2_X1 U570 ( .A1(n529), .A2(n541), .ZN(n669) );
  NAND2_X1 U571 ( .A1(n479), .A2(G221), .ZN(n480) );
  XNOR2_X1 U572 ( .A(n480), .B(KEYINPUT94), .ZN(n482) );
  INV_X1 U573 ( .A(KEYINPUT21), .ZN(n481) );
  XNOR2_X1 U574 ( .A(n482), .B(n481), .ZN(n558) );
  INV_X1 U575 ( .A(n558), .ZN(n676) );
  NOR2_X1 U576 ( .A1(n669), .A2(n676), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U578 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n490) );
  NAND2_X1 U579 ( .A1(n743), .A2(G224), .ZN(n489) );
  XNOR2_X1 U580 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U581 ( .A(n492), .B(n491), .ZN(n496) );
  XNOR2_X1 U582 ( .A(n493), .B(n494), .ZN(n495) );
  XNOR2_X1 U583 ( .A(n496), .B(n495), .ZN(n497) );
  NAND2_X1 U584 ( .A1(n615), .A2(n499), .ZN(n503) );
  NOR2_X1 U585 ( .A1(G237), .A2(G902), .ZN(n500) );
  XNOR2_X1 U586 ( .A(n500), .B(KEYINPUT73), .ZN(n504) );
  NAND2_X1 U587 ( .A1(n504), .A2(G210), .ZN(n501) );
  XNOR2_X1 U588 ( .A(n501), .B(KEYINPUT79), .ZN(n502) );
  XNOR2_X2 U589 ( .A(n503), .B(n502), .ZN(n599) );
  NAND2_X1 U590 ( .A1(n504), .A2(G214), .ZN(n665) );
  NAND2_X1 U591 ( .A1(G237), .A2(G234), .ZN(n505) );
  XNOR2_X1 U592 ( .A(n505), .B(KEYINPUT88), .ZN(n506) );
  XNOR2_X1 U593 ( .A(KEYINPUT14), .B(n506), .ZN(n507) );
  NAND2_X1 U594 ( .A1(G952), .A2(n507), .ZN(n699) );
  NOR2_X1 U595 ( .A1(G953), .A2(n699), .ZN(n555) );
  NAND2_X1 U596 ( .A1(n507), .A2(G902), .ZN(n552) );
  XNOR2_X1 U597 ( .A(KEYINPUT89), .B(G898), .ZN(n732) );
  NAND2_X1 U598 ( .A1(G953), .A2(n732), .ZN(n727) );
  NOR2_X1 U599 ( .A1(n552), .A2(n727), .ZN(n508) );
  OR2_X1 U600 ( .A1(n555), .A2(n508), .ZN(n509) );
  XNOR2_X1 U601 ( .A(n509), .B(KEYINPUT90), .ZN(n510) );
  INV_X1 U602 ( .A(KEYINPUT64), .ZN(n511) );
  XNOR2_X1 U603 ( .A(n511), .B(KEYINPUT0), .ZN(n512) );
  XNOR2_X1 U604 ( .A(n516), .B(KEYINPUT32), .ZN(n753) );
  INV_X1 U605 ( .A(KEYINPUT100), .ZN(n519) );
  AND2_X1 U606 ( .A1(n566), .A2(n677), .ZN(n522) );
  XNOR2_X1 U607 ( .A(n523), .B(KEYINPUT86), .ZN(n533) );
  XOR2_X1 U608 ( .A(KEYINPUT102), .B(KEYINPUT33), .Z(n527) );
  XNOR2_X1 U609 ( .A(n527), .B(n526), .ZN(n700) );
  XNOR2_X1 U610 ( .A(n535), .B(KEYINPUT91), .ZN(n538) );
  NOR2_X1 U611 ( .A1(n700), .A2(n538), .ZN(n528) );
  XNOR2_X1 U612 ( .A(n528), .B(KEYINPUT34), .ZN(n531) );
  OR2_X1 U613 ( .A1(n541), .A2(n529), .ZN(n587) );
  XOR2_X1 U614 ( .A(n587), .B(KEYINPUT76), .Z(n530) );
  NAND2_X1 U615 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U616 ( .A(n534), .B(KEYINPUT44), .ZN(n548) );
  AND2_X1 U617 ( .A1(n535), .A2(n690), .ZN(n537) );
  INV_X1 U618 ( .A(KEYINPUT31), .ZN(n536) );
  XNOR2_X1 U619 ( .A(n537), .B(n536), .ZN(n653) );
  OR2_X1 U620 ( .A1(n682), .A2(n538), .ZN(n539) );
  NOR2_X1 U621 ( .A1(n564), .A2(n539), .ZN(n639) );
  OR2_X1 U622 ( .A1(n653), .A2(n639), .ZN(n543) );
  NAND2_X1 U623 ( .A1(n541), .A2(n540), .ZN(n575) );
  NOR2_X1 U624 ( .A1(n541), .A2(n540), .ZN(n652) );
  NAND2_X1 U625 ( .A1(n543), .A2(n592), .ZN(n546) );
  AND2_X1 U626 ( .A1(n574), .A2(n556), .ZN(n544) );
  AND2_X1 U627 ( .A1(n358), .A2(n544), .ZN(n636) );
  INV_X1 U628 ( .A(n636), .ZN(n545) );
  AND2_X1 U629 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U630 ( .A1(n548), .A2(n547), .ZN(n551) );
  INV_X1 U631 ( .A(KEYINPUT84), .ZN(n549) );
  XNOR2_X1 U632 ( .A(n549), .B(KEYINPUT45), .ZN(n550) );
  INV_X1 U633 ( .A(n729), .ZN(n607) );
  OR2_X1 U634 ( .A1(n743), .A2(n552), .ZN(n553) );
  NOR2_X1 U635 ( .A1(G900), .A2(n553), .ZN(n554) );
  NAND2_X1 U636 ( .A1(n558), .A2(n557), .ZN(n578) );
  NOR2_X1 U637 ( .A1(n566), .A2(n578), .ZN(n559) );
  XNOR2_X1 U638 ( .A(n559), .B(KEYINPUT28), .ZN(n560) );
  XNOR2_X1 U639 ( .A(n599), .B(KEYINPUT38), .ZN(n570) );
  INV_X1 U640 ( .A(n570), .ZN(n666) );
  NAND2_X1 U641 ( .A1(n666), .A2(n665), .ZN(n670) );
  NOR2_X1 U642 ( .A1(n670), .A2(n669), .ZN(n562) );
  XNOR2_X1 U643 ( .A(KEYINPUT104), .B(KEYINPUT41), .ZN(n561) );
  XNOR2_X1 U644 ( .A(n562), .B(n561), .ZN(n701) );
  NOR2_X1 U645 ( .A1(n584), .A2(n701), .ZN(n563) );
  XNOR2_X1 U646 ( .A(n563), .B(KEYINPUT42), .ZN(n758) );
  XNOR2_X1 U647 ( .A(n565), .B(KEYINPUT75), .ZN(n567) );
  XNOR2_X1 U648 ( .A(n569), .B(n568), .ZN(n586) );
  INV_X1 U649 ( .A(n586), .ZN(n571) );
  NAND2_X1 U650 ( .A1(n571), .A2(n666), .ZN(n572) );
  XNOR2_X1 U651 ( .A(n572), .B(KEYINPUT39), .ZN(n602) );
  NOR2_X1 U652 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U653 ( .A1(n576), .A2(n665), .ZN(n577) );
  NOR2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n596) );
  NAND2_X1 U655 ( .A1(n596), .A2(n599), .ZN(n579) );
  XNOR2_X1 U656 ( .A(n579), .B(KEYINPUT36), .ZN(n580) );
  XNOR2_X1 U657 ( .A(n580), .B(KEYINPUT105), .ZN(n581) );
  NAND2_X1 U658 ( .A1(n581), .A2(n684), .ZN(n656) );
  INV_X1 U659 ( .A(n582), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n585), .A2(KEYINPUT47), .ZN(n590) );
  NOR2_X1 U661 ( .A1(n586), .A2(n587), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n588), .A2(n599), .ZN(n635) );
  XNOR2_X1 U663 ( .A(n635), .B(KEYINPUT82), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U665 ( .A(n592), .ZN(n671) );
  NOR2_X1 U666 ( .A1(KEYINPUT47), .A2(n671), .ZN(n593) );
  XOR2_X1 U667 ( .A(KEYINPUT71), .B(n593), .Z(n594) );
  NAND2_X1 U668 ( .A1(n594), .A2(n646), .ZN(n595) );
  INV_X1 U669 ( .A(n596), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n684), .A2(n597), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT43), .ZN(n600) );
  NOR2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U673 ( .A(n601), .B(KEYINPUT103), .ZN(n751) );
  NAND2_X1 U674 ( .A1(n652), .A2(n602), .ZN(n603) );
  XNOR2_X1 U675 ( .A(KEYINPUT106), .B(n603), .ZN(n756) );
  NAND2_X1 U676 ( .A1(n756), .A2(KEYINPUT2), .ZN(n604) );
  XOR2_X1 U677 ( .A(KEYINPUT80), .B(n604), .Z(n605) );
  AND2_X1 U678 ( .A1(n609), .A2(n605), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n609), .A2(n756), .ZN(n658) );
  NOR2_X1 U680 ( .A1(n658), .A2(n729), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n714), .A2(G210), .ZN(n617) );
  XOR2_X1 U682 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT87), .ZN(n614) );
  XNOR2_X1 U684 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U685 ( .A(n617), .B(n616), .ZN(n619) );
  INV_X1 U686 ( .A(G952), .ZN(n618) );
  AND2_X1 U687 ( .A1(n618), .A2(G953), .ZN(n723) );
  NOR2_X2 U688 ( .A1(n619), .A2(n723), .ZN(n620) );
  XNOR2_X1 U689 ( .A(n620), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U690 ( .A1(n714), .A2(G478), .ZN(n622) );
  XNOR2_X1 U691 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X2 U692 ( .A1(n623), .A2(n723), .ZN(n625) );
  XNOR2_X1 U693 ( .A(n625), .B(n624), .ZN(G63) );
  NAND2_X1 U694 ( .A1(n714), .A2(G472), .ZN(n629) );
  XOR2_X1 U695 ( .A(KEYINPUT107), .B(KEYINPUT62), .Z(n626) );
  XNOR2_X1 U696 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U697 ( .A(n629), .B(n628), .ZN(n630) );
  NOR2_X2 U698 ( .A1(n630), .A2(n723), .ZN(n632) );
  XNOR2_X1 U699 ( .A(n632), .B(n631), .ZN(G57) );
  XOR2_X1 U700 ( .A(G110), .B(n633), .Z(G12) );
  XNOR2_X1 U701 ( .A(G143), .B(KEYINPUT110), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n635), .B(n634), .ZN(G45) );
  XOR2_X1 U703 ( .A(G101), .B(n636), .Z(n637) );
  XNOR2_X1 U704 ( .A(KEYINPUT108), .B(n637), .ZN(G3) );
  NAND2_X1 U705 ( .A1(n639), .A2(n650), .ZN(n638) );
  XNOR2_X1 U706 ( .A(n638), .B(G104), .ZN(G6) );
  XOR2_X1 U707 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n641) );
  NAND2_X1 U708 ( .A1(n639), .A2(n652), .ZN(n640) );
  XNOR2_X1 U709 ( .A(n641), .B(n640), .ZN(n643) );
  XOR2_X1 U710 ( .A(G107), .B(KEYINPUT109), .Z(n642) );
  XNOR2_X1 U711 ( .A(n643), .B(n642), .ZN(G9) );
  XOR2_X1 U712 ( .A(G128), .B(KEYINPUT29), .Z(n645) );
  NAND2_X1 U713 ( .A1(n652), .A2(n646), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n645), .B(n644), .ZN(G30) );
  XOR2_X1 U715 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n648) );
  NAND2_X1 U716 ( .A1(n650), .A2(n646), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U718 ( .A(G146), .B(n649), .ZN(G48) );
  NAND2_X1 U719 ( .A1(n653), .A2(n650), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n651), .B(G113), .ZN(G15) );
  NAND2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n654), .B(G116), .ZN(G18) );
  XOR2_X1 U723 ( .A(G125), .B(KEYINPUT37), .Z(n655) );
  XNOR2_X1 U724 ( .A(n656), .B(n655), .ZN(G27) );
  INV_X1 U725 ( .A(n657), .ZN(n660) );
  INV_X1 U726 ( .A(KEYINPUT2), .ZN(n661) );
  AND2_X1 U727 ( .A1(n661), .A2(n742), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U729 ( .A1(n351), .A2(n661), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT83), .B(n662), .Z(n663) );
  NAND2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n705) );
  NOR2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U733 ( .A(KEYINPUT119), .B(n667), .Z(n668) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n673) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U737 ( .A(n674), .B(KEYINPUT120), .ZN(n675) );
  NOR2_X1 U738 ( .A1(n700), .A2(n675), .ZN(n695) );
  XOR2_X1 U739 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n679) );
  NAND2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U741 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U742 ( .A(n680), .B(KEYINPUT115), .ZN(n681) );
  NOR2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U744 ( .A(KEYINPUT117), .B(n683), .ZN(n688) );
  NOR2_X1 U745 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U746 ( .A(KEYINPUT50), .B(n686), .ZN(n687) );
  NOR2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U749 ( .A(KEYINPUT51), .B(n691), .Z(n692) );
  XNOR2_X1 U750 ( .A(n692), .B(KEYINPUT118), .ZN(n693) );
  NOR2_X1 U751 ( .A1(n701), .A2(n693), .ZN(n694) );
  NOR2_X1 U752 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U753 ( .A(KEYINPUT52), .B(n696), .Z(n697) );
  XNOR2_X1 U754 ( .A(n697), .B(KEYINPUT121), .ZN(n698) );
  NOR2_X1 U755 ( .A1(n699), .A2(n698), .ZN(n703) );
  NOR2_X1 U756 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U757 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U758 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U759 ( .A1(n706), .A2(G953), .ZN(n707) );
  XNOR2_X1 U760 ( .A(n707), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U761 ( .A1(n714), .A2(G469), .ZN(n712) );
  XOR2_X1 U762 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n710) );
  XNOR2_X1 U763 ( .A(n708), .B(KEYINPUT122), .ZN(n709) );
  XNOR2_X1 U764 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n723), .A2(n713), .ZN(G54) );
  NAND2_X1 U767 ( .A1(n714), .A2(G475), .ZN(n717) );
  XOR2_X1 U768 ( .A(n715), .B(KEYINPUT59), .Z(n716) );
  XNOR2_X1 U769 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X2 U770 ( .A1(n718), .A2(n723), .ZN(n719) );
  XNOR2_X1 U771 ( .A(n719), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U772 ( .A1(n714), .A2(G217), .ZN(n721) );
  XNOR2_X1 U773 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U774 ( .A1(n723), .A2(n722), .ZN(G66) );
  XOR2_X1 U775 ( .A(n724), .B(G101), .Z(n725) );
  XNOR2_X1 U776 ( .A(n726), .B(n725), .ZN(n728) );
  NAND2_X1 U777 ( .A1(n728), .A2(n727), .ZN(n738) );
  NOR2_X1 U778 ( .A1(n351), .A2(G953), .ZN(n736) );
  XOR2_X1 U779 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n731) );
  NAND2_X1 U780 ( .A1(G224), .A2(G953), .ZN(n730) );
  XNOR2_X1 U781 ( .A(n731), .B(n730), .ZN(n733) );
  NOR2_X1 U782 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U783 ( .A(KEYINPUT125), .B(n734), .Z(n735) );
  NOR2_X1 U784 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U785 ( .A(n738), .B(n737), .ZN(G69) );
  XNOR2_X1 U786 ( .A(n739), .B(KEYINPUT126), .ZN(n740) );
  XNOR2_X1 U787 ( .A(n741), .B(n740), .ZN(n745) );
  XNOR2_X1 U788 ( .A(n745), .B(n742), .ZN(n744) );
  NAND2_X1 U789 ( .A1(n744), .A2(n743), .ZN(n749) );
  XNOR2_X1 U790 ( .A(G227), .B(n745), .ZN(n746) );
  NAND2_X1 U791 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U792 ( .A1(G953), .A2(n747), .ZN(n748) );
  NAND2_X1 U793 ( .A1(n749), .A2(n748), .ZN(G72) );
  XOR2_X1 U794 ( .A(G122), .B(n750), .Z(G24) );
  XNOR2_X1 U795 ( .A(G140), .B(KEYINPUT114), .ZN(n752) );
  XNOR2_X1 U796 ( .A(n752), .B(n751), .ZN(G42) );
  XOR2_X1 U797 ( .A(n753), .B(G119), .Z(G21) );
  XNOR2_X1 U798 ( .A(G131), .B(KEYINPUT127), .ZN(n755) );
  XNOR2_X1 U799 ( .A(n755), .B(n754), .ZN(G33) );
  XOR2_X1 U800 ( .A(G134), .B(n756), .Z(n757) );
  XNOR2_X1 U801 ( .A(KEYINPUT113), .B(n757), .ZN(G36) );
  XOR2_X1 U802 ( .A(G137), .B(n758), .Z(G39) );
endmodule

