//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  AOI21_X1  g005(.A(G128), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(KEYINPUT1), .A3(G146), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT71), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT71), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n193), .B(new_n196), .C1(new_n197), .C2(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n200), .A3(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G134), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT68), .B(G134), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(new_n203), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT70), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT68), .A2(G134), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT68), .A2(G134), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n203), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n204), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT70), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G131), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n208), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g030(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n205), .A2(new_n203), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n203), .A2(KEYINPUT11), .A3(G134), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n205), .B2(new_n203), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n207), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n202), .A2(new_n216), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n225));
  OAI211_X1 g039(.A(KEYINPUT0), .B(G128), .C1(new_n197), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n189), .A2(new_n191), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(KEYINPUT66), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  OR3_X1    g044(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n220), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n209), .A2(new_n210), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G137), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n217), .A2(new_n218), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n211), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT69), .A2(G131), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n237), .B2(new_n239), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n234), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n224), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT2), .B(G113), .Z(new_n245));
  XNOR2_X1  g059(.A(G116), .B(G119), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n187), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n247), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n224), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n247), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n202), .A2(new_n216), .A3(new_n223), .A4(KEYINPUT72), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n243), .A4(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n248), .B(new_n249), .C1(new_n254), .C2(new_n187), .ZN(new_n255));
  NOR2_X1   g069(.A1(G237), .A2(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G210), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n257), .B(KEYINPUT27), .Z(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n258), .B(new_n259), .Z(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  OR2_X1    g075(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n251), .A2(KEYINPUT30), .A3(new_n243), .A4(new_n253), .ZN(new_n264));
  XOR2_X1   g078(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n265));
  NAND2_X1  g079(.A1(new_n244), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n247), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n254), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n261), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n262), .A2(new_n263), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT75), .ZN(new_n271));
  INV_X1    g085(.A(new_n248), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n251), .A2(new_n243), .A3(new_n253), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n247), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n254), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n275), .B2(KEYINPUT28), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n261), .A2(new_n263), .ZN(new_n277));
  AOI21_X1  g091(.A(G902), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n262), .A2(new_n269), .A3(new_n279), .A4(new_n263), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n271), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G472), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n255), .A2(new_n261), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n267), .A2(new_n260), .A3(new_n254), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT31), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n255), .A2(KEYINPUT74), .A3(new_n261), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n267), .A2(new_n291), .A3(new_n260), .A4(new_n254), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(KEYINPUT73), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(G472), .A2(G902), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n283), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n292), .B(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n283), .B(new_n295), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n282), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G217), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(G234), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT22), .B(G137), .ZN(new_n307));
  INV_X1    g121(.A(G953), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n308), .A2(G221), .A3(G234), .ZN(new_n309));
  XOR2_X1   g123(.A(new_n307), .B(new_n309), .Z(new_n310));
  INV_X1    g124(.A(G128), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G119), .ZN(new_n312));
  INV_X1    g126(.A(G119), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G128), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT24), .B(G110), .ZN(new_n316));
  OR3_X1    g130(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT76), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT76), .B1(new_n315), .B2(new_n316), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n312), .A2(KEYINPUT77), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n313), .B2(G128), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n320), .A2(KEYINPUT77), .ZN(new_n322));
  OAI22_X1  g136(.A1(new_n319), .A2(new_n321), .B1(new_n322), .B2(new_n312), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n317), .A2(new_n318), .B1(G110), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G140), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n328), .A3(KEYINPUT16), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n327), .A2(KEYINPUT16), .A3(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G146), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(G146), .B1(new_n329), .B2(new_n330), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT78), .A4(G146), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n324), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n315), .A2(new_n316), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n323), .B2(G110), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n326), .A2(new_n328), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n188), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n331), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(KEYINPUT79), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n338), .B2(new_n343), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n310), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n310), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n344), .B2(KEYINPUT79), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n304), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n348), .A2(KEYINPUT25), .A3(new_n304), .A4(new_n350), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n306), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n348), .A2(new_n350), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n356), .A2(G902), .A3(new_n305), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(G210), .B1(G237), .B2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G107), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(G104), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n363));
  INV_X1    g177(.A(G104), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(G107), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n362), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(G104), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(KEYINPUT3), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n367), .B(KEYINPUT3), .C1(new_n364), .C2(G107), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n366), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(G101), .ZN(new_n374));
  INV_X1    g188(.A(G101), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n366), .B(new_n375), .C1(new_n369), .C2(new_n371), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT4), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n364), .A2(G107), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n378), .B1(new_n368), .B2(KEYINPUT3), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT81), .B1(new_n365), .B2(new_n363), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(new_n370), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n375), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n247), .B(new_n374), .C1(new_n377), .C2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n375), .B1(new_n368), .B2(new_n378), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(new_n381), .B2(new_n375), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n313), .A2(G116), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(KEYINPUT5), .ZN(new_n387));
  INV_X1    g201(.A(G113), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G116), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G119), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n386), .A2(new_n391), .A3(KEYINPUT5), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n389), .A2(new_n392), .B1(new_n246), .B2(new_n245), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n385), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n383), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G110), .B(G122), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n383), .A2(new_n396), .A3(new_n394), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT6), .A4(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(G125), .B1(new_n199), .B2(new_n201), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n327), .B1(new_n230), .B2(new_n233), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G224), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(G953), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n404), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n399), .A2(KEYINPUT6), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n395), .A2(new_n397), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n401), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT7), .B1(new_n405), .B2(G953), .ZN(new_n412));
  XOR2_X1   g226(.A(new_n396), .B(KEYINPUT8), .Z(new_n413));
  NAND2_X1  g227(.A1(new_n245), .A2(new_n246), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n392), .A2(KEYINPUT84), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n389), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n392), .A2(KEYINPUT84), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n413), .B1(new_n418), .B2(new_n385), .ZN(new_n419));
  INV_X1    g233(.A(new_n384), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n376), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n393), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n404), .A2(new_n412), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT85), .B1(new_n404), .B2(new_n412), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n425));
  INV_X1    g239(.A(new_n412), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n425), .B(new_n426), .C1(new_n402), .C2(new_n403), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n423), .A2(new_n424), .A3(new_n400), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n304), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n360), .B1(new_n411), .B2(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n410), .A2(new_n304), .A3(new_n359), .A4(new_n428), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(KEYINPUT86), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(KEYINPUT86), .ZN(new_n433));
  INV_X1    g247(.A(new_n429), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n359), .B1(new_n434), .B2(new_n410), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G214), .B1(G237), .B2(G902), .ZN(new_n437));
  NAND2_X1  g251(.A1(G234), .A2(G237), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(G952), .A3(new_n308), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(G902), .A3(G953), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(G898), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n432), .A2(new_n436), .A3(new_n437), .A4(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n341), .B(new_n188), .ZN(new_n447));
  INV_X1    g261(.A(G237), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n308), .A3(G214), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n190), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n256), .A2(G143), .A3(G214), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT18), .A3(G131), .ZN(new_n453));
  NAND2_X1  g267(.A1(KEYINPUT18), .A2(G131), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n447), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G113), .B(G122), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT88), .B(G104), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n457), .B(new_n458), .Z(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  AND4_X1   g274(.A1(G143), .A2(new_n448), .A3(new_n308), .A4(G214), .ZN(new_n461));
  AOI21_X1  g275(.A(G143), .B1(new_n256), .B2(G214), .ZN(new_n462));
  OAI211_X1 g276(.A(KEYINPUT17), .B(G131), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT89), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT89), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n452), .A2(new_n465), .A3(KEYINPUT17), .A4(G131), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n329), .A2(G146), .A3(new_n330), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n334), .B1(new_n468), .B2(KEYINPUT78), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n467), .A2(KEYINPUT90), .A3(new_n333), .A4(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n452), .B(new_n207), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n337), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT90), .B1(new_n475), .B2(new_n467), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n456), .B(new_n460), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n464), .A2(new_n466), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n480), .B1(new_n481), .B2(new_n337), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n473), .A3(new_n470), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n483), .A2(KEYINPUT91), .A3(new_n456), .A4(new_n460), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n456), .B1(new_n474), .B2(new_n476), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT92), .B1(new_n486), .B2(new_n459), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(KEYINPUT92), .A3(new_n459), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n304), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G475), .ZN(new_n492));
  NAND2_X1  g306(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n341), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g308(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n495));
  OAI21_X1  g309(.A(new_n494), .B1(new_n341), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n331), .B1(new_n496), .B2(G146), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n497), .A2(new_n471), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n460), .B1(new_n498), .B2(new_n456), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n485), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n502));
  NOR2_X1   g316(.A1(G475), .A2(G902), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n499), .B1(new_n479), .B2(new_n484), .ZN(new_n505));
  INV_X1    g319(.A(new_n503), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT20), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(G478), .B1(KEYINPUT93), .B2(KEYINPUT15), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XOR2_X1   g326(.A(G116), .B(G122), .Z(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G107), .ZN(new_n514));
  XNOR2_X1  g328(.A(G116), .B(G122), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n361), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT13), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n311), .B2(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n311), .A2(G143), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n190), .A2(G128), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(new_n518), .ZN(new_n523));
  OAI21_X1  g337(.A(G134), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n236), .A2(new_n522), .A3(new_n520), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n517), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n520), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n205), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n390), .A2(KEYINPUT14), .A3(G122), .ZN(new_n530));
  OAI211_X1 g344(.A(G107), .B(new_n530), .C1(new_n513), .C2(KEYINPUT14), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n531), .A3(new_n516), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT9), .B(G234), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n533), .A2(new_n303), .A3(G953), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n526), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n526), .B2(new_n532), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n537), .A2(new_n304), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT94), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n539), .A3(new_n304), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n512), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n511), .A3(new_n510), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n492), .A2(new_n508), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G469), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n201), .B(new_n193), .C1(G128), .C2(new_n197), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n385), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n202), .B2(new_n385), .ZN(new_n551));
  INV_X1    g365(.A(new_n242), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n222), .A2(new_n240), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n551), .A2(KEYINPUT12), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT12), .B1(new_n551), .B2(new_n554), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n308), .A2(G227), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT80), .ZN(new_n559));
  XNOR2_X1  g373(.A(G110), .B(G140), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT82), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n552), .B2(new_n553), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT82), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT10), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n550), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n234), .B(new_n374), .C1(new_n377), .C2(new_n382), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n202), .A2(KEYINPUT10), .A3(new_n385), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n561), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n557), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n565), .A2(new_n569), .A3(new_n568), .A4(new_n570), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n554), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n561), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n548), .B(new_n304), .C1(new_n573), .C2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n548), .A2(new_n304), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n561), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n566), .A2(new_n571), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(new_n557), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n574), .A2(new_n575), .A3(new_n561), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(G469), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n577), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G221), .B1(new_n533), .B2(G902), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n446), .A2(new_n547), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n302), .A2(new_n358), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  OAI21_X1  g404(.A(new_n304), .B1(new_n298), .B2(new_n299), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT95), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n591), .A2(new_n595), .A3(G472), .ZN(new_n596));
  INV_X1    g410(.A(new_n358), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n587), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n593), .A2(new_n594), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT33), .B1(new_n536), .B2(KEYINPUT97), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n537), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G478), .ZN(new_n602));
  INV_X1    g416(.A(G478), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n304), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n538), .B2(new_n603), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n492), .B2(new_n508), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n434), .A2(KEYINPUT96), .A3(new_n359), .A4(new_n410), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n437), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n435), .A2(KEYINPUT96), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n431), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n607), .A2(new_n611), .A3(KEYINPUT98), .A4(new_n445), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n502), .B1(new_n501), .B2(new_n503), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n505), .A2(KEYINPUT20), .A3(new_n506), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT92), .ZN(new_n616));
  AOI211_X1 g430(.A(new_n616), .B(new_n460), .C1(new_n483), .C2(new_n456), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n487), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n618), .B2(new_n485), .ZN(new_n619));
  INV_X1    g433(.A(G475), .ZN(new_n620));
  OAI22_X1  g434(.A1(new_n614), .A2(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n606), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n608), .A2(new_n437), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n430), .A2(new_n625), .A3(new_n431), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(new_n626), .A3(new_n445), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n613), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n599), .B1(new_n612), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT34), .B(G104), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  AOI22_X1  g445(.A1(new_n592), .A2(KEYINPUT95), .B1(new_n295), .B2(new_n294), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n621), .A2(new_n546), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(new_n596), .A3(new_n598), .A4(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n627), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT35), .B(G107), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  AND2_X1   g451(.A1(new_n585), .A2(new_n586), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n349), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n344), .B(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n640), .A2(new_n304), .A3(new_n306), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n353), .A2(new_n354), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n641), .B1(new_n642), .B2(new_n305), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n645), .A2(new_n547), .A3(new_n446), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(new_n596), .A3(new_n632), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n440), .B1(new_n442), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AND4_X1   g467(.A1(new_n492), .A2(new_n508), .A3(new_n545), .A4(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n650), .B1(new_n654), .B2(new_n611), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n492), .A2(new_n508), .A3(new_n545), .A4(new_n653), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n624), .A2(new_n626), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT99), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n594), .A2(KEYINPUT32), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n300), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n645), .B1(new_n661), .B2(new_n282), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XOR2_X1   g478(.A(new_n652), .B(KEYINPUT39), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n638), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT101), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT40), .Z(new_n668));
  NAND2_X1  g482(.A1(new_n275), .A2(new_n261), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n669), .A2(new_n287), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n670), .B2(G902), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n661), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n432), .A2(new_n436), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n621), .A2(new_n545), .ZN(new_n676));
  INV_X1    g490(.A(new_n437), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n676), .A2(new_n677), .A3(new_n644), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n668), .A2(new_n672), .A3(new_n675), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  NAND3_X1  g494(.A1(new_n607), .A2(new_n611), .A3(new_n653), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n302), .A2(new_n682), .A3(new_n638), .A4(new_n644), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT102), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n662), .A2(new_n685), .A3(new_n682), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  NAND2_X1  g502(.A1(new_n628), .A2(new_n612), .ZN(new_n689));
  INV_X1    g503(.A(new_n576), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n574), .B(new_n561), .C1(new_n555), .C2(new_n556), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n548), .B1(new_n692), .B2(new_n304), .ZN(new_n693));
  INV_X1    g507(.A(new_n577), .ZN(new_n694));
  INV_X1    g508(.A(new_n586), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n689), .A2(new_n302), .A3(new_n358), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NOR3_X1   g513(.A1(new_n627), .A2(new_n621), .A3(new_n546), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n302), .A2(new_n358), .A3(new_n696), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  NAND2_X1  g516(.A1(new_n696), .A2(new_n611), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n547), .A2(new_n444), .A3(new_n643), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n302), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  OAI21_X1  g521(.A(new_n288), .B1(new_n276), .B2(new_n260), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n295), .B1(new_n298), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(G902), .B1(new_n290), .B2(new_n293), .ZN(new_n710));
  INV_X1    g524(.A(G472), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n358), .B(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n696), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n444), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n546), .B1(new_n492), .B2(new_n508), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n611), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n717), .B1(new_n716), .B2(new_n611), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n713), .B(new_n715), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NAND4_X1  g536(.A1(new_n607), .A2(new_n696), .A3(new_n611), .A4(new_n653), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n644), .B(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n327), .ZN(G27));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n660), .A2(new_n300), .B1(G472), .B2(new_n281), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n727), .B1(new_n728), .B2(new_n597), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n302), .A2(KEYINPUT105), .A3(new_n358), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n587), .A2(KEYINPUT104), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n677), .B1(new_n432), .B2(new_n436), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n585), .A2(new_n733), .A3(new_n586), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n607), .A2(new_n653), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n729), .A2(new_n730), .A3(new_n738), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n740));
  INV_X1    g554(.A(new_n736), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n302), .A2(new_n740), .A3(new_n358), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n737), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NAND4_X1  g559(.A1(new_n302), .A2(new_n740), .A3(new_n358), .A4(new_n654), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  INV_X1    g561(.A(new_n621), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n622), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT43), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n643), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n632), .A2(new_n596), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT44), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n732), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n582), .A2(new_n583), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(KEYINPUT45), .ZN(new_n756));
  OAI21_X1  g570(.A(G469), .B1(new_n755), .B2(KEYINPUT45), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n578), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n577), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n586), .A3(new_n665), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n753), .A2(new_n754), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n751), .A2(KEYINPUT44), .A3(new_n752), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  NAND2_X1  g581(.A1(new_n762), .A2(new_n586), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT47), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n728), .A2(new_n597), .A3(new_n741), .A4(new_n732), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n325), .ZN(G42));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n773));
  AND4_X1   g587(.A1(new_n697), .A2(new_n701), .A3(new_n706), .A4(new_n721), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n645), .A2(new_n547), .A3(new_n652), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n302), .A3(new_n732), .ZN(new_n776));
  INV_X1    g590(.A(new_n724), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n740), .A3(new_n741), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n746), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n774), .A2(new_n744), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n623), .A2(new_n446), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n632), .A2(new_n596), .A3(new_n598), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT106), .B1(new_n783), .B2(new_n589), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n647), .B1(new_n634), .B2(new_n446), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n783), .A2(new_n589), .A3(KEYINPUT106), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n781), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n725), .B1(new_n659), .B2(new_n662), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT107), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n643), .B2(new_n653), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n355), .A2(KEYINPUT107), .A3(new_n641), .A4(new_n652), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n638), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(KEYINPUT108), .B(new_n638), .C1(new_n793), .C2(new_n794), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n720), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n718), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n801), .A3(new_n672), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n685), .B1(new_n662), .B2(new_n682), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n728), .A2(new_n681), .A3(KEYINPUT102), .A4(new_n645), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n791), .B(new_n802), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n807), .B1(KEYINPUT109), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n805), .A2(new_n810), .A3(new_n806), .ZN(new_n811));
  OAI211_X1 g625(.A(KEYINPUT53), .B(new_n790), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n687), .A2(KEYINPUT52), .A3(new_n791), .A4(new_n802), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n808), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n790), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n813), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI211_X1 g632(.A(KEYINPUT110), .B(KEYINPUT53), .C1(new_n790), .C2(new_n815), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n773), .B(new_n812), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n790), .B1(new_n809), .B2(new_n811), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n817), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n779), .B1(new_n739), .B2(new_n743), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n784), .A2(new_n786), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n825), .A3(new_n788), .A4(new_n774), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n814), .B2(new_n808), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT53), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n773), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n821), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n729), .A2(new_n730), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n754), .A2(new_n714), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n750), .A2(new_n439), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT48), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n834), .B2(KEYINPUT48), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n832), .A2(new_n358), .A3(new_n440), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n672), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n607), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n308), .A2(G952), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n750), .A2(new_n439), .A3(new_n712), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n842), .B2(new_n704), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n837), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n836), .A2(new_n834), .A3(KEYINPUT48), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n693), .A2(new_n694), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n769), .B1(new_n586), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n842), .A2(new_n732), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n675), .A2(new_n714), .A3(new_n437), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n842), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g665(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n852));
  AOI22_X1  g666(.A1(new_n848), .A2(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OR3_X1    g667(.A1(new_n851), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n839), .A2(new_n748), .A3(new_n606), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n833), .A2(new_n777), .A3(new_n832), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT51), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n830), .A2(new_n846), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(G952), .B2(G953), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n847), .B(KEYINPUT49), .Z(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n358), .A3(new_n437), .A4(new_n586), .ZN(new_n862));
  OR4_X1    g676(.A1(new_n672), .A2(new_n862), .A3(new_n675), .A4(new_n749), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n860), .A2(new_n863), .ZN(G75));
  OAI21_X1  g678(.A(KEYINPUT110), .B1(new_n827), .B2(KEYINPUT53), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n816), .A2(new_n813), .A3(new_n817), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n304), .B1(new_n867), .B2(new_n812), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT56), .B1(new_n868), .B2(G210), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n401), .A2(new_n409), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(new_n407), .Z(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT55), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n308), .A2(G952), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n869), .B2(new_n873), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n874), .A2(new_n877), .ZN(G51));
  AOI21_X1  g692(.A(new_n773), .B1(new_n867), .B2(new_n812), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n821), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n578), .B(KEYINPUT113), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT57), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n692), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n812), .B1(new_n818), .B2(new_n819), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(G902), .A3(new_n758), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT114), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n875), .B1(new_n883), .B2(new_n886), .ZN(G54));
  NAND3_X1  g701(.A1(new_n868), .A2(KEYINPUT58), .A3(G475), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n888), .A2(new_n505), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n505), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n889), .A2(new_n890), .A3(new_n875), .ZN(G60));
  XOR2_X1   g705(.A(KEYINPUT115), .B(KEYINPUT59), .Z(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n604), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n601), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(new_n879), .B2(new_n821), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n897), .A3(new_n876), .ZN(new_n898));
  INV_X1    g712(.A(new_n895), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n820), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT116), .B1(new_n901), .B2(new_n875), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n601), .B1(new_n830), .B2(new_n894), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n898), .A2(new_n902), .A3(new_n903), .ZN(G63));
  XNOR2_X1  g718(.A(KEYINPUT117), .B(KEYINPUT60), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n303), .A2(new_n304), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n884), .A2(new_n640), .A3(new_n907), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n884), .A2(new_n907), .ZN(new_n909));
  INV_X1    g723(.A(new_n356), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n876), .B(new_n908), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT61), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n911), .B(new_n913), .ZN(G66));
  INV_X1    g728(.A(new_n443), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n308), .B1(new_n915), .B2(G224), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n825), .A2(new_n788), .A3(new_n774), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(new_n308), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n870), .B1(G898), .B2(new_n308), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT119), .Z(new_n920));
  XNOR2_X1  g734(.A(new_n918), .B(new_n920), .ZN(G69));
  NAND2_X1  g735(.A1(new_n651), .A2(G953), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT124), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n746), .B1(new_n769), .B2(new_n770), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n763), .B1(new_n718), .B2(new_n800), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n831), .B2(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n687), .A2(new_n791), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n927), .A2(new_n744), .A3(new_n766), .A4(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n924), .B1(new_n929), .B2(new_n308), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n264), .A2(new_n266), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n496), .B(KEYINPUT120), .Z(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n931), .A2(new_n932), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n308), .B1(G227), .B2(G900), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT125), .B1(new_n930), .B2(new_n935), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n679), .A2(new_n928), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n940), .A2(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(KEYINPUT62), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n633), .A2(new_n607), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n943), .A2(KEYINPUT121), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n667), .A2(new_n944), .A3(new_n754), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(KEYINPUT121), .B2(new_n943), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n946), .A2(new_n728), .A3(new_n597), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n771), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n941), .A2(new_n766), .A3(new_n942), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n936), .B1(new_n949), .B2(new_n308), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n937), .B(new_n938), .C1(new_n939), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n931), .A2(new_n936), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n950), .A2(KEYINPUT122), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n950), .A2(KEYINPUT122), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n938), .B(KEYINPUT123), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n951), .A2(new_n956), .ZN(G72));
  XNOR2_X1  g771(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n711), .A2(new_n304), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n958), .B(new_n959), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n949), .B2(new_n917), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n268), .B(KEYINPUT127), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n260), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n961), .B1(new_n929), .B2(new_n917), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n260), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(new_n967), .A3(new_n876), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n823), .A2(new_n828), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n960), .B1(new_n269), .B2(new_n287), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(G57));
endmodule


