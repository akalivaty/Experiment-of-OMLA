//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT30), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n190), .A2(G137), .ZN(new_n193));
  OAI21_X1  g007(.A(G131), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n190), .B2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  INV_X1    g012(.A(G131), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .A4(new_n191), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(G128), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G143), .B(G146), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n214));
  OAI22_X1  g028(.A1(G128), .A2(new_n213), .B1(new_n214), .B2(new_n205), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n215), .B2(KEYINPUT66), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n204), .A2(G146), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n202), .A2(G143), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n201), .B1(new_n216), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n196), .A2(new_n191), .A3(new_n198), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G131), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n228), .A2(new_n200), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n203), .A2(new_n205), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n213), .B2(new_n231), .ZN(new_n237));
  AND4_X1   g051(.A1(new_n236), .A2(new_n231), .A3(new_n203), .A4(new_n205), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n229), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n189), .B1(new_n226), .B2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(G116), .A2(G119), .ZN(new_n242));
  NOR2_X1   g056(.A1(G116), .A2(G119), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  INV_X1    g062(.A(G119), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(G116), .A2(G119), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT2), .A2(G113), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT2), .A2(G113), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n247), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n205), .B1(new_n208), .B2(new_n210), .ZN(new_n258));
  AOI21_X1  g072(.A(G128), .B1(new_n203), .B2(new_n205), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT66), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n213), .A2(new_n214), .A3(G128), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n225), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n201), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT64), .B1(new_n234), .B2(new_n230), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n213), .A2(new_n236), .A3(new_n231), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n265), .A2(new_n266), .B1(new_n234), .B2(new_n233), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n228), .A2(new_n200), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n264), .A2(KEYINPUT30), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n241), .A2(new_n257), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(G237), .A2(G953), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G210), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT26), .ZN(new_n276));
  INV_X1    g090(.A(G101), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n257), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n247), .A2(new_n256), .A3(KEYINPUT68), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n264), .A2(new_n269), .A3(new_n282), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT69), .B(KEYINPUT31), .Z(new_n284));
  NAND4_X1  g098(.A1(new_n271), .A2(new_n278), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT70), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n271), .A2(new_n283), .A3(new_n278), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT31), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n264), .A2(new_n269), .A3(new_n282), .ZN(new_n289));
  INV_X1    g103(.A(new_n257), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n264), .B2(new_n269), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT28), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT71), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n283), .A2(new_n296), .A3(new_n293), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n292), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n288), .B1(new_n298), .B2(new_n278), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n188), .B1(new_n286), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n292), .A2(new_n295), .A3(new_n297), .ZN(new_n303));
  INV_X1    g117(.A(new_n278), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n303), .A2(new_n304), .B1(new_n287), .B2(KEYINPUT31), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n285), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n285), .A2(new_n306), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT32), .A3(new_n188), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G472), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n295), .A2(KEYINPUT29), .A3(new_n297), .ZN(new_n313));
  INV_X1    g127(.A(new_n282), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n226), .B2(new_n240), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(new_n283), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n264), .A2(new_n282), .A3(KEYINPUT72), .A4(new_n269), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(KEYINPUT28), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n317), .A2(KEYINPUT73), .A3(KEYINPUT28), .A4(new_n318), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n313), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n298), .A2(KEYINPUT29), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n278), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n271), .A2(new_n283), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n326), .A2(KEYINPUT29), .A3(new_n278), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n327), .A2(G902), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n312), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n187), .B1(new_n311), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n188), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n285), .B(new_n306), .ZN(new_n333));
  AOI211_X1 g147(.A(new_n301), .B(new_n332), .C1(new_n333), .C2(new_n305), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT32), .B1(new_n309), .B2(new_n188), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n325), .A2(new_n329), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G472), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(KEYINPUT74), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G217), .ZN(new_n341));
  INV_X1    g155(.A(G902), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(G234), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n345));
  INV_X1    g159(.A(G953), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(G221), .A3(G234), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT22), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(G137), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT23), .B1(new_n217), .B2(G119), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n217), .A2(G119), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(KEYINPUT75), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT75), .B1(new_n249), .B2(G128), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n249), .A2(G128), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(KEYINPUT23), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G110), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT16), .ZN(new_n360));
  INV_X1    g174(.A(G140), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(G125), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(G125), .ZN(new_n363));
  INV_X1    g177(.A(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G140), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n362), .B1(new_n366), .B2(new_n360), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n202), .ZN(new_n368));
  OAI211_X1 g182(.A(G146), .B(new_n362), .C1(new_n366), .C2(new_n360), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n249), .A2(G128), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n352), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT24), .B(G110), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n359), .A2(new_n370), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G125), .B(G140), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n202), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n353), .A2(new_n356), .A3(new_n358), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n379), .A2(KEYINPUT76), .B1(new_n372), .B2(new_n373), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n357), .A2(new_n381), .A3(new_n358), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n378), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n350), .B1(new_n375), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n383), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n359), .A2(new_n370), .A3(new_n374), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n349), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n345), .B1(new_n388), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n345), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n384), .A2(new_n387), .A3(new_n342), .A4(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n344), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n344), .A2(new_n342), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT78), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n384), .A2(new_n387), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G214), .B1(G237), .B2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G210), .B1(G237), .B2(G902), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n239), .A2(G125), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n262), .B2(G125), .ZN(new_n402));
  INV_X1    g216(.A(G224), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G953), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n402), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G104), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT3), .B1(new_n407), .B2(G107), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT3), .ZN(new_n409));
  INV_X1    g223(.A(G107), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(G104), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(G107), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n408), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n413), .A2(G101), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n411), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n277), .A2(KEYINPUT79), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT79), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G101), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n418), .A3(new_n412), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT4), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT80), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n413), .A2(G101), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT80), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT79), .B(G101), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n424), .A2(new_n408), .A3(new_n411), .A4(new_n412), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n422), .A2(new_n423), .A3(new_n425), .A4(KEYINPUT4), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n413), .A2(new_n428), .A3(G101), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n257), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT5), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n249), .A3(G116), .ZN(new_n434));
  OAI211_X1 g248(.A(G113), .B(new_n434), .C1(new_n244), .C2(new_n433), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n245), .B2(new_n244), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n410), .A2(G104), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n412), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G101), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n425), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G122), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT6), .A4(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n430), .B1(new_n421), .B2(new_n426), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n444), .B(new_n446), .C1(new_n448), .C2(new_n441), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n443), .B2(new_n446), .ZN(new_n454));
  NOR4_X1   g268(.A1(new_n448), .A2(new_n453), .A3(new_n446), .A4(new_n441), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n443), .A2(new_n446), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n406), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n448), .A2(new_n441), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT83), .B1(new_n460), .B2(new_n445), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(new_n455), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n405), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n464), .B2(new_n405), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n402), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n402), .A2(new_n404), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n445), .B(KEYINPUT8), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n436), .A2(new_n440), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n441), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n402), .A2(new_n463), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n467), .A2(new_n468), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n342), .B1(new_n462), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n400), .B1(new_n459), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n406), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n460), .A2(new_n445), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n461), .A2(new_n477), .A3(new_n455), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n447), .A2(new_n451), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n454), .A2(new_n456), .ZN(new_n481));
  INV_X1    g295(.A(new_n473), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n399), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n398), .B1(new_n475), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(G475), .A2(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n272), .A2(G143), .A3(G214), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(G143), .B1(new_n272), .B2(G214), .ZN(new_n490));
  OAI21_X1  g304(.A(G131), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G237), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n346), .A3(G214), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n204), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n199), .A3(new_n488), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n376), .A2(KEYINPUT19), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n376), .A2(KEYINPUT19), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n496), .B(new_n369), .C1(G146), .C2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT88), .B1(new_n376), .B2(new_n202), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n366), .A2(new_n502), .A3(G146), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n377), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n494), .A2(new_n488), .ZN(new_n508));
  NAND2_X1  g322(.A1(KEYINPUT18), .A2(G131), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n494), .A2(KEYINPUT18), .A3(G131), .A4(new_n488), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n501), .A2(new_n503), .A3(new_n505), .A4(new_n377), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n507), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n500), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G113), .B(G122), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(new_n407), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n491), .A2(new_n520), .A3(new_n495), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n508), .A2(KEYINPUT17), .A3(G131), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n368), .A4(new_n369), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(new_n514), .A3(new_n517), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n487), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n526));
  OAI21_X1  g340(.A(KEYINPUT89), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT20), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(KEYINPUT90), .A3(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n523), .A2(new_n514), .A3(new_n517), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n517), .B1(new_n500), .B2(new_n514), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n486), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n533));
  INV_X1    g347(.A(new_n526), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n528), .B(new_n486), .C1(new_n530), .C2(new_n531), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT90), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n527), .A2(new_n529), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n517), .B1(new_n523), .B2(new_n514), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n342), .B1(new_n530), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(KEYINPUT91), .B(new_n342), .C1(new_n530), .C2(new_n540), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(G475), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G952), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(G953), .ZN(new_n548));
  INV_X1    g362(.A(G234), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n548), .B1(new_n549), .B2(new_n492), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AOI211_X1 g365(.A(new_n342), .B(new_n346), .C1(G234), .C2(G237), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT21), .B(G898), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G128), .B(G143), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT13), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n217), .A2(KEYINPUT13), .A3(G143), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(new_n190), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(new_n190), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n248), .B2(G122), .ZN(new_n562));
  INV_X1    g376(.A(G122), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(KEYINPUT92), .A3(G116), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n248), .A2(G122), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n565), .A2(new_n410), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n410), .B1(new_n565), .B2(new_n566), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n559), .B(new_n560), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(KEYINPUT14), .ZN(new_n570));
  OR3_X1    g384(.A1(new_n563), .A2(KEYINPUT14), .A3(G116), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n565), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G107), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n555), .B(new_n190), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n565), .A2(new_n410), .A3(new_n566), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT9), .B(G234), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n578), .A2(new_n341), .A3(G953), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n569), .A2(new_n576), .A3(new_n579), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(KEYINPUT93), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT93), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n577), .A2(new_n584), .A3(new_n580), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n342), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G478), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(KEYINPUT15), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n588), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n546), .A2(new_n554), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n485), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G221), .B1(new_n578), .B2(G902), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n213), .B2(G128), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n212), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n596), .B1(new_n599), .B2(new_n440), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT81), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n425), .B(new_n439), .C1(new_n212), .C2(new_n598), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT81), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n603), .A3(new_n596), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n427), .A2(new_n267), .A3(new_n429), .ZN(new_n606));
  INV_X1    g420(.A(new_n440), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n262), .A2(KEYINPUT10), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n605), .A2(new_n606), .A3(new_n229), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(G110), .B(G140), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n346), .A2(G227), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n602), .A2(new_n603), .A3(new_n596), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n603), .B1(new_n602), .B2(new_n596), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n608), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n267), .A2(new_n429), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n426), .B2(new_n421), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n268), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n602), .B1(new_n262), .B2(new_n607), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n268), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT82), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT12), .B1(new_n268), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n621), .A2(new_n268), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n609), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n614), .A2(new_n620), .B1(new_n629), .B2(new_n612), .ZN(new_n630));
  OAI21_X1  g444(.A(G469), .B1(new_n630), .B2(G902), .ZN(new_n631));
  INV_X1    g445(.A(G469), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n628), .A2(new_n613), .A3(new_n609), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n613), .B1(new_n620), .B2(new_n609), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n632), .B(new_n342), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n595), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n593), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n340), .A2(new_n396), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT94), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n424), .ZN(G3));
  AOI21_X1  g455(.A(new_n399), .B1(new_n480), .B2(new_n483), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n398), .B1(new_n642), .B2(KEYINPUT96), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT96), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n475), .A2(new_n484), .A3(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n539), .A2(new_n545), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n586), .A2(new_n587), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n581), .A2(KEYINPUT33), .A3(new_n582), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT33), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n583), .A2(new_n651), .A3(new_n585), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n583), .A2(KEYINPUT97), .A3(new_n651), .A4(new_n585), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n587), .A2(G902), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n648), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n646), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n643), .A2(new_n645), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(G469), .A2(G902), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n629), .A2(new_n612), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n620), .A2(new_n613), .A3(new_n609), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(G469), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n635), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n392), .A2(new_n395), .A3(new_n554), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n665), .A2(new_n666), .A3(new_n594), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n309), .A2(new_n342), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(KEYINPUT95), .A3(G472), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT95), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n309), .B(new_n342), .C1(new_n671), .C2(new_n312), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n660), .A2(new_n668), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT34), .B(G104), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G6));
  OAI211_X1 g490(.A(new_n527), .B(new_n535), .C1(new_n534), .C2(new_n532), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n677), .A2(new_n545), .A3(new_n591), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n643), .A2(new_n645), .A3(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n673), .A2(new_n668), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT35), .B(G107), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G9));
  NAND2_X1  g496(.A1(new_n385), .A2(new_n386), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n350), .A2(KEYINPUT36), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n685), .A2(new_n394), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n392), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n485), .A2(new_n636), .A3(new_n592), .A4(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n673), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT37), .B(G110), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  AND2_X1   g505(.A1(new_n677), .A2(new_n591), .ZN(new_n692));
  INV_X1    g506(.A(G900), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n552), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n550), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n545), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n331), .B2(new_n339), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n643), .A2(new_n645), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n636), .A2(new_n687), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT98), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n217), .ZN(G30));
  XOR2_X1   g518(.A(new_n695), .B(KEYINPUT39), .Z(new_n705));
  OR2_X1    g519(.A1(new_n637), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT40), .Z(new_n707));
  NAND3_X1  g521(.A1(new_n304), .A2(new_n318), .A3(new_n317), .ZN(new_n708));
  AOI21_X1  g522(.A(G902), .B1(new_n708), .B2(new_n287), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n302), .B(new_n310), .C1(new_n312), .C2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT99), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n475), .A2(new_n484), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT38), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n546), .A2(new_n591), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n714), .A2(new_n687), .A3(new_n398), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n707), .A2(new_n711), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  NAND2_X1  g531(.A1(new_n654), .A2(new_n655), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n649), .A3(new_n657), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n647), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n546), .A3(new_n695), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n699), .A2(new_n700), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n340), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT100), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n340), .A2(KEYINPUT100), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G146), .ZN(G48));
  INV_X1    g542(.A(new_n554), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n635), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n609), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n425), .A2(KEYINPUT10), .A3(new_n439), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n216), .B2(new_n225), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n601), .B2(new_n604), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n229), .B1(new_n735), .B2(new_n606), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n612), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n628), .A2(new_n613), .A3(new_n609), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n632), .B1(new_n739), .B2(new_n342), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n731), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n342), .B1(new_n633), .B2(new_n634), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n742), .A2(KEYINPUT101), .A3(G469), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n729), .B(new_n594), .C1(new_n741), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n660), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n311), .A2(new_n187), .A3(new_n330), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT74), .B1(new_n336), .B2(new_n338), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n396), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT41), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G113), .ZN(G15));
  NOR2_X1   g564(.A1(new_n744), .A2(new_n679), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n396), .B(new_n751), .C1(new_n746), .C2(new_n747), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G116), .ZN(G18));
  AND2_X1   g567(.A1(new_n643), .A2(new_n645), .ZN(new_n754));
  INV_X1    g568(.A(new_n743), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n742), .A2(G469), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n730), .A3(new_n635), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n595), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n592), .A2(new_n754), .A3(new_n687), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n340), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G119), .ZN(G21));
  AOI21_X1  g575(.A(new_n312), .B1(new_n309), .B2(new_n342), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n295), .A2(new_n297), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n321), .B2(new_n322), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n288), .B1(new_n764), .B2(new_n278), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT103), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(KEYINPUT103), .B(new_n288), .C1(new_n764), .C2(new_n278), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n333), .A3(new_n768), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n188), .B(KEYINPUT102), .Z(new_n770));
  AOI21_X1  g584(.A(new_n762), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n744), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n699), .A2(new_n714), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .A4(new_n396), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G122), .ZN(G24));
  NAND2_X1  g589(.A1(new_n755), .A2(new_n757), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n594), .ZN(new_n777));
  INV_X1    g591(.A(new_n687), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n699), .A3(new_n778), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n721), .B(new_n762), .C1(new_n769), .C2(new_n770), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G125), .ZN(G27));
  INV_X1    g596(.A(new_n396), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n665), .A2(KEYINPUT104), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT104), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n635), .A2(new_n785), .A3(new_n664), .A4(new_n661), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n595), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n712), .A2(new_n398), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT42), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n721), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n332), .B1(new_n333), .B2(new_n305), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT106), .B1(new_n792), .B2(KEYINPUT32), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT106), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n300), .A2(new_n794), .A3(new_n301), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n310), .A2(KEYINPUT105), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n330), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n793), .A2(new_n797), .A3(new_n795), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n783), .B(new_n791), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n721), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n787), .A2(new_n396), .A3(new_n802), .A4(new_n788), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT42), .B1(new_n804), .B2(new_n340), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n199), .ZN(G33));
  INV_X1    g621(.A(KEYINPUT107), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n787), .A2(new_n396), .A3(new_n788), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n698), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n808), .B1(new_n698), .B2(new_n809), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n190), .ZN(G36));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n658), .A2(new_n546), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(KEYINPUT43), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT109), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(KEYINPUT43), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT110), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n673), .A2(new_n687), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n814), .B1(new_n823), .B2(KEYINPUT44), .ZN(new_n824));
  INV_X1    g638(.A(new_n788), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n823), .B2(KEYINPUT44), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n662), .A2(new_n663), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT45), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n632), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT108), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n630), .A2(KEYINPUT45), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n661), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT46), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(KEYINPUT46), .A3(new_n661), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n635), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n594), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n705), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT44), .ZN(new_n842));
  OAI211_X1 g656(.A(KEYINPUT111), .B(new_n842), .C1(new_n821), .C2(new_n822), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n824), .A2(new_n826), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(G137), .ZN(G39));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n839), .A2(KEYINPUT112), .A3(new_n594), .ZN(new_n848));
  AND2_X1   g662(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n849));
  NOR2_X1   g663(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n848), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT112), .B1(new_n839), .B2(new_n594), .ZN(new_n853));
  OAI22_X1  g667(.A1(new_n852), .A2(new_n853), .B1(KEYINPUT113), .B2(KEYINPUT47), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n340), .A2(new_n396), .A3(new_n721), .A4(new_n825), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n851), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(G140), .ZN(G42));
  AOI22_X1  g671(.A1(new_n698), .A2(new_n701), .B1(new_n779), .B2(new_n780), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n686), .B(new_n392), .C1(new_n550), .C2(new_n694), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT115), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n860), .A2(new_n787), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n711), .A3(new_n773), .ZN(new_n862));
  INV_X1    g676(.A(new_n726), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT100), .B1(new_n340), .B2(new_n722), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n858), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n727), .A2(KEYINPUT52), .A3(new_n858), .A4(new_n862), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n810), .A2(new_n811), .B1(new_n801), .B2(new_n805), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n667), .A2(new_n485), .A3(new_n672), .A4(new_n670), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT114), .B1(new_n646), .B2(new_n658), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n646), .A2(new_n591), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n720), .A2(new_n874), .A3(new_n546), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n871), .A2(new_n876), .B1(new_n673), .B2(new_n688), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n340), .B2(new_n759), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n340), .B(new_n396), .C1(new_n745), .C2(new_n751), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n639), .A3(new_n774), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n825), .A2(new_n778), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n590), .A2(new_n696), .A3(new_n589), .A4(new_n677), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n340), .A2(new_n636), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n780), .A2(new_n787), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n870), .A2(new_n880), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n869), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(KEYINPUT117), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n865), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n868), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(new_n887), .A3(KEYINPUT53), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n869), .B2(new_n887), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(KEYINPUT117), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT54), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(KEYINPUT118), .B(KEYINPUT54), .C1(new_n895), .C2(new_n897), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n758), .A2(new_n788), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n821), .A2(new_n550), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n783), .B1(new_n799), .B2(new_n800), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT48), .Z(new_n906));
  NOR4_X1   g720(.A1(new_n711), .A2(new_n902), .A3(new_n783), .A4(new_n550), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n659), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n777), .A2(new_n699), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n550), .B1(new_n818), .B2(new_n820), .ZN(new_n911));
  INV_X1    g725(.A(new_n771), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n783), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n908), .B(new_n548), .C1(new_n910), .C2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n906), .A2(new_n915), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n713), .A2(new_n777), .A3(new_n397), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n911), .A2(new_n913), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT50), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n912), .A2(new_n778), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n720), .A2(new_n546), .ZN(new_n922));
  AOI22_X1  g736(.A1(new_n903), .A2(new_n921), .B1(new_n907), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n851), .A2(new_n854), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n776), .A2(KEYINPUT119), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n776), .A2(KEYINPUT119), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n927), .A2(new_n928), .A3(new_n594), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n914), .A2(new_n825), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n924), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n916), .B1(new_n933), .B2(KEYINPUT51), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n929), .B1(new_n851), .B2(new_n854), .ZN(new_n935));
  INV_X1    g749(.A(new_n932), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT51), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n920), .A2(KEYINPUT120), .A3(new_n923), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT120), .B1(new_n920), .B2(new_n923), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n698), .A2(new_n808), .A3(new_n809), .ZN(new_n942));
  INV_X1    g756(.A(new_n697), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n340), .A2(new_n943), .A3(new_n809), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT107), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n746), .A2(new_n747), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n789), .B1(new_n946), .B2(new_n803), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n799), .A2(new_n800), .ZN(new_n948));
  INV_X1    g762(.A(new_n791), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(new_n396), .A3(new_n949), .ZN(new_n950));
  AOI22_X1  g764(.A1(new_n942), .A2(new_n945), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n877), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n760), .A2(new_n639), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n748), .A2(new_n752), .A3(new_n774), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n886), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n951), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n868), .B2(new_n892), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(KEYINPUT53), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n888), .A2(new_n889), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT54), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n900), .A2(new_n901), .A3(new_n941), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n547), .A2(new_n346), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n776), .B(KEYINPUT49), .Z(new_n967));
  NAND4_X1  g781(.A1(new_n815), .A2(new_n396), .A3(new_n397), .A4(new_n594), .ZN(new_n968));
  OR4_X1    g782(.A1(new_n711), .A2(new_n967), .A3(new_n713), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(new_n969), .ZN(G75));
  NOR2_X1   g784(.A1(new_n346), .A2(G952), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n478), .A2(new_n476), .A3(new_n479), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(new_n459), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT55), .ZN(new_n974));
  OAI211_X1 g788(.A(G210), .B(G902), .C1(new_n959), .C2(new_n960), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT56), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n976), .A3(new_n974), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT121), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n975), .A2(KEYINPUT121), .A3(new_n976), .A4(new_n974), .ZN(new_n981));
  AOI211_X1 g795(.A(new_n971), .B(new_n977), .C1(new_n980), .C2(new_n981), .ZN(G51));
  XOR2_X1   g796(.A(new_n661), .B(KEYINPUT57), .Z(new_n983));
  OR2_X1    g797(.A1(new_n958), .A2(KEYINPUT53), .ZN(new_n984));
  INV_X1    g798(.A(new_n960), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n962), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT54), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n739), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n984), .A2(new_n985), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(G902), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n991), .A2(new_n834), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n971), .B1(new_n989), .B2(new_n992), .ZN(G54));
  NAND2_X1  g807(.A1(new_n519), .A2(new_n524), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(KEYINPUT58), .A2(G475), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n971), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n991), .A2(new_n995), .A3(new_n996), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(G60));
  NAND2_X1  g815(.A1(G478), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT59), .Z(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n656), .B(new_n1004), .C1(new_n986), .C2(new_n987), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n998), .ZN(new_n1006));
  AOI22_X1  g820(.A1(KEYINPUT117), .A2(new_n896), .B1(new_n958), .B2(KEYINPUT53), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n888), .A2(new_n889), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT117), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n962), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n963), .B1(new_n1011), .B2(KEYINPUT118), .ZN(new_n1012));
  INV_X1    g826(.A(new_n901), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1004), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n656), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1006), .B1(new_n1014), .B2(new_n1015), .ZN(G63));
  NAND2_X1  g830(.A1(G217), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT122), .Z(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT60), .Z(new_n1019));
  NAND3_X1  g833(.A1(new_n990), .A2(new_n685), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1019), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n388), .B1(new_n961), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1020), .A2(new_n1022), .A3(new_n998), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT61), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1023), .B(new_n1024), .ZN(G66));
  NOR3_X1   g839(.A1(new_n553), .A2(new_n403), .A3(new_n346), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n955), .B2(new_n346), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n452), .B(new_n458), .C1(G898), .C2(new_n346), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(G69));
  NAND2_X1  g843(.A1(new_n241), .A2(new_n270), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n499), .B(KEYINPUT123), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(G900), .B2(G953), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n727), .A2(new_n858), .ZN(new_n1034));
  AND2_X1   g848(.A1(new_n844), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n841), .A2(new_n773), .A3(new_n904), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n1035), .A2(new_n856), .A3(new_n951), .A4(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1033), .B1(new_n1037), .B2(G953), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1034), .A2(new_n716), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(KEYINPUT62), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1040), .B(KEYINPUT125), .ZN(new_n1041));
  OR2_X1    g855(.A1(new_n1039), .A2(KEYINPUT62), .ZN(new_n1042));
  NOR3_X1   g856(.A1(new_n706), .A2(new_n825), .A3(new_n876), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1043), .A2(new_n340), .A3(new_n396), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n1042), .A2(new_n844), .A3(new_n856), .A4(new_n1044), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1046), .A2(G953), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1032), .B(KEYINPUT124), .Z(new_n1048));
  OAI21_X1  g862(.A(new_n1038), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n346), .B1(G227), .B2(G900), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g865(.A(new_n1050), .ZN(new_n1052));
  OAI211_X1 g866(.A(new_n1038), .B(new_n1052), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1051), .A2(new_n1053), .ZN(G72));
  NAND2_X1  g868(.A1(G472), .A2(G902), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1055), .B(KEYINPUT63), .Z(new_n1056));
  OAI21_X1  g870(.A(new_n1056), .B1(new_n1037), .B2(new_n880), .ZN(new_n1057));
  XNOR2_X1  g871(.A(new_n326), .B(KEYINPUT126), .ZN(new_n1058));
  NOR2_X1   g872(.A1(new_n1058), .A2(new_n278), .ZN(new_n1059));
  XOR2_X1   g873(.A(new_n1059), .B(KEYINPUT127), .Z(new_n1060));
  AOI21_X1  g874(.A(new_n971), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g875(.A(new_n1056), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1062), .B1(new_n1046), .B2(new_n955), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1058), .A2(new_n278), .ZN(new_n1064));
  OAI21_X1  g878(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n326), .A2(new_n304), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n1062), .B1(new_n1067), .B2(new_n287), .ZN(new_n1068));
  AOI21_X1  g882(.A(new_n1065), .B1(new_n1066), .B2(new_n1068), .ZN(G57));
endmodule


