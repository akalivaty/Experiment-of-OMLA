

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606;

  XNOR2_X1 U328 ( .A(n425), .B(n563), .ZN(n584) );
  XNOR2_X2 U329 ( .A(n424), .B(n423), .ZN(n563) );
  AND2_X1 U330 ( .A1(G226GAT), .A2(G233GAT), .ZN(n296) );
  XOR2_X1 U331 ( .A(G218GAT), .B(G92GAT), .Z(n297) );
  XNOR2_X1 U332 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U333 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U334 ( .A(n400), .B(n296), .ZN(n335) );
  XNOR2_X1 U335 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U336 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U337 ( .A(n408), .B(n407), .ZN(n411) );
  XNOR2_X1 U338 ( .A(n382), .B(n297), .ZN(n342) );
  XNOR2_X1 U339 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U340 ( .A(n443), .B(n422), .ZN(n423) );
  INV_X1 U341 ( .A(G43GAT), .ZN(n462) );
  XNOR2_X1 U342 ( .A(n345), .B(n453), .ZN(n565) );
  XNOR2_X1 U343 ( .A(n462), .B(KEYINPUT40), .ZN(n463) );
  XNOR2_X1 U344 ( .A(n464), .B(n463), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(G120GAT), .B(G71GAT), .Z(n445) );
  XOR2_X1 U346 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n299) );
  XNOR2_X1 U347 ( .A(KEYINPUT84), .B(KEYINPUT17), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n336) );
  XOR2_X1 U349 ( .A(n445), .B(n336), .Z(n301) );
  XNOR2_X1 U350 ( .A(G190GAT), .B(G99GAT), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n306) );
  XNOR2_X1 U352 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n302), .B(G127GAT), .ZN(n326) );
  XOR2_X1 U354 ( .A(n326), .B(G183GAT), .Z(n304) );
  NAND2_X1 U355 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U357 ( .A(n306), .B(n305), .Z(n314) );
  XOR2_X1 U358 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n308) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(G134GAT), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U361 ( .A(G176GAT), .B(KEYINPUT20), .Z(n310) );
  XNOR2_X1 U362 ( .A(G169GAT), .B(G15GAT), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n575) );
  XNOR2_X1 U366 ( .A(KEYINPUT37), .B(KEYINPUT100), .ZN(n428) );
  XOR2_X1 U367 ( .A(KEYINPUT88), .B(KEYINPUT1), .Z(n316) );
  XNOR2_X1 U368 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n334) );
  XOR2_X1 U370 ( .A(G148GAT), .B(G120GAT), .Z(n318) );
  XNOR2_X1 U371 ( .A(G29GAT), .B(G141GAT), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U373 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n320) );
  XNOR2_X1 U374 ( .A(G1GAT), .B(G57GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U376 ( .A(n322), .B(n321), .Z(n332) );
  XNOR2_X1 U377 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n323), .B(KEYINPUT2), .ZN(n347) );
  XOR2_X1 U379 ( .A(n347), .B(KEYINPUT4), .Z(n325) );
  NAND2_X1 U380 ( .A1(G225GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n330) );
  XOR2_X1 U382 ( .A(G134GAT), .B(KEYINPUT74), .Z(n421) );
  XOR2_X1 U383 ( .A(n421), .B(G85GAT), .Z(n328) );
  XNOR2_X1 U384 ( .A(n326), .B(G162GAT), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U388 ( .A(n334), .B(n333), .Z(n568) );
  INV_X1 U389 ( .A(n568), .ZN(n507) );
  XOR2_X1 U390 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n370) );
  XOR2_X1 U391 ( .A(G169GAT), .B(G8GAT), .Z(n438) );
  XOR2_X1 U392 ( .A(G190GAT), .B(KEYINPUT75), .Z(n400) );
  XOR2_X1 U393 ( .A(n337), .B(KEYINPUT91), .Z(n341) );
  XOR2_X1 U394 ( .A(G204GAT), .B(G211GAT), .Z(n339) );
  XNOR2_X1 U395 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n363) );
  XNOR2_X1 U397 ( .A(G36GAT), .B(n363), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n343) );
  XOR2_X1 U399 ( .A(G183GAT), .B(KEYINPUT77), .Z(n382) );
  XNOR2_X1 U400 ( .A(n438), .B(n344), .ZN(n345) );
  XNOR2_X1 U401 ( .A(G176GAT), .B(G64GAT), .ZN(n453) );
  NOR2_X1 U402 ( .A1(n575), .A2(n565), .ZN(n346) );
  XOR2_X1 U403 ( .A(KEYINPUT94), .B(n346), .Z(n368) );
  XOR2_X1 U404 ( .A(n347), .B(KEYINPUT22), .Z(n349) );
  XOR2_X1 U405 ( .A(G141GAT), .B(G22GAT), .Z(n431) );
  XNOR2_X1 U406 ( .A(G50GAT), .B(n431), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n367) );
  INV_X1 U408 ( .A(G162GAT), .ZN(n350) );
  NAND2_X1 U409 ( .A1(n350), .A2(G106GAT), .ZN(n353) );
  INV_X1 U410 ( .A(G106GAT), .ZN(n351) );
  NAND2_X1 U411 ( .A1(n351), .A2(G162GAT), .ZN(n352) );
  NAND2_X1 U412 ( .A1(n353), .A2(n352), .ZN(n355) );
  XNOR2_X1 U413 ( .A(G218GAT), .B(KEYINPUT73), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n401) );
  XOR2_X1 U415 ( .A(n401), .B(KEYINPUT23), .Z(n357) );
  NAND2_X1 U416 ( .A1(G228GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U418 ( .A(KEYINPUT24), .B(KEYINPUT85), .Z(n359) );
  XNOR2_X1 U419 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U421 ( .A(n361), .B(n360), .Z(n365) );
  XNOR2_X1 U422 ( .A(G78GAT), .B(KEYINPUT72), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n362), .B(G148GAT), .ZN(n450) );
  XNOR2_X1 U424 ( .A(n450), .B(n363), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U426 ( .A(n367), .B(n366), .Z(n571) );
  NAND2_X1 U427 ( .A1(n368), .A2(n571), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n374) );
  INV_X1 U429 ( .A(n575), .ZN(n512) );
  NOR2_X1 U430 ( .A1(n512), .A2(n571), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n371), .B(KEYINPUT26), .ZN(n591) );
  INV_X1 U432 ( .A(n591), .ZN(n372) );
  XNOR2_X1 U433 ( .A(KEYINPUT27), .B(n565), .ZN(n376) );
  NOR2_X1 U434 ( .A1(n372), .A2(n376), .ZN(n373) );
  NOR2_X1 U435 ( .A1(n374), .A2(n373), .ZN(n375) );
  NOR2_X1 U436 ( .A1(n507), .A2(n375), .ZN(n381) );
  NOR2_X1 U437 ( .A1(n568), .A2(n376), .ZN(n377) );
  XOR2_X1 U438 ( .A(KEYINPUT92), .B(n377), .Z(n536) );
  XNOR2_X1 U439 ( .A(n571), .B(KEYINPUT28), .ZN(n538) );
  INV_X1 U440 ( .A(n538), .ZN(n515) );
  NOR2_X1 U441 ( .A1(n536), .A2(n515), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n378), .B(KEYINPUT93), .ZN(n379) );
  NOR2_X1 U443 ( .A1(n512), .A2(n379), .ZN(n380) );
  NOR2_X1 U444 ( .A1(n381), .A2(n380), .ZN(n465) );
  XOR2_X1 U445 ( .A(G57GAT), .B(KEYINPUT13), .Z(n444) );
  XOR2_X1 U446 ( .A(n382), .B(n444), .Z(n384) );
  XNOR2_X1 U447 ( .A(G78GAT), .B(G211GAT), .ZN(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U449 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n386) );
  NAND2_X1 U450 ( .A1(G231GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U452 ( .A(n388), .B(n387), .Z(n390) );
  XOR2_X1 U453 ( .A(G15GAT), .B(G1GAT), .Z(n433) );
  XNOR2_X1 U454 ( .A(n433), .B(KEYINPUT14), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n390), .B(n389), .ZN(n398) );
  XOR2_X1 U456 ( .A(G155GAT), .B(G71GAT), .Z(n392) );
  XNOR2_X1 U457 ( .A(G22GAT), .B(G127GAT), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U459 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n394) );
  XNOR2_X1 U460 ( .A(G8GAT), .B(G64GAT), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U462 ( .A(n396), .B(n395), .Z(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n602) );
  INV_X1 U464 ( .A(n602), .ZN(n560) );
  INV_X1 U465 ( .A(KEYINPUT76), .ZN(n425) );
  INV_X1 U466 ( .A(n401), .ZN(n399) );
  NAND2_X1 U467 ( .A1(n399), .A2(n400), .ZN(n404) );
  INV_X1 U468 ( .A(n400), .ZN(n402) );
  NAND2_X1 U469 ( .A1(n402), .A2(n401), .ZN(n403) );
  NAND2_X1 U470 ( .A1(n404), .A2(n403), .ZN(n408) );
  NAND2_X1 U471 ( .A1(G232GAT), .A2(G233GAT), .ZN(n406) );
  INV_X1 U472 ( .A(KEYINPUT67), .ZN(n405) );
  XNOR2_X1 U473 ( .A(G99GAT), .B(G85GAT), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n409), .B(G92GAT), .ZN(n449) );
  XNOR2_X1 U475 ( .A(n449), .B(KEYINPUT9), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n412) );
  NAND2_X1 U477 ( .A1(n412), .A2(KEYINPUT11), .ZN(n416) );
  INV_X1 U478 ( .A(n412), .ZN(n414) );
  INV_X1 U479 ( .A(KEYINPUT11), .ZN(n413) );
  NAND2_X1 U480 ( .A1(n414), .A2(n413), .ZN(n415) );
  NAND2_X1 U481 ( .A1(n416), .A2(n415), .ZN(n424) );
  XNOR2_X1 U482 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n417) );
  XNOR2_X1 U483 ( .A(n417), .B(G29GAT), .ZN(n418) );
  XOR2_X1 U484 ( .A(n418), .B(KEYINPUT8), .Z(n420) );
  XNOR2_X1 U485 ( .A(G43GAT), .B(G50GAT), .ZN(n419) );
  XOR2_X1 U486 ( .A(n420), .B(n419), .Z(n443) );
  XOR2_X1 U487 ( .A(n421), .B(KEYINPUT10), .Z(n422) );
  XNOR2_X1 U488 ( .A(KEYINPUT36), .B(n584), .ZN(n520) );
  NAND2_X1 U489 ( .A1(n560), .A2(n520), .ZN(n426) );
  NOR2_X1 U490 ( .A1(n465), .A2(n426), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n506) );
  XOR2_X1 U492 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n430) );
  XNOR2_X1 U493 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n429) );
  XNOR2_X1 U494 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n437) );
  XOR2_X1 U496 ( .A(n433), .B(KEYINPUT70), .Z(n435) );
  NAND2_X1 U497 ( .A1(G229GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U498 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U500 ( .A(n439), .B(n438), .Z(n441) );
  XNOR2_X1 U501 ( .A(G197GAT), .B(G113GAT), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U503 ( .A(n443), .B(n442), .Z(n593) );
  XNOR2_X1 U504 ( .A(KEYINPUT71), .B(n593), .ZN(n576) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n458) );
  XOR2_X1 U506 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n447) );
  NAND2_X1 U507 ( .A1(G230GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U509 ( .A(n448), .B(KEYINPUT31), .Z(n452) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n456) );
  XNOR2_X1 U513 ( .A(G204GAT), .B(G106GAT), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U515 ( .A(n458), .B(n457), .ZN(n598) );
  INV_X1 U516 ( .A(n598), .ZN(n459) );
  NAND2_X1 U517 ( .A1(n576), .A2(n459), .ZN(n471) );
  NOR2_X1 U518 ( .A1(n506), .A2(n471), .ZN(n461) );
  XNOR2_X1 U519 ( .A(KEYINPUT38), .B(KEYINPUT101), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n461), .B(n460), .ZN(n488) );
  NOR2_X1 U521 ( .A1(n575), .A2(n488), .ZN(n464) );
  XOR2_X1 U522 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n473) );
  INV_X1 U523 ( .A(n465), .ZN(n470) );
  XNOR2_X1 U524 ( .A(KEYINPUT16), .B(KEYINPUT81), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n466), .B(KEYINPUT80), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n560), .A2(n584), .ZN(n467) );
  XOR2_X1 U527 ( .A(n468), .B(n467), .Z(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n495) );
  NOR2_X1 U529 ( .A1(n471), .A2(n495), .ZN(n481) );
  NAND2_X1 U530 ( .A1(n481), .A2(n507), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U532 ( .A(G1GAT), .B(n474), .Z(G1324GAT) );
  INV_X1 U533 ( .A(n565), .ZN(n509) );
  NAND2_X1 U534 ( .A1(n481), .A2(n509), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n475), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n477) );
  XNOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n512), .A2(n481), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n478), .B(KEYINPUT97), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  NAND2_X1 U542 ( .A1(n481), .A2(n515), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U544 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n484) );
  NOR2_X1 U545 ( .A1(n568), .A2(n488), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(n485), .ZN(G1328GAT) );
  NOR2_X1 U548 ( .A1(n488), .A2(n565), .ZN(n487) );
  XNOR2_X1 U549 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(G1329GAT) );
  NOR2_X1 U551 ( .A1(n488), .A2(n538), .ZN(n489) );
  XOR2_X1 U552 ( .A(KEYINPUT104), .B(n489), .Z(n490) );
  XNOR2_X1 U553 ( .A(G50GAT), .B(n490), .ZN(G1331GAT) );
  XNOR2_X1 U554 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n491), .B(KEYINPUT107), .ZN(n492) );
  XOR2_X1 U556 ( .A(KEYINPUT106), .B(n492), .Z(n497) );
  XNOR2_X1 U557 ( .A(n598), .B(KEYINPUT64), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n493), .B(KEYINPUT41), .ZN(n554) );
  INV_X1 U559 ( .A(n554), .ZN(n578) );
  NAND2_X1 U560 ( .A1(n578), .A2(n593), .ZN(n494) );
  XOR2_X1 U561 ( .A(KEYINPUT105), .B(n494), .Z(n505) );
  NOR2_X1 U562 ( .A1(n505), .A2(n495), .ZN(n501) );
  NAND2_X1 U563 ( .A1(n501), .A2(n507), .ZN(n496) );
  XNOR2_X1 U564 ( .A(n497), .B(n496), .ZN(G1332GAT) );
  NAND2_X1 U565 ( .A1(n501), .A2(n509), .ZN(n498) );
  XNOR2_X1 U566 ( .A(n498), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U567 ( .A1(n512), .A2(n501), .ZN(n499) );
  XNOR2_X1 U568 ( .A(n499), .B(KEYINPUT108), .ZN(n500) );
  XNOR2_X1 U569 ( .A(G71GAT), .B(n500), .ZN(G1334GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n503) );
  NAND2_X1 U571 ( .A1(n501), .A2(n515), .ZN(n502) );
  XNOR2_X1 U572 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U573 ( .A(G78GAT), .B(n504), .Z(G1335GAT) );
  NOR2_X1 U574 ( .A1(n506), .A2(n505), .ZN(n516) );
  NAND2_X1 U575 ( .A1(n516), .A2(n507), .ZN(n508) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(n508), .ZN(G1336GAT) );
  XNOR2_X1 U577 ( .A(G92GAT), .B(KEYINPUT110), .ZN(n511) );
  NAND2_X1 U578 ( .A1(n509), .A2(n516), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n511), .B(n510), .ZN(G1337GAT) );
  XOR2_X1 U580 ( .A(G99GAT), .B(KEYINPUT111), .Z(n514) );
  NAND2_X1 U581 ( .A1(n516), .A2(n512), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n518) );
  NAND2_X1 U584 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U586 ( .A(G106GAT), .B(n519), .Z(G1339GAT) );
  NAND2_X1 U587 ( .A1(n520), .A2(n602), .ZN(n524) );
  XOR2_X1 U588 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n522) );
  INV_X1 U589 ( .A(KEYINPUT66), .ZN(n521) );
  NOR2_X1 U590 ( .A1(n525), .A2(n598), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n526), .B(KEYINPUT115), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n527), .A2(n576), .ZN(n534) );
  XOR2_X1 U593 ( .A(KEYINPUT113), .B(KEYINPUT47), .Z(n532) );
  NOR2_X1 U594 ( .A1(n554), .A2(n593), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n528), .B(KEYINPUT46), .ZN(n529) );
  NOR2_X1 U596 ( .A1(n602), .A2(n529), .ZN(n530) );
  NAND2_X1 U597 ( .A1(n530), .A2(n563), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  NOR2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n535), .B(KEYINPUT48), .ZN(n566) );
  NOR2_X1 U601 ( .A1(n566), .A2(n536), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(KEYINPUT116), .ZN(n552) );
  NAND2_X1 U603 ( .A1(n552), .A2(n538), .ZN(n539) );
  NOR2_X1 U604 ( .A1(n575), .A2(n539), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n576), .A2(n548), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n542) );
  NAND2_X1 U608 ( .A1(n548), .A2(n578), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT117), .Z(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n546) );
  NAND2_X1 U613 ( .A1(n548), .A2(n602), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n550) );
  NAND2_X1 U617 ( .A1(n548), .A2(n584), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(n551), .ZN(G1343GAT) );
  NAND2_X1 U620 ( .A1(n591), .A2(n552), .ZN(n562) );
  NOR2_X1 U621 ( .A1(n593), .A2(n562), .ZN(n553) );
  XOR2_X1 U622 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  NOR2_X1 U623 ( .A1(n554), .A2(n562), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n556) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n555) );
  XNOR2_X1 U626 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U627 ( .A(KEYINPUT52), .B(n557), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NOR2_X1 U629 ( .A1(n560), .A2(n562), .ZN(n561) );
  XOR2_X1 U630 ( .A(G155GAT), .B(n561), .Z(G1346GAT) );
  NOR2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U632 ( .A(G162GAT), .B(n564), .Z(G1347GAT) );
  INV_X1 U633 ( .A(KEYINPUT55), .ZN(n573) );
  NOR2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT54), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT65), .ZN(n590) );
  NAND2_X1 U638 ( .A1(n571), .A2(n590), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  NOR2_X2 U640 ( .A1(n575), .A2(n574), .ZN(n585) );
  NAND2_X1 U641 ( .A1(n576), .A2(n585), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G169GAT), .B(n577), .ZN(G1348GAT) );
  NAND2_X1 U643 ( .A1(n585), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G176GAT), .ZN(G1349GAT) );
  XOR2_X1 U647 ( .A(G183GAT), .B(KEYINPUT123), .Z(n583) );
  NAND2_X1 U648 ( .A1(n585), .A2(n602), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1350GAT) );
  XNOR2_X1 U650 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n587) );
  XOR2_X1 U652 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1351GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n592), .B(KEYINPUT126), .ZN(n597) );
  NOR2_X1 U657 ( .A1(n597), .A2(n593), .ZN(n595) );
  XNOR2_X1 U658 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(G197GAT), .B(n596), .ZN(G1352GAT) );
  XOR2_X1 U661 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n600) );
  INV_X1 U662 ( .A(n597), .ZN(n604) );
  NAND2_X1 U663 ( .A1(n598), .A2(n604), .ZN(n599) );
  XNOR2_X1 U664 ( .A(n600), .B(n599), .ZN(n601) );
  XOR2_X1 U665 ( .A(G204GAT), .B(n601), .Z(G1353GAT) );
  NAND2_X1 U666 ( .A1(n604), .A2(n602), .ZN(n603) );
  XNOR2_X1 U667 ( .A(n603), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U668 ( .A1(n604), .A2(n520), .ZN(n605) );
  XNOR2_X1 U669 ( .A(n605), .B(KEYINPUT62), .ZN(n606) );
  XNOR2_X1 U670 ( .A(G218GAT), .B(n606), .ZN(G1355GAT) );
endmodule

