//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n548, new_n549, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n596, new_n597,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145, new_n1146, new_n1147;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT68), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT69), .Z(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n464), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n476), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n474), .A2(G137), .A3(new_n475), .A4(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n466), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g057(.A1(new_n472), .A2(new_n479), .A3(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n477), .A2(new_n473), .A3(new_n475), .A4(new_n467), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT71), .ZN(new_n490));
  AND4_X1   g065(.A1(G2105), .A2(new_n477), .A3(new_n473), .A4(new_n467), .ZN(new_n491));
  AOI211_X1 g066(.A(new_n486), .B(new_n490), .C1(G124), .C2(new_n491), .ZN(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n477), .A2(new_n473), .A3(new_n494), .A4(new_n467), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n465), .A2(new_n467), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n493), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n495), .A2(KEYINPUT4), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(G114), .B2(new_n475), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n477), .A2(new_n473), .A3(G2105), .A4(new_n467), .ZN(new_n502));
  INV_X1    g077(.A(G126), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n498), .A2(new_n504), .ZN(G164));
  OR2_X1    g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n512), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT72), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(G543), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n516), .A2(new_n517), .A3(new_n508), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n511), .A2(new_n520), .A3(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND4_X1  g099(.A1(new_n516), .A2(G89), .A3(new_n508), .A4(new_n517), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n516), .A2(G51), .A3(G543), .A4(new_n517), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT7), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n530), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n508), .A2(new_n527), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n525), .A2(new_n526), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(G52), .A2(new_n519), .B1(new_n521), .B2(G90), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT73), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n510), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  NAND2_X1  g115(.A1(new_n521), .A2(G81), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n519), .A2(G43), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n541), .B(new_n542), .C1(new_n510), .C2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  OR3_X1    g126(.A1(new_n518), .A2(KEYINPUT9), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT9), .B1(new_n518), .B2(new_n551), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(new_n508), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(G651), .A2(new_n558), .B1(new_n521), .B2(G91), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n554), .A2(new_n559), .ZN(G299));
  NAND4_X1  g135(.A1(new_n516), .A2(G49), .A3(G543), .A4(new_n517), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n516), .A2(G87), .A3(new_n508), .A4(new_n517), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G288));
  INV_X1    g139(.A(G61), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n506), .B2(new_n507), .ZN(new_n566));
  AND2_X1   g141(.A1(G73), .A2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n516), .A2(G48), .A3(G543), .A4(new_n517), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n516), .A2(G86), .A3(new_n508), .A4(new_n517), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G305));
  NAND2_X1  g146(.A1(new_n519), .A2(G47), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n521), .A2(G85), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n572), .B(new_n573), .C1(new_n510), .C2(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(new_n521), .A2(G92), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT10), .Z(new_n577));
  NAND2_X1  g152(.A1(G79), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G66), .ZN(new_n581));
  OAI211_X1 g156(.A(KEYINPUT75), .B(new_n580), .C1(new_n556), .C2(new_n581), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n580), .B1(new_n556), .B2(new_n581), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n583), .A2(new_n586), .B1(G54), .B2(new_n519), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n577), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(G171), .B2(new_n589), .ZN(G284));
  OAI21_X1  g166(.A(new_n590), .B1(G171), .B2(new_n589), .ZN(G321));
  NAND2_X1  g167(.A1(G299), .A2(new_n589), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n589), .B2(G168), .ZN(G297));
  OAI21_X1  g169(.A(new_n593), .B1(new_n589), .B2(G168), .ZN(G280));
  INV_X1    g170(.A(new_n588), .ZN(new_n596));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G860), .ZN(G148));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n496), .A2(new_n480), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT12), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT13), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(G2100), .ZN(new_n606));
  INV_X1    g181(.A(new_n487), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n607), .A2(G135), .ZN(new_n608));
  INV_X1    g183(.A(G123), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n475), .A2(G111), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n502), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(G2096), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(G2096), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n606), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT76), .Z(G156));
  XNOR2_X1  g193(.A(G2427), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2430), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(KEYINPUT14), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2443), .B(G2446), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2451), .B(G2454), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT77), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n626), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G1341), .B(G1348), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT78), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT79), .Z(new_n634));
  INV_X1    g209(.A(G14), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n630), .B2(new_n632), .ZN(new_n636));
  AND2_X1   g211(.A1(new_n634), .A2(new_n636), .ZN(G401));
  XOR2_X1   g212(.A(G2067), .B(G2678), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT80), .ZN(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT17), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT81), .ZN(new_n648));
  INV_X1    g223(.A(new_n645), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n648), .B1(new_n642), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2096), .B(G2100), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1971), .B(G1976), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  AND2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT20), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n657), .A2(new_n658), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n655), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n655), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1981), .B(G1986), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT83), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G20), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT23), .Z(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(G299), .B2(G16), .ZN(new_n676));
  INV_X1    g251(.A(G1956), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G35), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G162), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT29), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n678), .B1(new_n682), .B2(G2090), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT94), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n673), .A2(G5), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G301), .B2(G16), .ZN(new_n686));
  INV_X1    g261(.A(G1961), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT93), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n673), .A2(G4), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n596), .B2(new_n673), .ZN(new_n691));
  INV_X1    g266(.A(G1348), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n545), .A2(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G16), .B2(G19), .ZN(new_n695));
  INV_X1    g270(.A(G1341), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n679), .A2(G27), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G164), .B2(new_n679), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G2078), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n679), .A2(G32), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT26), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n706), .A2(new_n707), .B1(G105), .B2(new_n480), .ZN(new_n708));
  INV_X1    g283(.A(G129), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n502), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n607), .B2(G141), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n703), .B1(new_n711), .B2(new_n679), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT27), .B(G1996), .Z(new_n713));
  AOI211_X1 g288(.A(new_n697), .B(new_n702), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT90), .Z(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n687), .B2(new_n686), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n689), .A2(new_n693), .A3(new_n714), .A4(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n682), .A2(G2090), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n607), .A2(G139), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT25), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n496), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n720), .B(new_n723), .C1(new_n475), .C2(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(G29), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n679), .B2(G33), .ZN(new_n727));
  INV_X1    g302(.A(G2072), .ZN(new_n728));
  INV_X1    g303(.A(G160), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n679), .B1(new_n730), .B2(G34), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(KEYINPUT89), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(G34), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n731), .B2(KEYINPUT89), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n729), .A2(new_n679), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G2084), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n727), .A2(new_n728), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n736), .B2(new_n735), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT31), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G11), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(G11), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(G28), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n679), .B1(new_n742), .B2(G28), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n740), .B(new_n741), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n613), .B2(G29), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n746), .B1(new_n700), .B2(G2078), .C1(new_n727), .C2(new_n728), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n738), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G286), .A2(new_n673), .ZN(new_n749));
  NOR2_X1   g324(.A1(G16), .A2(G21), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n749), .A2(KEYINPUT91), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(KEYINPUT91), .B2(new_n749), .ZN(new_n752));
  INV_X1    g327(.A(G1966), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT92), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n679), .A2(G26), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G128), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n475), .A2(G116), .ZN(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n502), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n607), .B2(G140), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n758), .B1(new_n763), .B2(new_n679), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2067), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n752), .B2(new_n753), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n748), .A2(new_n755), .A3(new_n766), .ZN(new_n767));
  NOR4_X1   g342(.A1(new_n684), .A2(new_n718), .A3(new_n719), .A4(new_n767), .ZN(new_n768));
  MUX2_X1   g343(.A(G6), .B(G305), .S(G16), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT32), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1981), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n673), .A2(G22), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT85), .Z(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G166), .B2(new_n673), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1971), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n673), .A2(G23), .ZN(new_n776));
  INV_X1    g351(.A(G288), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n673), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT33), .B(G1976), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n778), .B(new_n779), .Z(new_n780));
  NOR3_X1   g355(.A1(new_n771), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  MUX2_X1   g359(.A(G24), .B(G290), .S(G16), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1986), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n679), .A2(G25), .ZN(new_n787));
  INV_X1    g362(.A(G119), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n475), .A2(G107), .ZN(new_n789));
  OAI21_X1  g364(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n790));
  OAI22_X1  g365(.A1(new_n502), .A2(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n607), .B2(G131), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n787), .B1(new_n792), .B2(new_n679), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT35), .B(G1991), .Z(new_n794));
  XOR2_X1   g369(.A(new_n793), .B(new_n794), .Z(new_n795));
  NOR2_X1   g370(.A1(new_n786), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n783), .A2(new_n784), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT87), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT86), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n768), .B1(new_n800), .B2(KEYINPUT36), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT36), .B1(new_n797), .B2(new_n799), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n798), .B2(new_n799), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n801), .A2(new_n803), .ZN(G311));
  INV_X1    g379(.A(G311), .ZN(G150));
  NAND2_X1  g380(.A1(new_n596), .A2(G559), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT38), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n521), .A2(G93), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT95), .B(G55), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n808), .B1(new_n510), .B2(new_n809), .C1(new_n518), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n545), .B(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n807), .B(new_n812), .Z(new_n813));
  INV_X1    g388(.A(KEYINPUT39), .ZN(new_n814));
  AOI21_X1  g389(.A(G860), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT96), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n811), .A2(G860), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(G145));
  XNOR2_X1  g395(.A(new_n792), .B(KEYINPUT99), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(new_n604), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n725), .A2(KEYINPUT97), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n711), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n822), .B(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n763), .B(G164), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n491), .A2(G130), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT98), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n828), .A2(new_n475), .A3(G118), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n475), .B2(G118), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n830), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n827), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G142), .B2(new_n607), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n826), .B(new_n833), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n825), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n614), .B(G160), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G162), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n835), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT100), .B(G37), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g416(.A(new_n588), .B(G299), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT41), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n599), .B(new_n812), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n844), .A2(new_n842), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n843), .A2(KEYINPUT101), .A3(new_n844), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT42), .ZN(new_n851));
  XOR2_X1   g426(.A(G303), .B(KEYINPUT102), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(G290), .ZN(new_n853));
  XNOR2_X1  g428(.A(G305), .B(G288), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n853), .B(new_n854), .Z(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n850), .A2(KEYINPUT42), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n851), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n856), .B1(new_n851), .B2(new_n857), .ZN(new_n859));
  OAI21_X1  g434(.A(G868), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n811), .A2(new_n589), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(G295));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n861), .ZN(G331));
  INV_X1    g438(.A(new_n842), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n812), .B(G301), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(G286), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(G286), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  INV_X1    g444(.A(new_n843), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n855), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n856), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n839), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n871), .B2(new_n855), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n875), .A2(KEYINPUT43), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n882));
  NAND2_X1  g457(.A1(new_n872), .A2(new_n873), .ZN(new_n883));
  OAI21_X1  g458(.A(KEYINPUT44), .B1(new_n883), .B2(new_n877), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n876), .B1(new_n880), .B2(new_n874), .ZN(new_n885));
  OAI22_X1  g460(.A1(new_n881), .A2(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G397));
  INV_X1    g461(.A(KEYINPUT126), .ZN(new_n887));
  INV_X1    g462(.A(G1384), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n498), .B2(new_n504), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT45), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n471), .A2(new_n478), .A3(G40), .A4(new_n481), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G2067), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n763), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT104), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n711), .B(G1996), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n792), .B(new_n794), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT105), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(G290), .B(G1986), .Z(new_n903));
  AOI21_X1  g478(.A(new_n894), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n905));
  AND4_X1   g480(.A1(G40), .A2(new_n471), .A3(new_n478), .A4(new_n481), .ZN(new_n906));
  INV_X1    g481(.A(G114), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n499), .B1(new_n907), .B2(G2105), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(new_n491), .B2(G126), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n496), .A2(new_n497), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G1384), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT50), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n905), .B(new_n906), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n914), .B(new_n888), .C1(new_n498), .C2(new_n504), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n892), .B1(new_n889), .B2(KEYINPUT50), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(new_n905), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n677), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT57), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n554), .B2(new_n559), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n554), .A2(new_n921), .A3(new_n559), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(KEYINPUT45), .B(new_n888), .C1(new_n498), .C2(new_n504), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n891), .A2(new_n906), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT56), .B(G2072), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n920), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n889), .A2(KEYINPUT50), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n906), .A3(new_n916), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n918), .A2(KEYINPUT111), .A3(new_n916), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n692), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n889), .A2(new_n892), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n895), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n937), .B1(new_n936), .B2(new_n939), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(new_n588), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n925), .B1(new_n920), .B2(new_n929), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n930), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT60), .B1(new_n940), .B2(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n936), .A2(new_n939), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT112), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT60), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(new_n950), .A3(new_n596), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(KEYINPUT60), .B(new_n588), .C1(new_n940), .C2(new_n941), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT61), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n918), .A2(new_n905), .B1(new_n914), .B2(new_n913), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n931), .A2(new_n906), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT108), .ZN(new_n957));
  AOI21_X1  g532(.A(G1956), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n927), .A2(new_n928), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n923), .A2(new_n924), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n954), .B1(new_n961), .B2(new_n943), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n958), .B2(new_n959), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(new_n930), .A3(KEYINPUT61), .ZN(new_n964));
  NOR2_X1   g539(.A1(KEYINPUT114), .A2(KEYINPUT59), .ZN(new_n965));
  NAND2_X1  g540(.A1(KEYINPUT114), .A2(KEYINPUT59), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT58), .B(G1341), .Z(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n889), .B2(new_n892), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(KEYINPUT113), .B(new_n968), .C1(new_n889), .C2(new_n892), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n891), .A2(new_n906), .A3(new_n926), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n971), .B(new_n972), .C1(new_n973), .C2(G1996), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n965), .B(new_n967), .C1(new_n974), .C2(new_n545), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(KEYINPUT114), .A3(KEYINPUT59), .A4(new_n545), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n953), .A2(new_n962), .A3(new_n964), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n944), .B1(new_n952), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT115), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT61), .B1(new_n963), .B2(new_n930), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n974), .A2(new_n545), .ZN(new_n983));
  INV_X1    g558(.A(new_n965), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n966), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n976), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n951), .A2(new_n953), .A3(new_n987), .A4(new_n964), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n989), .A3(new_n944), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n934), .A2(new_n687), .A3(new_n935), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n891), .A2(KEYINPUT120), .A3(new_n906), .A4(new_n926), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT53), .ZN(new_n993));
  INV_X1    g568(.A(G2078), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n891), .A2(new_n994), .A3(new_n906), .A4(new_n926), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n927), .A2(KEYINPUT53), .A3(new_n992), .A4(new_n994), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n991), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(G171), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n927), .A2(KEYINPUT53), .A3(new_n994), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n991), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G171), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT119), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n1007), .A3(G171), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1000), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(KEYINPUT121), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT121), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT107), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n892), .B1(new_n913), .B2(KEYINPUT45), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1971), .B1(new_n1015), .B2(new_n891), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT106), .B(G2090), .Z(new_n1017));
  AND3_X1   g592(.A1(new_n918), .A2(new_n916), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1014), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G303), .A2(G8), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT55), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1971), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n913), .A2(KEYINPUT45), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n906), .A2(new_n926), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n918), .A2(new_n916), .A3(new_n1017), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(KEYINPUT107), .A3(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1019), .A2(new_n1022), .A3(G8), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n913), .A2(new_n906), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n561), .A2(new_n562), .A3(G1976), .A4(new_n563), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(G288), .B2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1030), .A2(G8), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(G8), .B(new_n1031), .C1(new_n889), .C2(new_n892), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT52), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G305), .A2(G1981), .ZN(new_n1037));
  INV_X1    g612(.A(G1981), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(KEYINPUT49), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1030), .A2(new_n1040), .A3(G8), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT49), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1034), .B(new_n1036), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT109), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1042), .ZN(new_n1045));
  INV_X1    g620(.A(G8), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n938), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1047), .A3(new_n1040), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1044), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n955), .A2(new_n957), .A3(new_n1017), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1046), .B1(new_n1052), .B2(new_n1026), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1029), .B(new_n1051), .C1(new_n1022), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G286), .A2(G8), .ZN(new_n1055));
  XOR2_X1   g630(.A(new_n1055), .B(KEYINPUT116), .Z(new_n1056));
  XNOR2_X1  g631(.A(new_n1055), .B(KEYINPUT116), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT51), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n932), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1060), .A2(new_n736), .B1(new_n973), .B2(new_n753), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1056), .B(new_n1059), .C1(new_n1061), .C2(new_n1046), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n1056), .B2(KEYINPUT117), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n1061), .B2(new_n1056), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n927), .A2(G1966), .B1(G2084), .B2(new_n932), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1057), .B1(new_n1066), .B2(G8), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1062), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1054), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n995), .B(KEYINPUT53), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(G301), .A3(new_n991), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1071), .A2(KEYINPUT54), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n998), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT122), .B1(new_n998), .B2(G171), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1013), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n981), .A2(new_n990), .A3(new_n1012), .A4(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1048), .A2(new_n1032), .A3(new_n777), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1039), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1047), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1029), .B2(new_n1043), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1066), .A2(G8), .A3(G168), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT63), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1085), .A2(new_n1029), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT110), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1019), .A2(G8), .A3(new_n1028), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n1087), .B(new_n1043), .C1(new_n1088), .C2(new_n1021), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1028), .A2(G8), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT107), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1021), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1043), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT110), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1086), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1084), .B1(new_n1054), .B2(new_n1083), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1082), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1029), .A2(new_n1051), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1053), .A2(new_n1022), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1068), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1068), .A2(new_n1102), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1008), .A2(new_n1006), .B1(new_n1068), .B2(new_n1102), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1104), .B1(new_n1108), .B2(new_n1100), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1097), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n904), .B1(new_n1078), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n894), .B1(new_n897), .B2(new_n711), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT46), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n894), .A2(G1996), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1114), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(KEYINPUT124), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT47), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n763), .A2(new_n895), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n792), .A2(new_n794), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n899), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n893), .B1(new_n899), .B2(new_n901), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n894), .A2(G1986), .A3(G290), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n893), .A2(new_n1123), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1120), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n887), .B1(new_n1112), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1129), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n1132));
  AOI211_X1 g707(.A(KEYINPUT119), .B(G301), .C1(new_n1070), .C2(new_n991), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1007), .B1(new_n1004), .B2(G171), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1133), .A2(new_n1134), .A3(new_n999), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1135), .B2(new_n1010), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1136), .A2(new_n1012), .A3(new_n1075), .A4(new_n1069), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n989), .B1(new_n988), .B2(new_n944), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1110), .B1(new_n1139), .B2(new_n990), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT126), .B(new_n1131), .C1(new_n1140), .C2(new_n904), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1130), .A2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g717(.A1(G227), .A2(new_n462), .ZN(new_n1144));
  AOI21_X1  g718(.A(new_n1144), .B1(new_n634), .B2(new_n636), .ZN(new_n1145));
  AOI21_X1  g719(.A(G229), .B1(new_n1145), .B2(KEYINPUT127), .ZN(new_n1146));
  OAI211_X1 g720(.A(new_n840), .B(new_n1146), .C1(KEYINPUT127), .C2(new_n1145), .ZN(new_n1147));
  NOR2_X1   g721(.A1(new_n881), .A2(new_n1147), .ZN(G308));
  INV_X1    g722(.A(G308), .ZN(G225));
endmodule


