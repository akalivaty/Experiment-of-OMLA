//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n450, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n554, new_n555, new_n556, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1258, new_n1259;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT69), .Z(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND3_X1   g039(.A1(KEYINPUT71), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT3), .B1(KEYINPUT71), .B2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n474), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n471), .B1(new_n481), .B2(G2105), .ZN(G160));
  OAI21_X1  g057(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n483), .A2(KEYINPUT72), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(KEYINPUT72), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n484), .A2(G124), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n465), .A2(new_n466), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n489), .B1(new_n491), .B2(G136), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n486), .A2(new_n492), .ZN(G162));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n465), .B2(new_n466), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n496), .A2(KEYINPUT4), .B1(new_n477), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n498), .A2(new_n502), .ZN(G164));
  OR2_X1    g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT73), .B(G651), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(G50), .A3(G543), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n506), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n512), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(new_n516), .A2(G89), .A3(new_n506), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n515), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g102(.A(G51), .B(G543), .C1(new_n527), .C2(new_n513), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n532), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n506), .A2(new_n529), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n522), .A2(new_n528), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  OAI211_X1 g111(.A(G90), .B(new_n506), .C1(new_n527), .C2(new_n513), .ZN(new_n537));
  OAI211_X1 g112(.A(G52), .B(G543), .C1(new_n527), .C2(new_n513), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n504), .B2(new_n505), .ZN(new_n540));
  AND2_X1   g115(.A1(G77), .A2(G543), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n511), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n537), .A2(new_n538), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND3_X1  g119(.A1(new_n516), .A2(G81), .A3(new_n506), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n516), .A2(G43), .A3(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n504), .B2(new_n505), .ZN(new_n548));
  AND2_X1   g123(.A1(G68), .A2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n511), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NOR2_X1   g132(.A1(new_n527), .A2(new_n513), .ZN(new_n558));
  NAND2_X1  g133(.A1(G53), .A2(G543), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n516), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n504), .B2(new_n505), .ZN(new_n565));
  AND2_X1   g140(.A1(G78), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g142(.A(G91), .B(new_n506), .C1(new_n527), .C2(new_n513), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(G299));
  NAND3_X1  g144(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n570), .B(new_n571), .C1(new_n519), .C2(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n506), .A2(G61), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n510), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT75), .B1(new_n579), .B2(new_n510), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n516), .A2(G86), .A3(new_n506), .ZN(new_n582));
  AND2_X1   g157(.A1(G48), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(new_n527), .B2(new_n513), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n510), .ZN(new_n588));
  XNOR2_X1  g163(.A(KEYINPUT76), .B(G47), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n516), .A2(G543), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n516), .A2(G85), .A3(new_n506), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  OAI211_X1 g168(.A(G54), .B(G543), .C1(new_n527), .C2(new_n513), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n504), .B2(new_n505), .ZN(new_n596));
  AND2_X1   g171(.A1(G79), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT77), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n594), .A2(new_n601), .A3(new_n598), .ZN(new_n602));
  OAI211_X1 g177(.A(G92), .B(new_n506), .C1(new_n527), .C2(new_n513), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n516), .A2(KEYINPUT10), .A3(G92), .A4(new_n506), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n600), .A2(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n593), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n593), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n568), .A2(new_n567), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n560), .B2(new_n562), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n610), .B1(new_n612), .B2(G868), .ZN(G297));
  OAI21_X1  g188(.A(new_n610), .B1(new_n612), .B2(G868), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n607), .B1(new_n615), .B2(G860), .ZN(G148));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n607), .B2(new_n615), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n605), .A2(new_n606), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n594), .A2(new_n601), .A3(new_n598), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n601), .B1(new_n594), .B2(new_n598), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR3_X1   g197(.A1(new_n622), .A2(KEYINPUT78), .A3(G559), .ZN(new_n623));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NOR3_X1   g199(.A1(new_n618), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(new_n624), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n477), .A2(new_n469), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT13), .Z(new_n630));
  INV_X1    g205(.A(KEYINPUT79), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G2100), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(KEYINPUT79), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n484), .A2(new_n485), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G123), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  INV_X1    g213(.A(G111), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n638), .B1(new_n639), .B2(G2105), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n491), .B2(G135), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n630), .A2(new_n631), .A3(G2100), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n642), .A2(G2096), .ZN(new_n645));
  NAND4_X1  g220(.A1(new_n634), .A2(new_n643), .A3(new_n644), .A4(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT80), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n654), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n654), .A2(new_n658), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n654), .A2(new_n658), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(G14), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT81), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT18), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n668), .A2(new_n669), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n676), .B(new_n680), .Z(G227));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT20), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n684), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n684), .B2(new_n690), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT82), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n698));
  XOR2_X1   g273(.A(new_n697), .B(new_n698), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n693), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n699), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n700), .A2(new_n704), .ZN(G229));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(KEYINPUT36), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G16), .B2(G24), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n710), .A2(G1986), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(G1986), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n711), .A2(new_n712), .B1(new_n706), .B2(KEYINPUT36), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G25), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT83), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G107), .B2(new_n464), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT85), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n491), .A2(G131), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT84), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n636), .A2(new_n723), .A3(G119), .ZN(new_n724));
  INV_X1    g299(.A(G119), .ZN(new_n725));
  OAI21_X1  g300(.A(KEYINPUT84), .B1(new_n635), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n722), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n716), .B1(new_n727), .B2(new_n714), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n728), .A2(new_n730), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n713), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G22), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G166), .B2(new_n734), .ZN(new_n736));
  INV_X1    g311(.A(G1971), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n581), .A2(new_n585), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G6), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT32), .B(G1981), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  MUX2_X1   g319(.A(G23), .B(G288), .S(G16), .Z(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT33), .B(G1976), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n740), .B(new_n742), .C1(G6), .C2(G16), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n738), .A2(new_n744), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n749), .A2(new_n751), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n707), .B(new_n733), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n607), .A2(G16), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G4), .B2(G16), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(KEYINPUT88), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(KEYINPUT88), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT89), .B(G1348), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OR3_X1    g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n714), .A2(G35), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G162), .B2(new_n714), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT29), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G2090), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n714), .A2(G32), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n484), .A2(G129), .A3(new_n485), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT26), .Z(new_n771));
  OAI211_X1 g346(.A(G141), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n469), .A2(G105), .ZN(new_n773));
  AND3_X1   g348(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n768), .B1(new_n776), .B2(new_n714), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(KEYINPUT91), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT27), .B(G1996), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(KEYINPUT91), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n767), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n766), .A2(G2090), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G11), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT94), .B(G28), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT30), .ZN(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n788), .B2(KEYINPUT30), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(new_n464), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT25), .ZN(new_n794));
  NAND2_X1  g369(.A1(G103), .A2(G2104), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G2105), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n491), .A2(G139), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G33), .B(new_n799), .S(G29), .Z(new_n800));
  OAI221_X1 g375(.A(new_n791), .B1(new_n642), .B2(new_n714), .C1(new_n800), .C2(G2072), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G21), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G168), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT92), .B(G1966), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n714), .A2(G27), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G164), .B2(new_n714), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2078), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G2072), .B2(new_n800), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n734), .A2(G19), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n551), .B2(new_n734), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G1341), .Z(new_n813));
  NOR2_X1   g388(.A1(G171), .A2(new_n734), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G5), .B2(new_n734), .ZN(new_n815));
  INV_X1    g390(.A(G1961), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n806), .A2(new_n810), .A3(new_n813), .A4(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT24), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n714), .B1(new_n821), .B2(G34), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n821), .B2(G34), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G160), .B2(G29), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(G2084), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT96), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(G2084), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n803), .A2(new_n804), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n815), .A2(new_n816), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n826), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n820), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n817), .A2(new_n818), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n714), .A2(G26), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n484), .A2(G128), .A3(new_n485), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n837));
  INV_X1    g412(.A(G116), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(G2105), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n491), .B2(G140), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n835), .B1(new_n841), .B2(G29), .ZN(new_n842));
  INV_X1    g417(.A(G2067), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n734), .A2(G20), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT23), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n612), .B2(new_n734), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G1956), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n832), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n763), .A2(new_n785), .A3(new_n831), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n754), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n707), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n752), .A2(new_n753), .ZN(new_n853));
  INV_X1    g428(.A(new_n733), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT97), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n858));
  NOR4_X1   g433(.A1(new_n855), .A2(new_n754), .A3(new_n850), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n857), .A2(new_n859), .ZN(G311));
  NAND2_X1  g435(.A1(new_n851), .A2(new_n856), .ZN(G150));
  NAND2_X1  g436(.A1(new_n607), .A2(G559), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT38), .Z(new_n863));
  NAND3_X1  g438(.A1(new_n516), .A2(G93), .A3(new_n506), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n516), .A2(G55), .A3(G543), .ZN(new_n865));
  INV_X1    g440(.A(G67), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n504), .B2(new_n505), .ZN(new_n867));
  AND2_X1   g442(.A1(G80), .A2(G543), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n511), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n864), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n551), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n864), .A2(new_n865), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n863), .B(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n877), .A2(new_n878), .A3(G860), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n873), .A2(G860), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT37), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n879), .A2(new_n881), .ZN(G145));
  NAND2_X1  g457(.A1(G162), .A2(G160), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n884));
  INV_X1    g459(.A(G160), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n486), .A2(new_n492), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n883), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n884), .B1(new_n883), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n642), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n887), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n885), .A2(new_n886), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT98), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n642), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n883), .A2(new_n884), .A3(new_n887), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n775), .A2(new_n799), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n769), .A2(new_n774), .A3(new_n793), .A4(new_n798), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n484), .A2(G130), .A3(new_n485), .ZN(new_n901));
  OAI21_X1  g476(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n902));
  INV_X1    g477(.A(G118), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(G2105), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n904), .B1(new_n491), .B2(G142), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n629), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n629), .A3(new_n905), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n900), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n898), .A3(new_n899), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n477), .A2(new_n497), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n499), .A2(new_n501), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n841), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n836), .A2(G164), .A3(new_n840), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n727), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n727), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n913), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n727), .A2(new_n921), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n926), .A2(new_n922), .A3(new_n912), .A4(new_n910), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n897), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G37), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n897), .B1(new_n927), .B2(new_n925), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT99), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n925), .A2(new_n927), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n896), .A3(new_n890), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT99), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n929), .A4(new_n928), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n939));
  OR3_X1    g514(.A1(new_n618), .A2(new_n623), .A3(new_n875), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n875), .B1(new_n618), .B2(new_n623), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n607), .A2(G299), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n622), .A2(new_n612), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT41), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n607), .B2(G299), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT100), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n622), .B2(new_n612), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n607), .A2(KEYINPUT100), .A3(G299), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n940), .B(new_n941), .C1(new_n944), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n940), .A2(new_n941), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT100), .B1(new_n607), .B2(G299), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n622), .A2(new_n948), .A3(new_n612), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n943), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(G303), .B(G288), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(G305), .A2(new_n708), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n739), .A2(G290), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(G305), .B(G290), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n958), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n962), .A2(new_n964), .A3(KEYINPUT42), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT42), .B1(new_n962), .B2(new_n964), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n952), .B(new_n957), .C1(new_n967), .C2(KEYINPUT102), .ZN(new_n968));
  INV_X1    g543(.A(new_n966), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n962), .A2(new_n964), .A3(KEYINPUT42), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT102), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n957), .A2(new_n952), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n967), .A2(KEYINPUT102), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n968), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G868), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n870), .A2(G868), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n939), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  AOI211_X1 g554(.A(KEYINPUT103), .B(new_n977), .C1(new_n975), .C2(G868), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(G295));
  NAND2_X1  g556(.A1(new_n976), .A2(new_n978), .ZN(G331));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n983));
  XNOR2_X1  g558(.A(G286), .B(G301), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n875), .B(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n951), .B2(new_n944), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n875), .A2(new_n984), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n875), .A2(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT104), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT104), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n875), .A2(new_n990), .A3(new_n984), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n956), .A2(new_n987), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n962), .A2(new_n964), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n986), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n929), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n986), .A2(new_n992), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n993), .B1(new_n996), .B2(KEYINPUT105), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n986), .A2(new_n992), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n995), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n983), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n989), .A2(new_n987), .A3(new_n991), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n950), .A2(new_n949), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n946), .B1(new_n1004), .B2(new_n943), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n942), .A2(KEYINPUT41), .A3(new_n943), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n956), .A2(new_n988), .A3(new_n987), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n993), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n995), .A2(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1010), .A2(KEYINPUT107), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT43), .B1(new_n1010), .B2(KEYINPUT107), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1002), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n996), .A2(KEYINPUT105), .ZN(new_n1015));
  INV_X1    g590(.A(new_n993), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n999), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n994), .A2(new_n929), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1001), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n995), .A2(new_n1009), .A3(KEYINPUT43), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1014), .B(new_n983), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1016), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1018), .A2(new_n1024), .A3(new_n1001), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1014), .B1(new_n1026), .B2(new_n983), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1013), .B1(new_n1022), .B2(new_n1027), .ZN(G397));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(G166), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G40), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n1034), .B(new_n471), .C1(new_n481), .C2(G2105), .ZN(new_n1035));
  INV_X1    g610(.A(G1384), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n498), .B2(new_n502), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT45), .B(new_n1036), .C1(new_n498), .C2(new_n502), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n737), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n918), .A2(new_n1043), .A3(new_n1036), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1037), .A2(KEYINPUT50), .ZN(new_n1045));
  INV_X1    g620(.A(G2090), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1035), .A2(new_n1044), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT110), .B(G8), .Z(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1033), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(G8), .A3(new_n1033), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT109), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1030), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT109), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(new_n1033), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1051), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1041), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2084), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1035), .A2(new_n1044), .A3(new_n1045), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1050), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(G286), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT112), .B(G1981), .Z(new_n1065));
  NAND3_X1  g640(.A1(new_n581), .A2(new_n585), .A3(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT113), .B(G86), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n506), .B(new_n1067), .C1(new_n527), .C2(new_n513), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1068), .A2(KEYINPUT114), .A3(new_n584), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT114), .B1(new_n1068), .B2(new_n584), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n576), .ZN(new_n1071));
  INV_X1    g646(.A(G1981), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT49), .B(new_n1066), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1070), .A2(new_n576), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1069), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G1981), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(KEYINPUT115), .A3(KEYINPUT49), .A4(new_n1066), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1066), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1072), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(G1384), .B1(new_n916), .B2(new_n917), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1049), .B1(new_n1035), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1075), .A2(new_n1080), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n1088));
  INV_X1    g663(.A(G1976), .ZN(new_n1089));
  OR2_X1    g664(.A1(G288), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1088), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT111), .B(G1976), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(G288), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1087), .A2(KEYINPUT117), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT117), .B1(new_n1087), .B2(new_n1095), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1057), .B(new_n1064), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1054), .A2(new_n1033), .ZN(new_n1101));
  NOR4_X1   g676(.A1(new_n1101), .A2(new_n1063), .A3(new_n1099), .A4(G286), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(new_n1087), .A3(new_n1095), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1066), .B(KEYINPUT116), .Z(new_n1106));
  NOR2_X1   g681(.A1(G288), .A2(G1976), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n1087), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1086), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1087), .A2(new_n1095), .ZN(new_n1110));
  OAI22_X1  g685(.A1(new_n1108), .A2(new_n1109), .B1(new_n1103), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G168), .A2(new_n1049), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(KEYINPUT51), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1063), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1030), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT51), .B1(new_n1115), .B2(new_n1112), .ZN(new_n1116));
  AOI211_X1 g691(.A(G168), .B(new_n1049), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1117));
  OAI211_X1 g692(.A(KEYINPUT62), .B(new_n1114), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1035), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n816), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G2078), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1035), .A2(new_n1039), .A3(new_n1122), .A4(new_n1040), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1124), .A3(KEYINPUT53), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1121), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(G301), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1118), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1062), .A2(G286), .A3(new_n1050), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1132), .B(KEYINPUT51), .C1(new_n1112), .C2(new_n1115), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT62), .B1(new_n1133), .B2(new_n1114), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1051), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1056), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1055), .B1(new_n1054), .B2(new_n1033), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1097), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1087), .A2(KEYINPUT117), .A3(new_n1095), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1111), .B1(new_n1135), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(new_n611), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n612), .B(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT56), .B(G2072), .Z(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1035), .A2(new_n1039), .A3(new_n1040), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(G1956), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1151), .A2(KEYINPUT119), .B1(new_n1152), .B2(new_n1119), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1147), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1085), .A2(G160), .A3(G40), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1035), .A2(KEYINPUT120), .A3(new_n1085), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n843), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1119), .A2(new_n759), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n622), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1156), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1119), .A2(new_n1152), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n1154), .B2(new_n1150), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1155), .ZN(new_n1168));
  XNOR2_X1  g743(.A(G299), .B(new_n1146), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1165), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1170), .B2(new_n1156), .ZN(new_n1173));
  XNOR2_X1  g748(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(G1341), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1159), .A2(new_n1160), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(G1996), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1035), .A2(new_n1039), .A3(new_n1177), .A4(new_n1040), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n551), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT59), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1182), .A3(new_n551), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1163), .ZN(new_n1185));
  AOI21_X1  g760(.A(G2067), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1185), .A2(new_n1186), .A3(new_n607), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT60), .B1(new_n1187), .B2(new_n1164), .ZN(new_n1188));
  OR4_X1    g763(.A1(KEYINPUT60), .A2(new_n1185), .A3(new_n1186), .A4(new_n622), .ZN(new_n1189));
  AND4_X1   g764(.A1(new_n1173), .A2(new_n1184), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1169), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1151), .A2(KEYINPUT119), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1192), .A2(new_n1147), .A3(new_n1155), .A4(new_n1166), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1191), .A2(KEYINPUT61), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT122), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1194), .B(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1171), .B1(new_n1190), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1121), .A2(KEYINPUT124), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1120), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1202));
  OAI21_X1  g777(.A(G171), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(KEYINPUT125), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1205), .B(G171), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT54), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1207), .B1(new_n1129), .B2(G301), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1204), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1133), .A2(new_n1114), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1211), .A2(G301), .A3(new_n1198), .A4(new_n1200), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1212), .B1(G301), .B2(new_n1129), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1210), .B1(new_n1213), .B2(new_n1207), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1209), .A2(new_n1142), .A3(new_n1214), .ZN(new_n1215));
  OAI211_X1 g790(.A(new_n1105), .B(new_n1143), .C1(new_n1197), .C2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1035), .A2(new_n1038), .A3(new_n1037), .ZN(new_n1217));
  NAND2_X1  g792(.A1(G290), .A2(G1986), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1218), .ZN(new_n1219));
  NOR2_X1   g794(.A1(G290), .A2(G1986), .ZN(new_n1220));
  NOR3_X1   g795(.A1(new_n1219), .A2(KEYINPUT108), .A3(new_n1220), .ZN(new_n1221));
  AOI211_X1 g796(.A(new_n1217), .B(new_n1221), .C1(KEYINPUT108), .C2(new_n1219), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1217), .ZN(new_n1223));
  OR2_X1    g798(.A1(new_n727), .A2(new_n729), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n727), .A2(new_n729), .ZN(new_n1225));
  XNOR2_X1  g800(.A(new_n841), .B(new_n843), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n775), .B(new_n1177), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1222), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1216), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g805(.A(new_n1217), .B1(new_n1226), .B2(new_n776), .ZN(new_n1231));
  OAI21_X1  g806(.A(KEYINPUT46), .B1(new_n1217), .B2(G1996), .ZN(new_n1232));
  OR3_X1    g807(.A1(new_n1217), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1231), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  XNOR2_X1  g809(.A(new_n1234), .B(KEYINPUT47), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1227), .A2(new_n1226), .ZN(new_n1236));
  AOI21_X1  g811(.A(new_n1225), .B1(new_n1236), .B2(new_n1223), .ZN(new_n1237));
  INV_X1    g812(.A(new_n841), .ZN(new_n1238));
  AOI21_X1  g813(.A(new_n1237), .B1(new_n843), .B2(new_n1238), .ZN(new_n1239));
  AND2_X1   g814(.A1(new_n1239), .A2(KEYINPUT126), .ZN(new_n1240));
  NOR2_X1   g815(.A1(new_n1239), .A2(KEYINPUT126), .ZN(new_n1241));
  NOR3_X1   g816(.A1(new_n1240), .A2(new_n1241), .A3(new_n1217), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n1228), .A2(new_n1223), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1223), .A2(new_n1220), .ZN(new_n1244));
  XNOR2_X1  g819(.A(new_n1244), .B(KEYINPUT48), .ZN(new_n1245));
  AOI211_X1 g820(.A(new_n1235), .B(new_n1242), .C1(new_n1243), .C2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1230), .A2(new_n1246), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g822(.A1(G227), .A2(new_n462), .ZN(new_n1249));
  AOI21_X1  g823(.A(new_n1249), .B1(new_n700), .B2(new_n704), .ZN(new_n1250));
  NAND2_X1  g824(.A1(new_n666), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g825(.A(new_n1251), .B1(new_n932), .B2(new_n936), .ZN(new_n1252));
  INV_X1    g826(.A(KEYINPUT127), .ZN(new_n1253));
  OAI211_X1 g827(.A(new_n1252), .B(new_n1253), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1254));
  INV_X1    g828(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g829(.A(new_n1253), .B1(new_n1026), .B2(new_n1252), .ZN(new_n1256));
  NOR2_X1   g830(.A1(new_n1255), .A2(new_n1256), .ZN(G308));
  NAND2_X1  g831(.A1(new_n1026), .A2(new_n1252), .ZN(new_n1258));
  NAND2_X1  g832(.A1(new_n1258), .A2(KEYINPUT127), .ZN(new_n1259));
  NAND2_X1  g833(.A1(new_n1259), .A2(new_n1254), .ZN(G225));
endmodule


