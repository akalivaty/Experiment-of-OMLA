//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n545, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G238), .A3(G237), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n464), .A2(new_n466), .A3(G137), .A4(new_n462), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n463), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n469), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n464), .A2(new_n466), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n462), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(KEYINPUT66), .A2(G138), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n464), .A2(new_n466), .A3(new_n484), .A4(new_n462), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n462), .A4(new_n484), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(G126), .A3(G2105), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n487), .A2(new_n489), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(G651), .ZN(new_n497));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT67), .A3(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n500), .A2(G50), .A3(G543), .A4(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n500), .A2(G88), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n503), .B(new_n505), .C1(new_n498), .C2(new_n506), .ZN(G303));
  INV_X1    g082(.A(G303), .ZN(G166));
  AOI21_X1  g083(.A(new_n501), .B1(new_n497), .B2(new_n499), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(G51), .A3(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n512));
  INV_X1    g087(.A(G89), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n510), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(KEYINPUT69), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(KEYINPUT69), .B1(new_n516), .B2(new_n517), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n516), .A2(new_n517), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n515), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(new_n525), .A3(new_n518), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n514), .A2(new_n527), .ZN(G168));
  INV_X1    g103(.A(new_n512), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G90), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n500), .A2(G543), .A3(new_n502), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT70), .B(G52), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n498), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n530), .A2(new_n534), .A3(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT71), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  AOI22_X1  g116(.A1(G43), .A2(new_n532), .B1(new_n529), .B2(G81), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n509), .A2(new_n550), .A3(G53), .A4(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT5), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT5), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT74), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G65), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n556), .A2(new_n558), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n563), .A2(KEYINPUT75), .A3(new_n564), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n567), .A2(G651), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT76), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n509), .A2(KEYINPUT73), .A3(new_n504), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT73), .B1(new_n509), .B2(new_n504), .ZN(new_n572));
  OAI21_X1  g147(.A(G91), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n567), .A2(new_n574), .A3(new_n568), .A4(G651), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n554), .A2(new_n570), .A3(new_n573), .A4(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  OAI21_X1  g152(.A(G87), .B1(new_n571), .B2(new_n572), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT78), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n500), .A2(G49), .A3(G543), .A4(new_n502), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n509), .A2(KEYINPUT77), .A3(G49), .A4(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n578), .A2(new_n580), .A3(new_n585), .ZN(G288));
  INV_X1    g161(.A(G48), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n531), .A2(new_n587), .B1(new_n588), .B2(new_n498), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT73), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n512), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n509), .A2(KEYINPUT73), .A3(new_n504), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n589), .B1(new_n593), .B2(G86), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n529), .A2(G85), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n532), .A2(G47), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n596), .B(new_n597), .C1(new_n498), .C2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(G92), .B1(new_n571), .B2(new_n572), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n593), .A2(new_n603), .A3(G92), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n504), .A2(G66), .ZN(new_n605));
  INV_X1    g180(.A(G79), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n555), .ZN(new_n607));
  AOI22_X1  g182(.A1(G54), .A2(new_n532), .B1(new_n607), .B2(G651), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n602), .A2(new_n604), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(KEYINPUT79), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n602), .A2(new_n604), .A3(new_n611), .A4(new_n608), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n600), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n600), .B1(new_n613), .B2(G868), .ZN(G321));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(G299), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n616), .B2(G168), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(new_n616), .B2(G168), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  OAI21_X1  g196(.A(KEYINPUT80), .B1(new_n543), .B2(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n613), .A2(new_n620), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  MUX2_X1   g199(.A(KEYINPUT80), .B(new_n622), .S(new_n624), .Z(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n488), .A2(new_n471), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT13), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n462), .A2(G111), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT81), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n478), .A2(G135), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n476), .A2(G123), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NOR2_X1   g212(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT82), .ZN(G156));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT15), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2435), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  AND2_X1   g226(.A1(new_n651), .A2(G14), .ZN(G401));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n657), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n655), .B2(new_n656), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  INV_X1    g239(.A(new_n655), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n656), .B(KEYINPUT17), .Z(new_n666));
  OAI21_X1  g241(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n657), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n661), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n673), .A2(new_n674), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n678), .A3(new_n680), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n683), .B(new_n684), .C1(new_n682), .C2(new_n681), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT88), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G229));
  INV_X1    g267(.A(KEYINPUT102), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT90), .B(G16), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n543), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n695), .A2(G19), .ZN(new_n697));
  OAI21_X1  g272(.A(KEYINPUT94), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(KEYINPUT94), .B2(new_n697), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(G1341), .Z(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G4), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n613), .B2(new_n701), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT93), .B(G1348), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G26), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n476), .A2(G128), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n478), .A2(G140), .ZN(new_n709));
  OR2_X1    g284(.A1(G104), .A2(G2105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n710), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n707), .B1(new_n713), .B2(new_n706), .ZN(new_n714));
  MUX2_X1   g289(.A(new_n707), .B(new_n714), .S(KEYINPUT28), .Z(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT95), .B(G2067), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n700), .A2(new_n705), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT96), .Z(new_n719));
  AND2_X1   g294(.A1(new_n706), .A2(G33), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n471), .A2(G103), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT25), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n478), .A2(G139), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(KEYINPUT97), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(KEYINPUT97), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n488), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  OAI22_X1  g303(.A1(new_n726), .A2(new_n727), .B1(new_n462), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n720), .B1(new_n729), .B2(G29), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT98), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n731), .ZN(new_n734));
  AND3_X1   g309(.A1(new_n733), .A2(G2072), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(G2072), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(G5), .A2(G16), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G301), .B2(new_n701), .ZN(new_n739));
  INV_X1    g314(.A(G1961), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT31), .B(G11), .Z(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT30), .B(G28), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n742), .B1(new_n706), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n636), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n706), .ZN(new_n746));
  NAND2_X1  g321(.A1(G164), .A2(G29), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G27), .B2(G29), .ZN(new_n748));
  INV_X1    g323(.A(G2078), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n741), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n739), .A2(new_n740), .ZN(new_n752));
  NOR2_X1   g327(.A1(G16), .A2(G21), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G168), .B2(G16), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(G1966), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n751), .A2(new_n752), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G29), .A2(G32), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n478), .A2(G141), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT99), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n471), .A2(G105), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT26), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n761), .B(new_n763), .C1(G129), .C2(new_n476), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n758), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT27), .B(G1996), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(KEYINPUT24), .A2(G34), .ZN(new_n770));
  NAND2_X1  g345(.A1(KEYINPUT24), .A2(G34), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n770), .A2(new_n706), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G160), .B2(new_n706), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2084), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n748), .A2(new_n749), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  NOR4_X1   g351(.A1(new_n757), .A2(new_n769), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n737), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT100), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n737), .A2(new_n777), .A3(KEYINPUT100), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(G299), .A2(G16), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n695), .A2(G20), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT101), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT23), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(G162), .A2(G29), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G29), .B2(G35), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT29), .B(G2090), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n782), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n693), .B1(new_n719), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n794), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n718), .B(KEYINPUT96), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n796), .A2(new_n797), .A3(KEYINPUT102), .ZN(new_n798));
  MUX2_X1   g373(.A(G23), .B(G288), .S(G16), .Z(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT33), .B(G1976), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n695), .A2(G22), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n695), .ZN(new_n803));
  INV_X1    g378(.A(G1971), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n701), .A2(G6), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n594), .B2(new_n701), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT32), .B(G1981), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n801), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT34), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n476), .A2(G119), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n478), .A2(G131), .ZN(new_n813));
  OR2_X1    g388(.A1(G95), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT89), .Z(new_n817));
  MUX2_X1   g392(.A(G25), .B(new_n817), .S(G29), .Z(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT35), .B(G1991), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n818), .B(new_n819), .Z(new_n820));
  MUX2_X1   g395(.A(G24), .B(G290), .S(new_n694), .Z(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT91), .B(G1986), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n811), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(KEYINPUT36), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n824), .A2(new_n826), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n825), .A2(KEYINPUT36), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n795), .A2(new_n798), .B1(new_n829), .B2(new_n830), .ZN(G311));
  OAI21_X1  g406(.A(new_n830), .B1(new_n827), .B2(new_n828), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n719), .A2(new_n693), .A3(new_n794), .ZN(new_n833));
  AOI21_X1  g408(.A(KEYINPUT102), .B1(new_n796), .B2(new_n797), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(G150));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n836), .A2(new_n531), .B1(new_n512), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT103), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(new_n498), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n613), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n543), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n541), .A2(new_n542), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n840), .A2(new_n849), .A3(new_n842), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT39), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n847), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n845), .B1(new_n853), .B2(G860), .ZN(G145));
  XNOR2_X1  g429(.A(new_n729), .B(new_n712), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n765), .B(G164), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n857), .A2(KEYINPUT105), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n476), .A2(G130), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n478), .A2(G142), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n462), .A2(G118), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n628), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n816), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n857), .A2(KEYINPUT105), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n858), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n865), .B(KEYINPUT104), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n857), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n482), .B(G160), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n636), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n867), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n857), .B(new_n868), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n874), .B2(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g452(.A(new_n623), .B(new_n851), .ZN(new_n878));
  XNOR2_X1  g453(.A(G299), .B(new_n609), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n879), .B(KEYINPUT41), .Z(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  XNOR2_X1  g461(.A(G288), .B(G290), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n594), .B(G303), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n885), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n885), .B2(new_n886), .ZN(new_n891));
  OAI21_X1  g466(.A(G868), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n843), .A2(new_n616), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(G295));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n893), .ZN(G331));
  NOR2_X1   g470(.A1(G171), .A2(KEYINPUT106), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(G286), .B1(KEYINPUT106), .B2(G171), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(new_n848), .A3(new_n850), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n848), .B2(new_n850), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n851), .A2(new_n898), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n896), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n879), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n882), .A2(new_n905), .A3(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n889), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n908), .A3(new_n889), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n911), .A2(new_n916), .A3(new_n912), .A4(new_n913), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(KEYINPUT107), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n920), .A3(KEYINPUT43), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n915), .A2(KEYINPUT44), .A3(new_n917), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(G397));
  INV_X1    g499(.A(G1384), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n493), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n926), .B(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT109), .B1(G160), .B2(G40), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n932));
  INV_X1    g507(.A(G40), .ZN(new_n933));
  NOR4_X1   g508(.A1(new_n469), .A2(new_n473), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n936), .A2(KEYINPUT110), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(KEYINPUT110), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT126), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n941));
  OAI22_X1  g516(.A1(new_n939), .A2(G1996), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n937), .A2(new_n938), .ZN(new_n943));
  INV_X1    g518(.A(G2067), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n712), .B(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1996), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n940), .A2(new_n941), .ZN(new_n947));
  NOR2_X1   g522(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n766), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n942), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT47), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n943), .A2(G1996), .A3(new_n765), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT111), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n943), .A2(new_n963), .A3(G1996), .A4(new_n765), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n945), .B1(G1996), .B2(new_n765), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n943), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n817), .A2(new_n819), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n962), .A2(new_n964), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(G2067), .B2(new_n712), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n943), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n962), .A2(new_n964), .ZN(new_n971));
  NOR2_X1   g546(.A1(G290), .A2(G1986), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n943), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT48), .ZN(new_n974));
  INV_X1    g549(.A(new_n816), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n819), .B(KEYINPUT112), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n939), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n975), .B2(new_n976), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n971), .A2(new_n974), .A3(new_n966), .A4(new_n978), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n960), .A2(new_n970), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n467), .A2(new_n468), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(G2105), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n470), .A2(new_n472), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n983), .A3(G40), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n932), .ZN(new_n985));
  NAND3_X1  g560(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n926), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n944), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n493), .B2(new_n925), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n493), .A2(new_n989), .A3(new_n925), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n935), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n988), .B1(new_n992), .B2(G1348), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT60), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n610), .A2(new_n994), .A3(new_n612), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n997));
  NAND2_X1  g572(.A1(new_n985), .A2(new_n986), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n926), .A2(new_n929), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n493), .A2(KEYINPUT45), .A3(new_n925), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n998), .A2(new_n946), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n493), .A2(new_n925), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n931), .B2(new_n934), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT58), .B(G1341), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n997), .B1(new_n1006), .B2(new_n543), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT59), .ZN(new_n1009));
  AOI211_X1 g584(.A(new_n849), .B(new_n1009), .C1(new_n1001), .C2(new_n1005), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n996), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n990), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n493), .A2(new_n989), .A3(new_n925), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n998), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1956), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT56), .B(G2072), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1017), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n563), .A2(KEYINPUT75), .A3(new_n564), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT75), .B1(new_n563), .B2(new_n564), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n574), .B1(new_n1021), .B2(G651), .ZN(new_n1022));
  INV_X1    g597(.A(new_n575), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n552), .A2(new_n553), .B1(new_n593), .B2(G91), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT57), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n570), .A2(new_n575), .ZN(new_n1027));
  INV_X1    g602(.A(new_n553), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n573), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1027), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1016), .B(new_n1018), .C1(new_n1026), .C2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G299), .A2(new_n1031), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1024), .A2(KEYINPUT57), .A3(new_n1025), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n991), .A2(new_n990), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1956), .B1(new_n1036), .B2(new_n998), .ZN(new_n1037));
  AND4_X1   g612(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1017), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1034), .B(new_n1035), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1033), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT61), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n610), .A2(new_n612), .ZN(new_n1043));
  INV_X1    g618(.A(G1348), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1014), .A2(new_n1044), .B1(new_n944), .B2(new_n987), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1348), .B1(new_n1036), .B2(new_n998), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1003), .A2(G2067), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n610), .B(new_n612), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT60), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1033), .A2(new_n1039), .A3(KEYINPUT61), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1011), .A2(new_n1042), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1039), .A2(new_n1049), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1033), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT120), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n514), .B2(new_n527), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT121), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1061), .B(G8), .C1(new_n514), .C2(new_n527), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT51), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1066));
  INV_X1    g641(.A(G1966), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G2084), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1036), .A2(new_n1069), .A3(new_n998), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1064), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1063), .A2(KEYINPUT51), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1072), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n992), .A2(new_n1069), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1074), .B(new_n1075), .C1(new_n1076), .C2(new_n1065), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(new_n1072), .ZN(new_n1080));
  AOI221_X4 g655(.A(KEYINPUT122), .B1(new_n1062), .B2(new_n1059), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1073), .B(new_n1077), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT49), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n589), .B1(G86), .B2(new_n529), .ZN(new_n1084));
  INV_X1    g659(.A(G1981), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g661(.A(G1981), .B(new_n589), .C1(G86), .C2(new_n593), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n594), .A2(new_n1085), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1089), .B(KEYINPUT49), .C1(new_n1085), .C2(new_n1084), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1065), .B1(new_n998), .B2(new_n1002), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1976), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT116), .B1(G288), .B2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n593), .A2(G87), .B1(new_n583), .B2(new_n584), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(G1976), .A4(new_n580), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT52), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1092), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1000), .B1(new_n931), .B2(new_n934), .ZN(new_n1101));
  INV_X1    g676(.A(new_n999), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n804), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G2090), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1036), .A2(new_n1104), .A3(new_n998), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1065), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(G303), .A2(G8), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT55), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(G303), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1106), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n1116));
  NAND2_X1  g691(.A1(G288), .A2(new_n1093), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g694(.A(KEYINPUT117), .B(KEYINPUT52), .C1(G288), .C2(new_n1093), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1098), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1100), .A2(new_n1115), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT114), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1114), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1109), .A2(new_n1112), .A3(KEYINPUT114), .A4(new_n1113), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1106), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT115), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1106), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1066), .A2(G2078), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1132), .A2(new_n1133), .B1(new_n740), .B2(new_n1014), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1066), .A2(G2078), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT53), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G301), .B(KEYINPUT54), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1082), .A2(new_n1122), .A3(new_n1131), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1134), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n930), .A2(KEYINPUT53), .A3(new_n1000), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1142), .A2(G2078), .A3(new_n984), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1141), .A2(new_n1143), .A3(new_n1138), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1053), .A2(new_n1146), .A3(new_n1055), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1057), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1089), .B1(new_n1150), .B2(G288), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1091), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1121), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1153), .A2(new_n1099), .A3(new_n1092), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1152), .B1(new_n1131), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1122), .A2(new_n1131), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1071), .A2(G168), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT118), .B1(new_n1154), .B2(new_n1115), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1122), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1071), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1163), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1160), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1155), .B1(new_n1159), .B2(new_n1165), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1148), .A2(new_n1149), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1149), .B1(new_n1148), .B2(new_n1166), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1082), .A2(KEYINPUT62), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1169), .A2(G171), .A3(new_n1137), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1131), .B(new_n1122), .C1(new_n1082), .C2(KEYINPUT62), .ZN(new_n1171));
  OR3_X1    g746(.A1(new_n1170), .A2(KEYINPUT125), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(KEYINPUT125), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1167), .A2(new_n1168), .A3(new_n1174), .ZN(new_n1175));
  AND2_X1   g750(.A1(G290), .A2(G1986), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n943), .B1(new_n972), .B2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n971), .A2(new_n1177), .A3(new_n966), .A4(new_n978), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n980), .B1(new_n1175), .B2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g754(.A(G229), .B1(new_n651), .B2(G14), .ZN(new_n1181));
  AOI211_X1 g755(.A(new_n460), .B(G227), .C1(new_n873), .C2(new_n875), .ZN(new_n1182));
  NAND4_X1  g756(.A1(new_n918), .A2(new_n1181), .A3(new_n921), .A4(new_n1182), .ZN(G225));
  INV_X1    g757(.A(G225), .ZN(G308));
endmodule


