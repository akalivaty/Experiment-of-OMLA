//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT65), .B(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n214), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT1), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n212), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n213), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT64), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT0), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n231), .B(new_n235), .C1(new_n230), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n217), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT66), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(G68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n227), .A2(G50), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n248), .B(new_n253), .ZN(G351));
  AOI21_X1  g0054(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G274), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n255), .A2(new_n260), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n262), .B1(G226), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G222), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G223), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n270), .B(new_n255), .C1(G77), .C2(new_n266), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G179), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(G169), .B2(new_n272), .ZN(new_n275));
  INV_X1    g0075(.A(G1), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G13), .A3(G20), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G50), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n214), .A2(KEYINPUT67), .A3(G33), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n280), .B1(new_n213), .B2(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n279), .A2(new_n209), .A3(new_n282), .A4(new_n277), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n210), .A2(G1), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n283), .A2(new_n202), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n281), .A2(G20), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n287), .A2(new_n288), .B1(G150), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n290), .A2(new_n291), .B1(G20), .B2(new_n203), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n291), .B2(new_n290), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n279), .A2(new_n209), .A3(new_n282), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n278), .B(new_n285), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n275), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n295), .B(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n272), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(G190), .B2(new_n272), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n298), .A2(new_n304), .A3(new_n301), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n296), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n262), .B1(G244), .B2(new_n264), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n266), .A2(new_n268), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n308), .A2(new_n217), .B1(new_n222), .B2(new_n266), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n266), .A2(G1698), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n226), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n255), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT69), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT69), .B1(new_n307), .B2(new_n312), .ZN(new_n316));
  OAI21_X1  g0116(.A(G190), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  INV_X1    g0118(.A(new_n289), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n286), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n318), .B2(new_n319), .ZN(new_n321));
  INV_X1    g0121(.A(new_n288), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT15), .B(G87), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n321), .B1(new_n210), .B2(new_n218), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n277), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n324), .A2(new_n294), .B1(new_n218), .B2(new_n325), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n283), .A2(new_n218), .A3(new_n284), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n315), .A2(new_n316), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n317), .B(new_n330), .C1(new_n332), .C2(new_n299), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n332), .B2(new_n273), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n306), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n325), .A2(new_n227), .ZN(new_n339));
  XOR2_X1   g0139(.A(new_n339), .B(KEYINPUT12), .Z(new_n340));
  AOI22_X1  g0140(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n227), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n322), .B2(new_n218), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n342), .A2(new_n294), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n340), .B1(KEYINPUT11), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(KEYINPUT11), .B2(new_n343), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n283), .A2(new_n227), .A3(new_n284), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT72), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT3), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G33), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G1698), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT71), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n353), .A2(new_n268), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(G232), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n310), .A2(KEYINPUT71), .A3(new_n217), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n255), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n262), .B1(G238), .B2(new_n264), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT13), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(new_n365), .A3(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT14), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n368), .A3(G169), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n273), .B2(new_n367), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n368), .B1(new_n367), .B2(G169), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n349), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n348), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n299), .B1(new_n364), .B2(new_n366), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n338), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n283), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n286), .A2(new_n284), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n380), .A2(new_n381), .B1(new_n325), .B2(new_n286), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n294), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n216), .A2(new_n227), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n385), .A2(new_n201), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(G20), .B1(G159), .B2(new_n289), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n353), .A2(KEYINPUT73), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT73), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n350), .A2(new_n352), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n210), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT74), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n266), .A2(new_n393), .A3(G20), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n395), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n388), .B1(new_n400), .B2(G68), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n384), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n350), .A2(KEYINPUT75), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n352), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n350), .A2(KEYINPUT75), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT7), .B(new_n210), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n393), .B1(new_n266), .B2(G20), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n387), .B1(new_n408), .B2(new_n227), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n383), .B1(new_n402), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n255), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n268), .A2(G223), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n266), .A2(new_n414), .B1(G33), .B2(G87), .ZN(new_n415));
  AND2_X1   g0215(.A1(G226), .A2(G1698), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT76), .B1(new_n266), .B2(new_n416), .ZN(new_n417));
  AND4_X1   g0217(.A1(KEYINPUT76), .A2(new_n350), .A3(new_n352), .A4(new_n416), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT77), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n415), .B(KEYINPUT77), .C1(new_n417), .C2(new_n418), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n413), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n261), .B1(new_n217), .B2(new_n263), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(new_n299), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(G190), .B2(new_n425), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n412), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n412), .A2(KEYINPUT17), .A3(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n424), .A2(G179), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT78), .B1(new_n423), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n335), .B1(new_n423), .B2(new_n424), .ZN(new_n435));
  INV_X1    g0235(.A(new_n422), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n350), .A2(new_n352), .A3(new_n416), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT76), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n266), .A2(KEYINPUT76), .A3(new_n416), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT77), .B1(new_n441), .B2(new_n415), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n255), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT78), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n424), .A2(G179), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n434), .A2(new_n435), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n434), .A2(new_n435), .A3(new_n446), .A4(KEYINPUT79), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT18), .B1(new_n451), .B2(new_n412), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n392), .A2(new_n396), .A3(new_n393), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n396), .B1(new_n392), .B2(new_n393), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n453), .A2(new_n454), .A3(new_n398), .ZN(new_n455));
  OAI211_X1 g0255(.A(KEYINPUT16), .B(new_n387), .C1(new_n455), .C2(new_n227), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(new_n411), .A3(new_n294), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n382), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT18), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(new_n449), .A4(new_n450), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n452), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n452), .A2(KEYINPUT80), .A3(new_n460), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n432), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n379), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n281), .A2(G1), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n283), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G116), .ZN(new_n469));
  AOI21_X1  g0269(.A(G20), .B1(G33), .B2(G283), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n281), .A2(G97), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n470), .A2(new_n471), .B1(G20), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT20), .B1(new_n294), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n294), .A2(KEYINPUT20), .A3(new_n473), .ZN(new_n475));
  OAI221_X1 g0275(.A(new_n469), .B1(G116), .B2(new_n277), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n266), .A2(G257), .A3(new_n268), .ZN(new_n477));
  INV_X1    g0277(.A(G303), .ZN(new_n478));
  OAI221_X1 g0278(.A(new_n477), .B1(new_n478), .B2(new_n266), .C1(new_n310), .C2(new_n223), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n255), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT84), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n258), .A3(KEYINPUT5), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(KEYINPUT84), .B2(G41), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n259), .A2(G1), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n257), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n255), .B1(new_n486), .B2(new_n482), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G270), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n480), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n476), .A2(G169), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n490), .A2(new_n273), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n476), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n476), .A2(KEYINPUT21), .A3(new_n490), .A4(G169), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT23), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n210), .B2(G107), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n222), .A2(KEYINPUT23), .A3(G20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G116), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n499), .A2(new_n500), .B1(new_n502), .B2(new_n210), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n266), .A2(new_n210), .A3(G87), .ZN(new_n504));
  XOR2_X1   g0304(.A(KEYINPUT90), .B(KEYINPUT22), .Z(new_n505));
  AND2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n504), .A2(new_n505), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n384), .B1(new_n508), .B2(new_n509), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n283), .A2(new_n222), .A3(new_n467), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n325), .A2(KEYINPUT25), .A3(new_n222), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT25), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n277), .B2(G107), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(KEYINPUT91), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT91), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n517), .B(new_n514), .C1(new_n277), .C2(G107), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OR3_X1    g0319(.A1(new_n512), .A2(new_n519), .A3(KEYINPUT92), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT92), .B1(new_n512), .B2(new_n519), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n510), .A2(new_n511), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n266), .A2(G257), .A3(G1698), .ZN(new_n523));
  INV_X1    g0323(.A(G294), .ZN(new_n524));
  INV_X1    g0324(.A(G250), .ZN(new_n525));
  OAI221_X1 g0325(.A(new_n523), .B1(new_n281), .B2(new_n524), .C1(new_n308), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n255), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n488), .A2(G264), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n487), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n335), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(G179), .B2(new_n529), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n522), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n497), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n510), .A2(new_n511), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n520), .A2(new_n521), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n529), .A2(G200), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n373), .B2(new_n529), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n490), .A2(G200), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n490), .A2(new_n373), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n541), .A2(new_n542), .A3(new_n476), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n534), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n266), .A2(G238), .A3(new_n268), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(new_n501), .C1(new_n310), .C2(new_n219), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT87), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n357), .A2(G244), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT87), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n548), .A2(new_n549), .A3(new_n545), .A4(new_n501), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n413), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n413), .B(G250), .C1(G1), .C2(new_n259), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n257), .A2(new_n485), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n273), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n266), .A2(new_n210), .A3(G68), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT88), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT19), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n288), .A2(new_n559), .A3(G97), .ZN(new_n560));
  AOI21_X1  g0360(.A(G20), .B1(G33), .B2(G97), .ZN(new_n561));
  INV_X1    g0361(.A(G87), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G97), .A2(G107), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n560), .B1(new_n564), .B2(new_n559), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n558), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n557), .A2(KEYINPUT88), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n294), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n323), .A2(new_n325), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n323), .B(KEYINPUT89), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n468), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n335), .B1(new_n551), .B2(new_n554), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n556), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n554), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n547), .A2(new_n550), .ZN(new_n576));
  OAI211_X1 g0376(.A(G190), .B(new_n575), .C1(new_n576), .C2(new_n413), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n568), .A2(new_n569), .ZN(new_n578));
  INV_X1    g0378(.A(new_n468), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n562), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n577), .B(new_n581), .C1(new_n299), .C2(new_n555), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n574), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g0384(.A(G97), .B(G107), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT6), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G97), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n586), .A2(new_n588), .A3(G107), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n590), .A2(new_n210), .B1(new_n218), .B2(new_n319), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n222), .B1(new_n406), .B2(new_n407), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n294), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n468), .A2(G97), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n593), .B(new_n594), .C1(G97), .C2(new_n277), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n354), .A2(KEYINPUT81), .A3(G244), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n266), .A2(G244), .A3(new_n268), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT81), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g0399(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT4), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT83), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  OR3_X1    g0403(.A1(new_n597), .A2(KEYINPUT83), .A3(new_n602), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n357), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n601), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n255), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n488), .A2(G257), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n487), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n609), .A2(KEYINPUT85), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(KEYINPUT85), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n595), .B1(G200), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n606), .B2(new_n255), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n373), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT86), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n607), .A2(new_n610), .A3(new_n273), .A4(new_n611), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n595), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n614), .A2(G169), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OR2_X1    g0421(.A1(new_n614), .A2(G169), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n622), .A2(KEYINPUT86), .A3(new_n618), .A4(new_n595), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n616), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n544), .A2(new_n584), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n466), .A2(new_n626), .ZN(G372));
  INV_X1    g0427(.A(KEYINPUT93), .ZN(new_n628));
  INV_X1    g0428(.A(new_n447), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n458), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT18), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n458), .A2(new_n459), .A3(new_n629), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n376), .B1(new_n372), .B2(new_n337), .ZN(new_n634));
  INV_X1    g0434(.A(new_n432), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n303), .A2(new_n305), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n628), .B1(new_n638), .B2(new_n296), .ZN(new_n639));
  OAI221_X1 g0439(.A(KEYINPUT93), .B1(new_n295), .B2(new_n275), .C1(new_n636), .C2(new_n637), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n466), .ZN(new_n642));
  INV_X1    g0442(.A(new_n574), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n622), .A2(new_n618), .A3(new_n595), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n583), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n583), .B1(new_n621), .B2(new_n623), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n647), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n540), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(new_n532), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n624), .A2(new_n652), .A3(new_n583), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n642), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n641), .A2(new_n655), .ZN(G369));
  NAND3_X1  g0456(.A1(new_n276), .A2(new_n210), .A3(G13), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n476), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n497), .B(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n543), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  INV_X1    g0467(.A(new_n662), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n522), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n533), .B1(new_n669), .B2(new_n540), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n532), .A2(new_n668), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n497), .A2(new_n662), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n670), .A2(new_n675), .B1(new_n532), .B2(new_n668), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n232), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n563), .A2(new_n562), .A3(new_n472), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n679), .A2(new_n680), .A3(new_n276), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n208), .B2(new_n679), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT28), .Z(new_n683));
  INV_X1    g0483(.A(KEYINPUT29), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n684), .B(new_n668), .C1(new_n649), .C2(new_n653), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n648), .A2(new_n646), .ZN(new_n686));
  INV_X1    g0486(.A(new_n619), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n687), .A2(new_n574), .A3(new_n582), .A4(new_n622), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n643), .B1(new_n688), .B2(KEYINPUT26), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT96), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n653), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n686), .A2(new_n689), .A3(KEYINPUT96), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n662), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n685), .B1(new_n694), .B2(new_n684), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n527), .A2(new_n528), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n490), .A2(new_n696), .A3(new_n273), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(new_n555), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT30), .A4(new_n614), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(new_n555), .A3(new_n614), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT94), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n490), .A2(new_n529), .A3(new_n273), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n705), .B(new_n612), .C1(new_n551), .C2(new_n554), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n700), .A2(new_n703), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT31), .B1(new_n707), .B2(new_n662), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT95), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n544), .A2(new_n584), .A3(new_n625), .A4(new_n668), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n662), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT95), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n710), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n717), .A2(G330), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n695), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT97), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT97), .B1(new_n695), .B2(new_n718), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n683), .B1(new_n723), .B2(G1), .ZN(G364));
  INV_X1    g0524(.A(new_n666), .ZN(new_n725));
  INV_X1    g0525(.A(G330), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT98), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n210), .A2(G13), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n276), .B1(new_n729), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n679), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n667), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n725), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n209), .B1(G20), .B2(new_n335), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n373), .A2(G179), .A3(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n210), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n588), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n210), .A2(new_n273), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n373), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n743), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n747), .A2(G190), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n266), .B1(new_n746), .B2(new_n202), .C1(new_n218), .C2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n744), .A2(G190), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n742), .B(new_n750), .C1(G68), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n743), .A2(G190), .A3(new_n299), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT100), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT32), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n210), .A2(G190), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(new_n273), .A3(new_n299), .ZN(new_n759));
  INV_X1    g0559(.A(G159), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n759), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(KEYINPUT32), .A3(G159), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n756), .A2(G58), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT101), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(new_n299), .B2(G179), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n210), .A2(new_n373), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n273), .A2(KEYINPUT101), .A3(G200), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G87), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n766), .A2(new_n758), .A3(new_n768), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G107), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n752), .A2(new_n764), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(KEYINPUT102), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  INV_X1    g0577(.A(G329), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n749), .A2(new_n777), .B1(new_n759), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n753), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n266), .B(new_n779), .C1(G322), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n741), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G294), .A2(new_n782), .B1(new_n745), .B2(G326), .ZN(new_n783));
  INV_X1    g0583(.A(new_n751), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT103), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n786), .B2(new_n785), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G303), .A2(new_n770), .B1(new_n773), .B2(G283), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n781), .A2(new_n783), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n776), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n775), .A2(KEYINPUT102), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n739), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n737), .A2(new_n739), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n253), .A2(new_n259), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n389), .A2(new_n391), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n678), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n795), .B(new_n798), .C1(new_n259), .C2(new_n208), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n678), .A2(new_n353), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n800), .A2(G355), .B1(new_n472), .B2(new_n678), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  OAI21_X1  g0602(.A(new_n794), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n738), .A2(new_n793), .A3(new_n803), .A4(new_n732), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n734), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  OAI21_X1  g0606(.A(new_n668), .B1(new_n649), .B2(new_n653), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n329), .A2(new_n662), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n333), .A2(new_n808), .B1(new_n334), .B2(new_n336), .ZN(new_n809));
  AND3_X1   g0609(.A1(new_n334), .A2(new_n336), .A3(new_n668), .ZN(new_n810));
  OAI21_X1  g0610(.A(KEYINPUT105), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n333), .A2(new_n808), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n337), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT105), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n334), .A2(new_n336), .A3(new_n668), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n807), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n811), .A2(new_n816), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n654), .A2(new_n819), .A3(new_n668), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n718), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n732), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n718), .A2(new_n818), .A3(new_n820), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n739), .A2(new_n735), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(G77), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n796), .B1(new_n828), .B2(new_n759), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n773), .A2(G68), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n202), .B2(new_n769), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(G58), .C2(new_n782), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT104), .Z(new_n833));
  AOI22_X1  g0633(.A1(G159), .A2(new_n748), .B1(new_n745), .B2(G137), .ZN(new_n834));
  INV_X1    g0634(.A(G150), .ZN(new_n835));
  INV_X1    g0635(.A(G143), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n784), .C1(new_n755), .C2(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT34), .Z(new_n838));
  AOI21_X1  g0638(.A(new_n742), .B1(G303), .B2(new_n745), .ZN(new_n839));
  INV_X1    g0639(.A(G283), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n840), .B2(new_n784), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n749), .A2(new_n472), .B1(new_n759), .B2(new_n777), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n266), .B(new_n842), .C1(G294), .C2(new_n780), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n773), .A2(G87), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n770), .A2(G107), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n833), .A2(new_n838), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n733), .B(new_n827), .C1(new_n847), .C2(new_n739), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n819), .B2(new_n736), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n824), .A2(new_n849), .ZN(G384));
  INV_X1    g0650(.A(new_n590), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n851), .A2(KEYINPUT35), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(KEYINPUT35), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n852), .A2(G116), .A3(new_n211), .A4(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT36), .Z(new_n855));
  OR3_X1    g0655(.A1(new_n207), .A2(new_n218), .A3(new_n385), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n276), .B(G13), .C1(new_n856), .C2(new_n249), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n660), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n458), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n428), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n451), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT37), .B1(new_n862), .B2(new_n458), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n398), .B1(new_n394), .B2(KEYINPUT74), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n227), .B1(new_n864), .B2(new_n397), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n410), .B1(new_n865), .B2(new_n388), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n456), .A3(new_n294), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n382), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n859), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n629), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n870), .A3(new_n428), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n861), .A2(new_n863), .B1(new_n871), .B2(KEYINPUT37), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n465), .B2(new_n869), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(KEYINPUT38), .B(new_n873), .C1(new_n465), .C2(new_n869), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(KEYINPUT39), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n452), .A2(KEYINPUT80), .A3(new_n460), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT80), .B1(new_n452), .B2(new_n460), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n635), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n869), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n875), .B(new_n872), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n458), .B(new_n859), .C1(new_n432), .C2(new_n633), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n863), .A2(new_n861), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n428), .A2(new_n630), .A3(new_n860), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n879), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n372), .A2(new_n662), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n878), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n859), .B1(new_n631), .B2(new_n632), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n876), .A2(new_n877), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n348), .A2(new_n668), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n378), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n372), .B(new_n377), .C1(new_n348), .C2(new_n668), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n820), .B2(new_n815), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n895), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n894), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT106), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n695), .A2(new_n642), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n641), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n905), .B(new_n907), .Z(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n885), .A2(new_n889), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n875), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n877), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n711), .A2(new_n714), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n819), .A3(new_n900), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n909), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n914), .A2(new_n819), .A3(new_n900), .A4(new_n909), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n876), .B2(new_n877), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n642), .A2(new_n914), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(G330), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n908), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n276), .B2(new_n729), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n908), .A2(new_n924), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n858), .B1(new_n926), .B2(new_n927), .ZN(G367));
  OAI221_X1 g0728(.A(new_n794), .B1(new_n232), .B2(new_n323), .C1(new_n798), .C2(new_n243), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n733), .B1(new_n929), .B2(KEYINPUT108), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(KEYINPUT108), .B2(new_n929), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n266), .B1(new_n835), .B2(new_n753), .C1(new_n749), .C2(new_n202), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(G77), .B2(new_n773), .ZN(new_n933));
  INV_X1    g0733(.A(G137), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n769), .A2(new_n216), .B1(new_n759), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT109), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n784), .A2(new_n760), .B1(new_n746), .B2(new_n836), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n741), .A2(new_n227), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n933), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n935), .A2(KEYINPUT109), .ZN(new_n941));
  INV_X1    g0741(.A(G317), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n749), .A2(new_n840), .B1(new_n759), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n772), .A2(new_n588), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n943), .A2(new_n796), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n478), .B2(new_n755), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n784), .A2(new_n524), .B1(new_n746), .B2(new_n777), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G107), .B2(new_n782), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n770), .A2(KEYINPUT46), .A3(G116), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT46), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n769), .B2(new_n472), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n940), .A2(new_n941), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT47), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n931), .B1(new_n954), .B2(new_n739), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n662), .B1(new_n578), .B2(new_n580), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n584), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n574), .B2(new_n956), .ZN(new_n958));
  INV_X1    g0758(.A(new_n737), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n595), .A2(new_n662), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n625), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n687), .A2(new_n622), .A3(new_n662), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(new_n676), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n676), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n966), .A2(new_n674), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n674), .B1(new_n966), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n672), .B(new_n675), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n667), .B(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n972), .A2(new_n974), .B1(new_n721), .B2(new_n722), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT107), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n679), .B(KEYINPUT41), .Z(new_n977));
  OR3_X1    g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n976), .B1(new_n975), .B2(new_n977), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n731), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n672), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n964), .A2(new_n981), .A3(new_n675), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT42), .Z(new_n983));
  AOI21_X1  g0783(.A(new_n533), .B1(new_n962), .B2(new_n963), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n621), .A2(new_n623), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n668), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n983), .A2(new_n986), .B1(KEYINPUT43), .B2(new_n958), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n987), .B(new_n988), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n673), .A2(new_n964), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n960), .B1(new_n980), .B2(new_n991), .ZN(G387));
  INV_X1    g0792(.A(new_n974), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n721), .B2(new_n722), .ZN(new_n994));
  INV_X1    g0794(.A(new_n679), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n723), .B2(new_n974), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n796), .B1(new_n746), .B2(new_n760), .C1(new_n286), .C2(new_n784), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n570), .A2(new_n782), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n218), .B2(new_n769), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G50), .A2(new_n780), .B1(new_n762), .B2(G150), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n227), .B2(new_n749), .ZN(new_n1002));
  NOR4_X1   g0802(.A1(new_n998), .A2(new_n1000), .A3(new_n1002), .A4(new_n944), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G283), .A2(new_n782), .B1(new_n770), .B2(G294), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n755), .A2(new_n942), .B1(new_n478), .B2(new_n749), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT110), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(KEYINPUT110), .B1(new_n749), .B2(new_n478), .C1(new_n755), .C2(new_n942), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G311), .A2(new_n751), .B1(new_n745), .B2(G322), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT48), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1004), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT111), .Z(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT49), .Z(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT112), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n796), .B1(G326), .B2(new_n762), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n472), .B2(new_n772), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n1016), .B2(KEYINPUT112), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1003), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n739), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n286), .A2(G50), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT50), .ZN(new_n1025));
  AOI211_X1 g0825(.A(G45), .B(new_n680), .C1(G68), .C2(G77), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n798), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n259), .B2(new_n240), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n800), .A2(new_n680), .B1(new_n222), .B2(new_n678), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n733), .B1(new_n1030), .B2(new_n794), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n981), .B2(new_n959), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1023), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT113), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n997), .B(new_n1034), .C1(new_n730), .C2(new_n993), .ZN(G393));
  AOI21_X1  g0835(.A(new_n995), .B1(new_n994), .B2(new_n972), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n994), .B2(new_n972), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n972), .A2(new_n731), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n794), .B1(new_n588), .B2(new_n232), .C1(new_n798), .C2(new_n247), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT114), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n732), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n1040), .B2(new_n1039), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n353), .B1(new_n749), .B2(new_n524), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G322), .B2(new_n762), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G116), .A2(new_n782), .B1(new_n751), .B2(G303), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n770), .A2(G283), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1046), .A2(new_n774), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G317), .A2(new_n745), .B1(new_n780), .B2(G311), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G150), .A2(new_n745), .B1(new_n780), .B2(G159), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT51), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n741), .A2(new_n218), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G50), .B2(new_n751), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n748), .A2(new_n287), .B1(G143), .B2(new_n762), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(new_n796), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n844), .B1(new_n227), .B2(new_n769), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1054), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1052), .A2(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1044), .A2(KEYINPUT115), .B1(new_n739), .B2(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(KEYINPUT115), .B2(new_n1044), .C1(new_n964), .C2(new_n959), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1037), .A2(new_n1038), .A3(new_n1063), .ZN(G390));
  AOI21_X1  g0864(.A(new_n810), .B1(new_n694), .B2(new_n819), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n892), .B(new_n912), .C1(new_n1065), .C2(new_n901), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n717), .A2(G330), .A3(new_n819), .A4(new_n900), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n914), .A2(G330), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n819), .A2(new_n900), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT116), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1068), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(KEYINPUT39), .B1(new_n877), .B2(new_n911), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n882), .A2(new_n883), .ZN(new_n1076));
  AOI21_X1  g0876(.A(KEYINPUT38), .B1(new_n1076), .B2(new_n873), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n884), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1078), .B2(KEYINPUT39), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n815), .B1(new_n807), .B2(new_n817), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n893), .B1(new_n1080), .B2(new_n900), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1066), .B(new_n1074), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1072), .A2(KEYINPUT116), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1081), .B1(new_n878), .B2(new_n891), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n690), .A2(new_n691), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n653), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n1086), .A3(new_n693), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(new_n668), .A3(new_n819), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n901), .B1(new_n1088), .B2(new_n815), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n872), .B1(new_n882), .B2(new_n883), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n890), .B1(new_n1090), .B2(KEYINPUT38), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1089), .A2(new_n1091), .A3(new_n893), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1083), .B1(new_n1084), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1082), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(KEYINPUT117), .B1(new_n1094), .B2(new_n730), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT117), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1082), .A2(new_n1093), .A3(new_n1096), .A4(new_n731), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n466), .A2(new_n1069), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n906), .A2(new_n641), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n717), .A2(G330), .A3(new_n819), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1101), .A2(new_n901), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1080), .B1(new_n1102), .B2(new_n1071), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n901), .B1(new_n1069), .B2(new_n817), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1065), .A2(new_n1104), .A3(new_n1067), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1100), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1094), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n1082), .A3(new_n1093), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n679), .A3(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1079), .A2(new_n736), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n749), .A2(new_n588), .B1(new_n759), .B2(new_n524), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n266), .B(new_n1112), .C1(G116), .C2(new_n780), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1113), .A2(new_n771), .A3(new_n830), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1055), .B1(G283), .B2(new_n745), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n222), .B2(new_n784), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n770), .A2(G150), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT53), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n784), .A2(new_n934), .B1(new_n760), .B2(new_n741), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G128), .B2(new_n745), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n773), .A2(G50), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n353), .B1(new_n748), .B2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G132), .A2(new_n780), .B1(new_n762), .B2(G125), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1120), .A2(new_n1121), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1114), .A2(new_n1116), .B1(new_n1118), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n739), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1128), .B(new_n732), .C1(new_n287), .C2(new_n826), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1111), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT118), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1098), .A2(new_n1110), .A3(new_n1131), .ZN(G378));
  OAI21_X1  g0932(.A(KEYINPUT40), .B1(new_n1091), .B2(new_n915), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n909), .B(new_n916), .C1(new_n1077), .C2(new_n884), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n726), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n904), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(G330), .B1(new_n917), .B2(new_n919), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n894), .A3(new_n903), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1140));
  XNOR2_X1  g0940(.A(new_n306), .B(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n295), .A2(new_n660), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT119), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1141), .B(new_n1143), .Z(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1136), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n731), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n733), .B1(new_n202), .B2(new_n825), .ZN(new_n1149));
  INV_X1    g0949(.A(G128), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n749), .A2(new_n934), .B1(new_n753), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G132), .B2(new_n751), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G150), .A2(new_n782), .B1(new_n745), .B2(G125), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(new_n769), .C2(new_n1122), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n773), .A2(G159), .ZN(new_n1157));
  AOI211_X1 g0957(.A(G33), .B(G41), .C1(new_n762), .C2(G124), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n570), .A2(new_n748), .B1(G58), .B2(new_n773), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n258), .B1(new_n753), .B2(new_n222), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G283), .B2(new_n762), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(new_n218), .C2(new_n769), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n784), .A2(new_n588), .B1(new_n746), .B2(new_n472), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1163), .A2(new_n796), .A3(new_n938), .A4(new_n1164), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(KEYINPUT58), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(KEYINPUT58), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n796), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n258), .B1(new_n1168), .B2(new_n281), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n202), .ZN(new_n1170));
  AND4_X1   g0970(.A1(new_n1159), .A2(new_n1166), .A3(new_n1167), .A4(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1149), .B1(new_n1022), .B2(new_n1171), .C1(new_n1144), .C2(new_n736), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1148), .A2(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n906), .A2(new_n641), .A3(new_n1099), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1109), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1175), .A2(new_n1146), .A3(KEYINPUT57), .A4(new_n1147), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n679), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1136), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1144), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT57), .B1(new_n1180), .B2(new_n1175), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1173), .B1(new_n1177), .B2(new_n1181), .ZN(G375));
  AOI21_X1  g0982(.A(new_n1071), .B1(new_n901), .B2(new_n1101), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1080), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1105), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(new_n1174), .ZN(new_n1186));
  OR3_X1    g0986(.A1(new_n1186), .A2(new_n1106), .A3(new_n977), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n732), .B1(G68), .B2(new_n826), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n749), .A2(new_n222), .B1(new_n784), .B2(new_n472), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT121), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n746), .A2(new_n524), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n353), .B1(new_n759), .B2(new_n478), .C1(new_n753), .C2(new_n840), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n1190), .B2(new_n1189), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n999), .B1(new_n218), .B2(new_n772), .C1(new_n588), .C2(new_n769), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G150), .A2(new_n748), .B1(new_n782), .B2(G50), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT122), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT122), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1168), .B1(G128), .B2(new_n762), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G132), .A2(new_n745), .B1(new_n751), .B2(new_n1123), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n756), .A2(G137), .B1(G58), .B2(new_n773), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n760), .B2(new_n769), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n1195), .A2(new_n1196), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1188), .B1(new_n1206), .B2(new_n739), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT123), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n901), .A2(new_n735), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1209), .B2(KEYINPUT120), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(KEYINPUT120), .B2(new_n1209), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1185), .B2(new_n731), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1187), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(G381));
  NAND3_X1  g1014(.A1(new_n1175), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT57), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n679), .A3(new_n1176), .ZN(new_n1218));
  INV_X1    g1018(.A(G378), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1218), .A2(new_n1219), .A3(new_n1173), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G393), .A2(G396), .ZN(new_n1221));
  INV_X1    g1021(.A(G390), .ZN(new_n1222));
  INV_X1    g1022(.A(G384), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .A4(new_n1213), .ZN(new_n1224));
  OR3_X1    g1024(.A1(new_n1220), .A2(new_n1224), .A3(G387), .ZN(G407));
  INV_X1    g1025(.A(G213), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(G343), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1220), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT124), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G213), .B(G407), .C1(new_n1231), .C2(new_n1232), .ZN(G409));
  NAND2_X1  g1033(.A1(G375), .A2(G378), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT60), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1185), .B2(new_n1174), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(new_n1186), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1103), .A2(new_n1100), .A3(KEYINPUT60), .A4(new_n1105), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n679), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1212), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1223), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G384), .B(new_n1212), .C1(new_n1237), .C2(new_n1239), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n977), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1175), .A2(new_n1146), .A3(new_n1244), .A4(new_n1147), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1245), .A2(new_n1148), .A3(new_n1172), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1227), .B1(new_n1246), .B2(new_n1219), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1234), .A2(new_n1243), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT62), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT61), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT126), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1227), .A2(G2897), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1241), .A2(new_n1251), .A3(new_n1242), .A4(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1241), .A2(new_n1251), .A3(new_n1242), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1252), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1251), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1254), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1246), .A2(new_n1219), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1228), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1219), .B1(new_n1218), .B2(new_n1173), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1234), .A2(new_n1247), .A3(new_n1263), .A4(new_n1243), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1249), .A2(new_n1250), .A3(new_n1262), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G387), .A2(new_n1222), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G390), .B(new_n960), .C1(new_n980), .C2(new_n991), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(new_n805), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT127), .B1(G387), .B2(new_n1222), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1268), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1269), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1272), .A2(new_n1266), .A3(KEYINPUT127), .A4(new_n1267), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1265), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1234), .A2(new_n1247), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT61), .B1(new_n1277), .B2(new_n1258), .ZN(new_n1278));
  XOR2_X1   g1078(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1279));
  NAND2_X1  g1079(.A1(new_n1248), .A2(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1234), .A2(new_n1247), .A3(KEYINPUT63), .A4(new_n1243), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1276), .A2(new_n1278), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1275), .A2(new_n1282), .ZN(G405));
  INV_X1    g1083(.A(new_n1220), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1243), .B1(new_n1284), .B2(new_n1261), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1243), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1234), .A2(new_n1220), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(new_n1276), .ZN(G402));
endmodule


