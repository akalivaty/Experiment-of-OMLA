//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n213), .B(new_n218), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n232), .B(new_n233), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT66), .B(G50), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G222), .A2(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G223), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n247), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  OAI211_X1 g0053(.A(G1), .B(G13), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n251), .B(new_n255), .C1(G77), .C2(new_n247), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT67), .B(G45), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n260), .B2(G41), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G226), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n256), .A2(new_n261), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G200), .ZN(new_n267));
  INV_X1    g0067(.A(G190), .ZN(new_n268));
  INV_X1    g0068(.A(G13), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n269), .A2(new_n208), .A3(G1), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n216), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n208), .A2(G1), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(G50), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n269), .A2(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  OAI21_X1  g0078(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n279));
  INV_X1    g0079(.A(G150), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n208), .A2(new_n252), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G58), .ZN(new_n283));
  OR3_X1    g0083(.A1(new_n283), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT69), .B1(new_n283), .B2(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(KEYINPUT68), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT68), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G58), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT8), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n284), .B(new_n285), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n208), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n282), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n272), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n276), .B1(G50), .B2(new_n278), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n267), .B1(new_n268), .B2(new_n266), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT10), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n266), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n296), .B(new_n302), .C1(G179), .C2(new_n266), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n291), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n274), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(KEYINPUT76), .ZN(new_n307));
  INV_X1    g0107(.A(new_n273), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n306), .B2(KEYINPUT76), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n307), .A2(new_n309), .B1(new_n270), .B2(new_n305), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT68), .B(G58), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n202), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G159), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT72), .B1(new_n281), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G20), .A2(G33), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT72), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(G159), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n314), .A2(G20), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G33), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT7), .B1(new_n324), .B2(new_n208), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n208), .A2(KEYINPUT7), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n247), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(G68), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n320), .A2(new_n328), .A3(KEYINPUT16), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n272), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n324), .A2(new_n208), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT7), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n326), .B1(new_n334), .B2(KEYINPUT73), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n321), .A2(new_n323), .A3(new_n336), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n332), .A2(new_n333), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n320), .B1(new_n338), .B2(new_n313), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT16), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT74), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n335), .A2(new_n337), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n333), .B1(new_n247), .B2(G20), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n313), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n316), .A2(new_n319), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n201), .B1(new_n289), .B2(G68), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(new_n208), .ZN(new_n347));
  OAI211_X1 g0147(.A(KEYINPUT74), .B(new_n340), .C1(new_n344), .C2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n331), .B1(new_n341), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT75), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n340), .B1(new_n344), .B2(new_n347), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT74), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n348), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(KEYINPUT75), .A3(new_n331), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n311), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n261), .B1(new_n231), .B2(new_n263), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n249), .A2(G226), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n247), .B(new_n360), .C1(G223), .C2(G1698), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G87), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n254), .B1(new_n363), .B2(KEYINPUT77), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT77), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(new_n365), .A3(new_n362), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n359), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G179), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n301), .B2(new_n367), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT18), .B1(new_n358), .B2(new_n370), .ZN(new_n371));
  AOI211_X1 g0171(.A(new_n351), .B(new_n330), .C1(new_n355), .C2(new_n348), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT75), .B1(new_n356), .B2(new_n331), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n310), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT18), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(new_n369), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT17), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n367), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(G190), .B2(new_n367), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n358), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n310), .C1(new_n372), .C2(new_n373), .ZN(new_n382));
  XOR2_X1   g0182(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n371), .B(new_n376), .C1(new_n381), .C2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G238), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n261), .B1(new_n388), .B2(new_n263), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n231), .A2(G1698), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n247), .B(new_n390), .C1(G226), .C2(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G97), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n254), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT13), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n394), .A2(G190), .ZN(new_n395));
  INV_X1    g0195(.A(new_n393), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n264), .A2(G238), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n261), .A4(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n317), .A2(G50), .B1(G20), .B2(new_n313), .ZN(new_n400));
  INV_X1    g0200(.A(G77), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(new_n292), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n272), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT11), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT12), .B1(new_n278), .B2(G68), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT12), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n270), .A2(new_n407), .A3(new_n313), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n274), .A2(new_n313), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n406), .A2(new_n408), .B1(new_n273), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT71), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n402), .A2(KEYINPUT11), .A3(new_n272), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n405), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n405), .A2(new_n412), .A3(new_n410), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT71), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n395), .A2(new_n399), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT70), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n399), .A2(new_n394), .A3(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(KEYINPUT70), .B(KEYINPUT13), .C1(new_n389), .C2(new_n393), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n418), .A2(G200), .A3(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(G169), .A3(new_n419), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT14), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n418), .A2(new_n424), .A3(G169), .A4(new_n419), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n399), .A2(new_n394), .A3(G179), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n415), .A2(new_n413), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n421), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n247), .A2(G238), .A3(G1698), .ZN(new_n431));
  INV_X1    g0231(.A(G107), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n247), .A2(new_n249), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n431), .B1(new_n432), .B2(new_n247), .C1(new_n433), .C2(new_n231), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n255), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n264), .A2(G244), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n436), .A2(new_n261), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n301), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n273), .A2(G77), .A3(new_n275), .ZN(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT8), .B(G58), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n441), .A2(new_n281), .B1(new_n208), .B2(new_n401), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT15), .B(G87), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n442), .B1(new_n293), .B2(new_n444), .ZN(new_n445));
  OAI221_X1 g0245(.A(new_n440), .B1(G77), .B2(new_n278), .C1(new_n445), .C2(new_n295), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n438), .ZN(new_n448));
  INV_X1    g0248(.A(G179), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n446), .B1(new_n448), .B2(G190), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n438), .A2(G200), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n447), .A2(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n304), .A2(new_n387), .A3(new_n430), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n207), .B(G45), .C1(new_n253), .C2(KEYINPUT5), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT80), .B1(new_n458), .B2(new_n253), .ZN(new_n459));
  AND2_X1   g0259(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n460));
  NOR2_X1   g0260(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n461));
  OAI211_X1 g0261(.A(KEYINPUT80), .B(new_n253), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n457), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n254), .ZN(new_n465));
  INV_X1    g0265(.A(G257), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT81), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n321), .A2(new_n323), .A3(G250), .A4(G1698), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n321), .A2(new_n323), .A3(G244), .A4(new_n249), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT4), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n468), .B(new_n469), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n470), .A2(new_n471), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n255), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n253), .B1(new_n460), .B2(new_n461), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT80), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n456), .B1(new_n477), .B2(new_n462), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n255), .A2(new_n257), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n478), .A2(new_n255), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(G257), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n467), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G200), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT82), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n338), .A2(new_n432), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n432), .A2(KEYINPUT6), .A3(G97), .ZN(new_n490));
  INV_X1    g0290(.A(G97), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n432), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n204), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n490), .B1(new_n493), .B2(KEYINPUT6), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(G20), .B1(G77), .B2(new_n317), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n295), .B1(new_n489), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n270), .A2(new_n491), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n207), .A2(G33), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n273), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n499), .B2(new_n491), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n467), .A2(new_n481), .A3(new_n484), .A4(G190), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n485), .A2(KEYINPUT82), .A3(G200), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n488), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n501), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n485), .A2(G169), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n485), .A2(new_n449), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(G45), .ZN(new_n511));
  OAI21_X1  g0311(.A(G250), .B1(new_n511), .B2(G1), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n258), .A2(G45), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n255), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n247), .A2(G244), .A3(G1698), .ZN(new_n515));
  INV_X1    g0315(.A(G116), .ZN(new_n516));
  OAI221_X1 g0316(.A(new_n515), .B1(new_n252), .B2(new_n516), .C1(new_n433), .C2(new_n388), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n517), .B2(new_n255), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G190), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n247), .A2(new_n208), .A3(G68), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT19), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n208), .B1(new_n392), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(G87), .B2(new_n205), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n292), .B2(new_n491), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n525), .A2(new_n272), .B1(new_n270), .B2(new_n443), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n273), .A2(G87), .A3(new_n498), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n519), .B(new_n528), .C1(new_n378), .C2(new_n518), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n518), .A2(new_n449), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n526), .B1(new_n443), .B2(new_n499), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(new_n531), .C1(G169), .C2(new_n518), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n505), .A2(new_n510), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT83), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT83), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n505), .A2(new_n510), .A3(new_n537), .A4(new_n534), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT84), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n321), .A2(new_n323), .A3(G264), .A4(G1698), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n321), .A2(new_n323), .A3(G257), .A4(new_n249), .ZN(new_n541));
  INV_X1    g0341(.A(G303), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(new_n247), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n255), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n480), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(G270), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n478), .A2(new_n546), .A3(new_n255), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n539), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n478), .A2(new_n479), .B1(new_n543), .B2(new_n255), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n464), .A2(G270), .A3(new_n254), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT84), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n378), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT85), .B1(new_n499), .B2(new_n516), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT85), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n273), .A2(new_n554), .A3(G116), .A4(new_n498), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n468), .B(new_n208), .C1(G33), .C2(new_n491), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n516), .A2(G20), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n272), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT20), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  INV_X1    g0362(.A(new_n558), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n561), .A2(new_n562), .B1(new_n277), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n556), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT88), .B1(new_n552), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n551), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT84), .B1(new_n549), .B2(new_n550), .ZN(new_n568));
  OAI21_X1  g0368(.A(G200), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT88), .ZN(new_n570));
  INV_X1    g0370(.A(new_n565), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n548), .A2(G190), .A3(new_n551), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n566), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n321), .A2(new_n323), .A3(G257), .A4(G1698), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n321), .A2(new_n323), .A3(G250), .A4(new_n249), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G294), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n255), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n482), .B2(G264), .ZN(new_n581));
  AOI21_X1  g0381(.A(G169), .B1(new_n581), .B2(new_n480), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n464), .A2(G264), .A3(new_n254), .ZN(new_n583));
  AND4_X1   g0383(.A1(new_n449), .A2(new_n583), .A3(new_n480), .A4(new_n579), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n270), .A2(KEYINPUT25), .A3(new_n432), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT25), .B1(new_n270), .B2(new_n432), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n499), .A2(new_n432), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n321), .A2(new_n323), .A3(new_n208), .A4(G87), .ZN(new_n588));
  AND2_X1   g0388(.A1(KEYINPUT89), .A2(KEYINPUT22), .ZN(new_n589));
  NOR2_X1   g0389(.A1(KEYINPUT89), .A2(KEYINPUT22), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n247), .A2(new_n208), .A3(G87), .A4(new_n589), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT23), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n208), .B2(G107), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n432), .A2(KEYINPUT23), .A3(G20), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n252), .A2(new_n516), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n595), .A2(new_n596), .B1(new_n597), .B2(new_n208), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n592), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT24), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n592), .A2(new_n593), .A3(new_n598), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n587), .B1(new_n603), .B2(new_n272), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n582), .A2(new_n584), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n581), .A2(new_n480), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G200), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT90), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n583), .A2(G190), .A3(new_n480), .A4(new_n579), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .A4(new_n604), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(new_n609), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n378), .B1(new_n581), .B2(new_n480), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT90), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n605), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n301), .B1(new_n556), .B2(new_n564), .ZN(new_n615));
  OAI211_X1 g0415(.A(KEYINPUT21), .B(new_n615), .C1(new_n567), .C2(new_n568), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT86), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n548), .A2(new_n551), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT86), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(KEYINPUT21), .A4(new_n615), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n615), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n545), .A2(new_n547), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(G179), .A3(new_n565), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT87), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT87), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n624), .A2(new_n627), .A3(new_n565), .A4(G179), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n622), .A2(new_n623), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n574), .A2(new_n614), .A3(new_n621), .A4(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n455), .A2(new_n536), .A3(new_n538), .A4(new_n630), .ZN(G372));
  NAND2_X1  g0431(.A1(new_n382), .A2(KEYINPUT17), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n352), .A2(new_n357), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(new_n310), .A3(new_n380), .A4(new_n383), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n427), .A2(new_n429), .ZN(new_n636));
  INV_X1    g0436(.A(new_n421), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n450), .A2(new_n446), .A3(new_n439), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT92), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n447), .A2(KEYINPUT92), .A3(new_n450), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n635), .B1(new_n636), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n371), .A2(new_n376), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n300), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n303), .ZN(new_n646));
  INV_X1    g0446(.A(new_n605), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n629), .A2(new_n621), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n610), .A2(new_n613), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n505), .A2(new_n510), .A3(new_n650), .A4(new_n534), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n532), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n510), .A2(new_n653), .A3(new_n533), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n507), .B1(new_n449), .B2(new_n485), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT91), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n501), .B1(new_n655), .B2(new_n656), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(new_n534), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n654), .B1(new_n659), .B2(new_n653), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n646), .B1(new_n454), .B2(new_n661), .ZN(G369));
  NAND2_X1  g0462(.A1(new_n629), .A2(new_n621), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n277), .A2(new_n208), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT94), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n605), .A2(new_n669), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT93), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n614), .B1(new_n604), .B2(new_n670), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n605), .A2(new_n670), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n571), .A2(new_n670), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n663), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n681), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n574), .A2(new_n621), .A3(new_n629), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n685), .A2(new_n676), .A3(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n211), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n215), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(new_n690), .ZN(new_n694));
  XOR2_X1   g0494(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n695));
  XNOR2_X1  g0495(.A(new_n694), .B(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n670), .B1(new_n652), .B2(new_n660), .ZN(new_n697));
  XNOR2_X1  g0497(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n653), .B1(new_n510), .B2(new_n533), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT97), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT26), .A4(new_n534), .ZN(new_n703));
  OAI211_X1 g0503(.A(KEYINPUT97), .B(new_n653), .C1(new_n510), .C2(new_n533), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI211_X1 g0506(.A(KEYINPUT29), .B(new_n670), .C1(new_n706), .C2(new_n652), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G330), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n630), .A2(new_n536), .A3(new_n538), .A4(new_n670), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n624), .A2(G179), .A3(new_n518), .A4(new_n581), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  OR3_X1    g0512(.A1(new_n711), .A2(new_n712), .A3(new_n485), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n518), .A2(G179), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n618), .A2(new_n485), .A3(new_n606), .A4(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n712), .B1(new_n711), .B2(new_n485), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT31), .B1(new_n717), .B2(new_n669), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n709), .B1(new_n710), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n708), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n696), .B1(new_n722), .B2(G1), .ZN(G364));
  NOR2_X1   g0523(.A1(new_n269), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n207), .B1(new_n724), .B2(G45), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n689), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n685), .B2(G330), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G330), .B2(new_n685), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT98), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n211), .B(new_n247), .C1(new_n730), .C2(G355), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT98), .B1(new_n205), .B2(G87), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n731), .A2(new_n732), .B1(G116), .B2(new_n211), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n242), .A2(G45), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n688), .B(new_n247), .C1(new_n215), .C2(new_n259), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n216), .B1(G20), .B2(new_n301), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n727), .B1(new_n736), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n208), .A2(new_n449), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G190), .A3(G200), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT100), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n745), .A2(new_n746), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n268), .A2(G179), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n208), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n751), .A2(G326), .B1(G294), .B2(new_n754), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT101), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(KEYINPUT101), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n208), .A2(G179), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(new_n268), .A3(G200), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n758), .A2(new_n760), .B1(new_n761), .B2(new_n542), .ZN(new_n762));
  INV_X1    g0562(.A(new_n744), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n763), .A2(G190), .A3(new_n378), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT33), .B(G317), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G311), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G190), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n744), .A2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n763), .A2(new_n268), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G322), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n324), .B1(new_n767), .B2(new_n769), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n759), .A2(new_n768), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT102), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n773), .B1(G329), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n756), .A2(new_n757), .A3(new_n766), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n760), .A2(new_n432), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT32), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n774), .A2(new_n315), .ZN(new_n781));
  INV_X1    g0581(.A(new_n764), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n779), .B1(new_n780), .B2(new_n781), .C1(new_n782), .C2(new_n313), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G50), .B2(new_n751), .ZN(new_n784));
  INV_X1    g0584(.A(G87), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n761), .A2(new_n785), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n247), .B1(new_n769), .B2(new_n401), .C1(new_n753), .C2(new_n491), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(new_n780), .C2(new_n781), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n770), .B(KEYINPUT99), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n784), .B(new_n788), .C1(new_n312), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n777), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n743), .B1(new_n791), .B2(new_n740), .ZN(new_n792));
  INV_X1    g0592(.A(new_n739), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n685), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n729), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(G396));
  NAND2_X1  g0596(.A1(new_n638), .A2(KEYINPUT104), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT104), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n447), .A2(new_n798), .A3(new_n450), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n446), .A2(new_n669), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n451), .B2(new_n452), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n797), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(KEYINPUT105), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n640), .A2(new_n641), .A3(new_n800), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT105), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n797), .A2(new_n799), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n697), .B(new_n807), .Z(new_n808));
  INV_X1    g0608(.A(new_n721), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n727), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n809), .B2(new_n808), .ZN(new_n811));
  INV_X1    g0611(.A(new_n740), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n738), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n727), .B1(new_n813), .B2(G77), .ZN(new_n814));
  INV_X1    g0614(.A(G294), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n324), .B1(new_n771), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n769), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n816), .B1(G116), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n751), .A2(G303), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n753), .A2(new_n491), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n785), .A2(new_n760), .B1(new_n761), .B2(new_n432), .ZN(new_n821));
  XOR2_X1   g0621(.A(KEYINPUT103), .B(G283), .Z(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n820), .B(new_n821), .C1(new_n764), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n775), .A2(G311), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n818), .A2(new_n819), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n782), .A2(new_n280), .B1(new_n769), .B2(new_n315), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n750), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n789), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n827), .B(new_n829), .C1(G143), .C2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n831), .A2(KEYINPUT34), .ZN(new_n832));
  INV_X1    g0632(.A(new_n760), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n324), .B1(new_n833), .B2(G68), .ZN(new_n834));
  INV_X1    g0634(.A(G50), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n835), .B2(new_n761), .C1(new_n312), .C2(new_n753), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G132), .B2(new_n775), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n831), .B2(KEYINPUT34), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n826), .B1(new_n832), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n814), .B1(new_n839), .B2(new_n740), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n807), .B2(new_n738), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n811), .A2(new_n841), .ZN(G384));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n374), .A2(new_n369), .ZN(new_n844));
  INV_X1    g0644(.A(new_n667), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n374), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n844), .A2(new_n846), .A3(new_n847), .A4(new_n382), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT16), .B1(new_n320), .B2(new_n328), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n310), .B1(new_n330), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n369), .B2(new_n845), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n382), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n845), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI221_X4 g0655(.A(new_n843), .B1(new_n848), .B2(new_n853), .C1(new_n386), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n855), .B1(new_n635), .B2(new_n644), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n848), .A2(new_n853), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT38), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT39), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n857), .A2(KEYINPUT38), .A3(new_n858), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT39), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n358), .A2(new_n667), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n382), .B1(new_n358), .B2(new_n370), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n864), .B2(new_n863), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n386), .A2(new_n863), .B1(new_n865), .B2(new_n848), .ZN(new_n866));
  XNOR2_X1  g0666(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n861), .B(new_n862), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n860), .A2(KEYINPUT106), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n636), .A2(new_n669), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n371), .A2(new_n376), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n632), .A2(new_n634), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n854), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n848), .A2(new_n853), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n843), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n861), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT106), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT39), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n869), .A2(new_n870), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n428), .A2(new_n670), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n880), .B(new_n421), .C1(new_n427), .C2(new_n429), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n429), .B(new_n669), .C1(new_n427), .C2(new_n421), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n670), .B(new_n807), .C1(new_n652), .C2(new_n660), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n797), .A2(new_n799), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(new_n669), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n884), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n889), .A2(new_n876), .B1(new_n644), .B2(new_n667), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n879), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT108), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n879), .A2(KEYINPUT108), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n455), .A2(new_n707), .A3(new_n699), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n646), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT109), .Z(new_n898));
  XNOR2_X1  g0698(.A(new_n895), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n807), .B1(new_n881), .B2(new_n883), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n710), .B2(new_n720), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n876), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n386), .A2(new_n863), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n865), .A2(new_n848), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n867), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n901), .B(KEYINPUT40), .C1(new_n856), .C2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n454), .B1(new_n710), .B2(new_n720), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n909), .A2(new_n910), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n912), .A2(new_n709), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n899), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n899), .A2(new_n914), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n207), .B2(new_n724), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n915), .B1(new_n917), .B2(KEYINPUT110), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(KEYINPUT110), .B2(new_n917), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n494), .A2(KEYINPUT35), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n920), .A2(G116), .A3(new_n217), .A4(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT36), .ZN(new_n923));
  OAI21_X1  g0723(.A(G77), .B1(new_n312), .B2(new_n313), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n693), .A2(new_n924), .B1(G50), .B2(new_n313), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(G1), .A3(new_n269), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n919), .A2(new_n923), .A3(new_n926), .ZN(G367));
  INV_X1    g0727(.A(new_n727), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n688), .A2(new_n247), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n237), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n742), .B1(new_n688), .B2(new_n444), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n532), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n528), .A2(new_n670), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n533), .B2(new_n934), .ZN(new_n936));
  INV_X1    g0736(.A(G317), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n324), .B1(new_n774), .B2(new_n937), .C1(new_n822), .C2(new_n769), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n764), .A2(G294), .B1(G97), .B2(new_n833), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n432), .B2(new_n753), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n938), .B(new_n940), .C1(G303), .C2(new_n830), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT46), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n761), .B2(new_n516), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT114), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n751), .A2(G311), .B1(new_n944), .B2(new_n943), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n761), .A2(new_n942), .A3(new_n516), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT113), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n941), .A2(new_n945), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n754), .A2(G68), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n771), .B2(new_n280), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT115), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(KEYINPUT115), .ZN(new_n953));
  INV_X1    g0753(.A(G143), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n952), .B(new_n953), .C1(new_n954), .C2(new_n750), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT116), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n247), .B1(new_n774), .B2(new_n828), .C1(new_n835), .C2(new_n769), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n782), .A2(new_n315), .B1(new_n312), .B2(new_n761), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n958), .B(new_n959), .C1(G77), .C2(new_n833), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n955), .B2(new_n956), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n949), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  OAI221_X1 g0763(.A(new_n932), .B1(new_n793), .B2(new_n936), .C1(new_n963), .C2(new_n812), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT117), .ZN(new_n965));
  INV_X1    g0765(.A(new_n686), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n676), .B1(new_n685), .B2(G330), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(new_n672), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n672), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(KEYINPUT112), .A3(new_n722), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT112), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n708), .A2(new_n721), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n971), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT111), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n657), .A2(new_n658), .A3(new_n669), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n505), .B(new_n510), .C1(new_n501), .C2(new_n670), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n677), .A2(new_n678), .A3(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  INV_X1    g0785(.A(new_n981), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n679), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n679), .A2(KEYINPUT44), .A3(new_n986), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n984), .A2(new_n985), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n978), .B1(new_n991), .B2(new_n686), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n984), .A2(new_n985), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n989), .A2(new_n990), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(KEYINPUT111), .A3(new_n966), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n991), .A2(new_n686), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n977), .A2(new_n992), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n998), .A2(new_n722), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n689), .B(KEYINPUT41), .Z(new_n1000));
  OAI21_X1  g0800(.A(new_n725), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n672), .A2(new_n676), .A3(new_n981), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT42), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n981), .A2(new_n605), .B1(new_n506), .B2(new_n655), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n669), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1003), .A2(KEYINPUT42), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1002), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n966), .A2(new_n981), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1010), .B(new_n1011), .Z(new_n1012));
  AOI21_X1  g0812(.A(new_n965), .B1(new_n1001), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(G387));
  AOI21_X1  g0814(.A(new_n690), .B1(new_n973), .B2(new_n976), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT119), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1015), .A2(KEYINPUT119), .B1(new_n975), .B2(new_n971), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n972), .A2(new_n726), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n211), .A2(new_n247), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1020), .A2(new_n691), .B1(G107), .B2(new_n211), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n234), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n441), .A2(G50), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT50), .Z(new_n1024));
  OAI211_X1 g0824(.A(new_n691), .B(new_n511), .C1(new_n313), .C2(new_n401), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n929), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1022), .A2(new_n260), .B1(KEYINPUT118), .B2(new_n1026), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(KEYINPUT118), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1021), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n727), .B1(new_n1029), .B2(new_n742), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n771), .A2(new_n835), .B1(new_n769), .B2(new_n313), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n774), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n324), .B(new_n1031), .C1(G150), .C2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n401), .A2(new_n761), .B1(new_n760), .B2(new_n491), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n753), .A2(new_n443), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n751), .A2(G159), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n291), .A2(new_n764), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1033), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n247), .B1(new_n1032), .B2(G326), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n753), .A2(new_n822), .B1(new_n761), .B2(new_n815), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n764), .A2(G311), .B1(G303), .B2(new_n817), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n772), .B2(new_n750), .C1(new_n789), .C2(new_n937), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n1043), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT49), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1040), .B1(new_n516), .B2(new_n760), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1039), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1030), .B1(new_n1050), .B2(new_n740), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n676), .B2(new_n793), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1019), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1018), .A2(new_n1054), .ZN(G393));
  NAND2_X1  g0855(.A1(new_n995), .A2(new_n966), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n997), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n973), .A2(new_n976), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n690), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1059), .A2(new_n998), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n741), .B1(new_n491), .B2(new_n211), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n929), .B2(new_n245), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n750), .A2(new_n280), .B1(new_n315), .B2(new_n771), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT51), .Z(new_n1064));
  OAI22_X1  g0864(.A1(new_n782), .A2(new_n835), .B1(new_n760), .B2(new_n785), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n247), .B1(new_n774), .B2(new_n954), .C1(new_n441), .C2(new_n769), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n753), .A2(new_n401), .B1(new_n761), .B2(new_n313), .ZN(new_n1067));
  OR3_X1    g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n750), .A2(new_n937), .B1(new_n767), .B2(new_n771), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT52), .Z(new_n1070));
  INV_X1    g0870(.A(new_n761), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n823), .A2(new_n1071), .B1(new_n1032), .B2(G322), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT120), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n247), .B(new_n778), .C1(G294), .C2(new_n817), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(KEYINPUT120), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G303), .A2(new_n764), .B1(new_n754), .B2(G116), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1064), .A2(new_n1068), .B1(new_n1070), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n928), .B(new_n1062), .C1(new_n1078), .C2(new_n740), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n981), .B2(new_n793), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n1057), .B2(new_n725), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1060), .A2(new_n1081), .ZN(G390));
  OAI21_X1  g0882(.A(new_n727), .B1(new_n291), .B2(new_n813), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n761), .A2(new_n280), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n751), .B2(G128), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n782), .A2(new_n828), .B1(new_n315), .B2(new_n753), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G50), .B2(new_n833), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n775), .A2(G125), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT54), .B(G143), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n769), .A2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n324), .B(new_n1092), .C1(G132), .C2(new_n770), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n782), .A2(new_n432), .B1(new_n769), .B2(new_n491), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n751), .B2(G283), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT122), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n247), .B(new_n786), .C1(G116), .C2(new_n770), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n775), .A2(G294), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n754), .A2(G77), .B1(new_n833), .B2(G68), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1094), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1083), .B1(new_n1102), .B2(new_n740), .ZN(new_n1103));
  AOI211_X1 g0903(.A(KEYINPUT106), .B(new_n862), .C1(new_n875), .C2(new_n861), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n877), .B1(new_n876), .B2(KEYINPUT39), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n868), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1103), .B1(new_n1106), .B2(new_n738), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n721), .B(new_n807), .C1(new_n881), .C2(new_n883), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n670), .B(new_n807), .C1(new_n706), .C2(new_n652), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n884), .B1(new_n1109), .B2(new_n888), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n856), .A2(new_n907), .ZN(new_n1111));
  OR3_X1    g0911(.A1(new_n1110), .A2(new_n870), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n889), .A2(new_n870), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1108), .B(new_n1112), .C1(new_n1106), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1108), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1113), .B1(new_n869), .B2(new_n878), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1110), .A2(new_n1111), .A3(new_n870), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1107), .B1(new_n1119), .B2(new_n725), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n896), .B(new_n646), .C1(new_n454), .C2(new_n809), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n721), .A2(new_n807), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n884), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1108), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n885), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n887), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1123), .A2(new_n888), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1121), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1114), .A2(new_n1118), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1128), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n690), .B1(new_n1119), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1120), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(G378));
  INV_X1    g0933(.A(KEYINPUT57), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1121), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n710), .A2(new_n720), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n880), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n430), .A2(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n806), .A2(new_n804), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1139), .A2(new_n882), .B1(new_n1140), .B2(new_n803), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n861), .B2(new_n875), .ZN(new_n1143));
  OAI211_X1 g0943(.A(G330), .B(new_n908), .C1(new_n1143), .C2(KEYINPUT40), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n296), .A2(new_n845), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n304), .A2(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n300), .A2(new_n303), .A3(new_n1145), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OR3_X1    g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1149), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1144), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n904), .A2(G330), .A3(new_n908), .A4(new_n1152), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(new_n893), .A3(new_n894), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n879), .A2(KEYINPUT108), .A3(new_n890), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT108), .B1(new_n879), .B2(new_n890), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1134), .B1(new_n1136), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1164), .A2(KEYINPUT57), .A3(new_n1157), .A4(new_n1161), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n689), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1162), .A2(new_n725), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n727), .B1(new_n813), .B2(G50), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n770), .A2(G107), .B1(new_n444), .B2(new_n817), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n764), .A2(G97), .B1(new_n289), .B2(new_n833), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n1170), .A3(new_n950), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G283), .B2(new_n775), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n253), .B(new_n324), .C1(new_n761), .C2(new_n401), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT123), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(new_n516), .C2(new_n750), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT58), .ZN(new_n1176));
  AOI21_X1  g0976(.A(G50), .B1(new_n252), .B2(new_n253), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n247), .B2(G41), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n751), .A2(G125), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n764), .A2(G132), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n770), .A2(G128), .B1(G137), .B2(new_n817), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1091), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n754), .A2(G150), .B1(new_n1071), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n833), .A2(G159), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G33), .B(G41), .C1(new_n1032), .C2(G124), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1176), .B(new_n1178), .C1(new_n1185), .C2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1168), .B1(new_n1190), .B2(new_n740), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1152), .B2(new_n738), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT124), .Z(new_n1193));
  NOR2_X1   g0993(.A1(new_n1167), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1166), .A2(new_n1194), .ZN(G375));
  NAND2_X1  g0995(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1121), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1000), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n1199), .A3(new_n1130), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n727), .B1(new_n813), .B2(G68), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n754), .A2(G50), .B1(new_n1071), .B2(G159), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n782), .B2(new_n1091), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G132), .B2(new_n751), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n247), .B1(new_n769), .B2(new_n280), .C1(new_n312), .C2(new_n760), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G128), .B2(new_n775), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n828), .C2(new_n789), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n753), .A2(new_n443), .B1(new_n760), .B2(new_n401), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n324), .B1(new_n432), .B2(new_n769), .C1(new_n771), .C2(new_n758), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(G116), .C2(new_n764), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n815), .B2(new_n750), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n775), .A2(G303), .B1(G97), .B2(new_n1071), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT125), .Z(new_n1213));
  OAI21_X1  g1013(.A(new_n1207), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1201), .B1(new_n1214), .B2(new_n740), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n884), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n738), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1197), .B2(new_n725), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1200), .A2(new_n1219), .ZN(G381));
  NAND3_X1  g1020(.A1(new_n1018), .A2(new_n795), .A3(new_n1054), .ZN(new_n1221));
  OR4_X1    g1021(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1166), .A2(new_n1132), .A3(new_n1194), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n1222), .A2(G387), .A3(new_n1223), .ZN(G407));
  NAND2_X1  g1024(.A1(new_n668), .A2(G213), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT126), .Z(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(new_n1223), .C2(new_n1227), .ZN(G409));
  INV_X1    g1028(.A(KEYINPUT61), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1166), .A2(G378), .A3(new_n1194), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1157), .A2(new_n1161), .A3(KEYINPUT127), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT127), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n725), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1164), .A2(new_n1199), .A3(new_n1157), .A4(new_n1161), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1192), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1132), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1226), .B1(new_n1230), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT60), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1198), .B1(new_n1238), .B2(new_n1128), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1196), .A2(new_n1135), .A3(new_n1238), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(new_n690), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1218), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(G384), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1242), .A2(G384), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G2897), .B(new_n1226), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1245), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1226), .A2(G2897), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1243), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1229), .B1(new_n1237), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT63), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1230), .A2(new_n1236), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1227), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1253), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G393), .A2(G396), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(G390), .A2(new_n1259), .A3(new_n1221), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1060), .A2(new_n1081), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n795), .B1(new_n1018), .B2(new_n1054), .ZN(new_n1262));
  AOI211_X1 g1062(.A(G396), .B(new_n1053), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1260), .A2(new_n1013), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1013), .B1(new_n1260), .B2(new_n1264), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1237), .A2(KEYINPUT63), .A3(new_n1256), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1252), .A2(new_n1258), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1237), .A2(new_n1270), .A3(new_n1256), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1237), .B2(new_n1256), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1271), .A2(new_n1251), .A3(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1269), .B1(new_n1273), .B2(new_n1267), .ZN(G405));
  AOI21_X1  g1074(.A(G378), .B1(new_n1166), .B2(new_n1194), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1276), .A2(new_n1257), .A3(new_n1230), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1257), .B1(new_n1276), .B2(new_n1230), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(new_n1267), .ZN(G402));
endmodule


