//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT89), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT13), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT16), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(G1gat), .B2(new_n205), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(G8gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n212), .A2(new_n217), .A3(G29gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(G36gat), .B1(new_n214), .B2(new_n215), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT15), .B1(new_n223), .B2(new_n220), .ZN(new_n224));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n225), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n227), .B(KEYINPUT15), .C1(new_n223), .C2(new_n220), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n211), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n210), .A2(new_n229), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n204), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n226), .A2(KEYINPUT17), .A3(new_n228), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT88), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n226), .A2(KEYINPUT88), .A3(new_n228), .A4(KEYINPUT17), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n210), .B1(new_n229), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n203), .A3(new_n232), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n233), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(G197gat), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT11), .B(G169gat), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n241), .A2(KEYINPUT18), .A3(new_n203), .A4(new_n232), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n244), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n249), .B1(new_n244), .B2(new_n250), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT32), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT27), .B(G183gat), .ZN(new_n255));
  INV_X1    g054(.A(G190gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(KEYINPUT28), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT27), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OR2_X1    g059(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n261));
  AOI21_X1  g060(.A(G190gat), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n257), .B1(new_n262), .B2(KEYINPUT28), .ZN(new_n263));
  NAND2_X1  g062(.A1(G183gat), .A2(G190gat), .ZN(new_n264));
  OR2_X1    g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT26), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n265), .A2(new_n266), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n272));
  INV_X1    g071(.A(KEYINPUT23), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(G176gat), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT65), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G169gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n268), .A2(KEYINPUT23), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n265), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n264), .A2(KEYINPUT24), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT24), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(G183gat), .A3(G190gat), .ZN(new_n285));
  INV_X1    g084(.A(G183gat), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n283), .A2(new_n285), .B1(new_n286), .B2(new_n256), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n272), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n283), .A2(new_n285), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n286), .ZN(new_n291));
  NAND2_X1  g090(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n256), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n291), .A2(new_n295), .A3(new_n256), .A4(new_n292), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n289), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n274), .A2(new_n275), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n298), .A3(KEYINPUT25), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n288), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G113gat), .B(G120gat), .Z(new_n301));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n303));
  XNOR2_X1  g102(.A(G127gat), .B(G134gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n301), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(G127gat), .B(G134gat), .Z(new_n306));
  NAND2_X1  g105(.A1(new_n303), .A2(new_n302), .ZN(new_n307));
  XNOR2_X1  g106(.A(G113gat), .B(G120gat), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n306), .B(new_n307), .C1(KEYINPUT1), .C2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n271), .A2(new_n300), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT69), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n271), .A2(new_n300), .A3(new_n313), .A4(new_n310), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n271), .A2(new_n300), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n305), .A2(new_n309), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n312), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(G227gat), .A2(G233gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n254), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT33), .ZN(new_n321));
  XNOR2_X1  g120(.A(G15gat), .B(G43gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(G71gat), .B(G99gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n320), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT33), .B1(new_n318), .B2(new_n319), .ZN(new_n326));
  NOR4_X1   g125(.A1(new_n320), .A2(new_n326), .A3(KEYINPUT70), .A4(new_n324), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT70), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n318), .A2(new_n319), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n324), .B1(new_n329), .B2(KEYINPUT32), .ZN(new_n330));
  INV_X1    g129(.A(new_n326), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n325), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n318), .A2(new_n319), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n336), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n338), .B(new_n325), .C1(new_n327), .C2(new_n332), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT36), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(KEYINPUT72), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n333), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(KEYINPUT36), .A3(new_n339), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G228gat), .ZN(new_n348));
  INV_X1    g147(.A(G233gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G141gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G148gat), .ZN(new_n352));
  INV_X1    g151(.A(G148gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G141gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n352), .A2(new_n354), .B1(KEYINPUT2), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  NOR2_X1   g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT78), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G155gat), .ZN(new_n360));
  INV_X1    g159(.A(G162gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(new_n355), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n355), .ZN(new_n366));
  XNOR2_X1  g165(.A(G141gat), .B(G148gat), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n355), .A2(KEYINPUT2), .ZN(new_n368));
  OAI211_X1 g167(.A(KEYINPUT78), .B(new_n366), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372));
  XNOR2_X1  g171(.A(G211gat), .B(G218gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G211gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT73), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT73), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G211gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT22), .B1(new_n379), .B2(G218gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(G197gat), .B(G204gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n374), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G218gat), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n376), .B2(new_n378), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n381), .B(new_n373), .C1(new_n385), .C2(KEYINPUT22), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n372), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI211_X1 g188(.A(KEYINPUT82), .B(KEYINPUT29), .C1(new_n383), .C2(new_n386), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n371), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n383), .A2(new_n386), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n370), .A2(new_n372), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n350), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n386), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT22), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT73), .B(G211gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(new_n384), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n373), .B1(new_n401), .B2(new_n381), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n393), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n370), .B1(new_n403), .B2(new_n372), .ZN(new_n404));
  INV_X1    g203(.A(new_n350), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n404), .A2(new_n395), .A3(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(KEYINPUT84), .B(G22gat), .C1(new_n397), .C2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408));
  INV_X1    g207(.A(G50gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n410), .B(new_n411), .Z(new_n412));
  INV_X1    g211(.A(new_n406), .ZN(new_n413));
  INV_X1    g212(.A(G22gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n403), .A2(KEYINPUT82), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n387), .A2(new_n388), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n416), .A3(new_n372), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n395), .B1(new_n417), .B2(new_n371), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n413), .B(new_n414), .C1(new_n418), .C2(new_n350), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n407), .A2(new_n412), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT3), .B1(new_n403), .B2(KEYINPUT82), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n370), .B1(new_n421), .B2(new_n416), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n405), .B1(new_n422), .B2(new_n395), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n413), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT84), .B1(new_n424), .B2(G22gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n423), .A2(new_n427), .A3(new_n414), .A4(new_n413), .ZN(new_n428));
  INV_X1    g227(.A(new_n412), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(G22gat), .B1(new_n397), .B2(new_n406), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(new_n419), .A3(KEYINPUT83), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n420), .A2(new_n426), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n365), .A2(new_n369), .A3(KEYINPUT3), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n394), .A2(new_n316), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G225gat), .A2(G233gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(KEYINPUT5), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n370), .A2(new_n305), .A3(new_n309), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT4), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n310), .A2(new_n441), .A3(new_n370), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n440), .A2(KEYINPUT80), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT80), .B1(new_n440), .B2(new_n442), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n435), .B(new_n438), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n371), .A2(new_n316), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n439), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n448), .B2(new_n437), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n440), .A2(KEYINPUT79), .A3(new_n442), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT79), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n439), .A2(new_n451), .A3(KEYINPUT4), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(new_n436), .A3(new_n435), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n449), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n445), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G1gat), .B(G29gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT0), .ZN(new_n457));
  XNOR2_X1  g256(.A(G57gat), .B(G85gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n459), .A3(new_n454), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n455), .A2(KEYINPUT6), .A3(new_n460), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n392), .ZN(new_n467));
  NAND2_X1  g266(.A1(G226gat), .A2(G233gat), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n468), .B(KEYINPUT74), .Z(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n470), .B1(new_n315), .B2(new_n393), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n469), .B1(new_n271), .B2(new_n300), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G8gat), .B(G36gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT75), .ZN(new_n475));
  XNOR2_X1  g274(.A(G64gat), .B(G92gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n315), .A2(new_n470), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT29), .B1(new_n271), .B2(new_n300), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n478), .B(new_n392), .C1(new_n479), .C2(new_n470), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n473), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT76), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n473), .A2(KEYINPUT76), .A3(new_n480), .A4(new_n477), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT77), .B(KEYINPUT30), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n477), .B1(new_n473), .B2(new_n480), .ZN(new_n487));
  INV_X1    g286(.A(new_n481), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(KEYINPUT30), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n433), .B1(new_n466), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n431), .A2(KEYINPUT83), .A3(new_n419), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n428), .A2(new_n429), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n407), .A2(new_n412), .A3(new_n419), .ZN(new_n494));
  OAI22_X1  g293(.A1(new_n492), .A2(new_n493), .B1(new_n494), .B2(new_n425), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n435), .B1(new_n443), .B2(new_n444), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n437), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(KEYINPUT39), .C1(new_n437), .C2(new_n448), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n498), .B(new_n459), .C1(KEYINPUT39), .C2(new_n497), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT40), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n500), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n461), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n486), .A2(new_n489), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n495), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n466), .A2(new_n483), .A3(new_n484), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n473), .A2(new_n480), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n477), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT38), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n507), .A2(new_n508), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n511), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n511), .B1(new_n509), .B2(new_n513), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n506), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n347), .B(new_n491), .C1(new_n505), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n464), .A2(new_n465), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n486), .A4(new_n489), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(new_n433), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n521), .A2(KEYINPUT86), .A3(new_n339), .A4(new_n337), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT86), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n495), .A2(new_n519), .A3(new_n518), .A4(new_n504), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n523), .B1(new_n340), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n466), .A2(new_n490), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n345), .A2(new_n527), .A3(new_n339), .A4(new_n495), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n253), .B1(new_n517), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G64gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G57gat), .ZN(new_n533));
  INV_X1    g332(.A(G57gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G64gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT9), .ZN(new_n536));
  NAND2_X1  g335(.A1(G71gat), .A2(G78gat), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n533), .A2(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(G71gat), .A2(G78gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n537), .B(KEYINPUT90), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(KEYINPUT9), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n537), .ZN(new_n545));
  INV_X1    g344(.A(new_n533), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT91), .B(G57gat), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(G64gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n534), .A2(KEYINPUT91), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G57gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n553), .A3(G64gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n533), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(KEYINPUT92), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n543), .B1(new_n550), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G127gat), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n541), .A2(new_n538), .A3(new_n539), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n555), .A2(KEYINPUT92), .B1(new_n537), .B2(new_n544), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n557), .A2(KEYINPUT94), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT21), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n211), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n562), .A2(new_n571), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(new_n360), .ZN(new_n576));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n572), .A2(new_n573), .A3(new_n578), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT41), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT95), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT96), .ZN(new_n587));
  XOR2_X1   g386(.A(G134gat), .B(G162gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G99gat), .B(G106gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT7), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(KEYINPUT97), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT8), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n594), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT7), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(KEYINPUT97), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n602), .A2(new_n603), .A3(G85gat), .A4(G92gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n591), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g404(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n595), .B2(new_n596), .ZN(new_n606));
  AND4_X1   g405(.A1(new_n591), .A2(new_n604), .A3(new_n594), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n608), .B1(new_n229), .B2(new_n239), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n238), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G190gat), .B(G218gat), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n600), .A2(new_n604), .ZN(new_n612));
  INV_X1    g411(.A(new_n591), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n600), .A2(new_n591), .A3(new_n604), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI22_X1  g415(.A1(new_n230), .A2(new_n616), .B1(new_n584), .B2(new_n583), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n610), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n617), .B1(new_n609), .B2(new_n238), .ZN(new_n619));
  INV_X1    g418(.A(new_n611), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n590), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n611), .B1(new_n610), .B2(new_n617), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n620), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n624), .A3(new_n589), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n613), .A2(KEYINPUT98), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n616), .B1(new_n557), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n566), .A2(new_n608), .A3(new_n628), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT10), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n616), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n568), .A3(new_n569), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G230gat), .A2(G233gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT99), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n639), .B1(new_n630), .B2(new_n631), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  NAND3_X1  g444(.A1(new_n640), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n638), .B1(new_n633), .B2(new_n635), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(new_n641), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n646), .A2(KEYINPUT100), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT100), .B1(new_n646), .B2(new_n649), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n582), .A2(new_n627), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n531), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n518), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT101), .B(G1gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1324gat));
  NOR2_X1   g457(.A1(new_n655), .A2(new_n504), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(G8gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n662), .B2(new_n659), .ZN(new_n663));
  MUX2_X1   g462(.A(new_n661), .B(new_n663), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g463(.A(G15gat), .B1(new_n655), .B2(new_n347), .ZN(new_n665));
  INV_X1    g464(.A(new_n340), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n531), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n653), .A2(G15gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(G1326gat));
  NOR2_X1   g468(.A1(new_n655), .A2(new_n495), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673));
  AOI221_X4 g472(.A(new_n673), .B1(new_n528), .B2(KEYINPUT35), .C1(new_n522), .C2(new_n525), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT102), .B1(new_n526), .B2(new_n529), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n517), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT103), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n517), .B(new_n678), .C1(new_n674), .C2(new_n675), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n627), .A2(KEYINPUT44), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n627), .B1(new_n517), .B2(new_n530), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n652), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n582), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n253), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n518), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n682), .A2(new_n689), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(G29gat), .A3(new_n518), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT45), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(G1328gat));
  NOR3_X1   g494(.A1(new_n692), .A2(G36gat), .A3(new_n504), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT46), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n690), .A2(new_n504), .ZN(new_n698));
  OAI21_X1  g497(.A(G36gat), .B1(new_n698), .B2(KEYINPUT104), .ZN(new_n699));
  INV_X1    g498(.A(new_n689), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n681), .B2(new_n684), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n701), .A2(KEYINPUT104), .A3(new_n490), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n697), .B1(new_n699), .B2(new_n702), .ZN(G1329gat));
  INV_X1    g502(.A(G43gat), .ZN(new_n704));
  INV_X1    g503(.A(new_n347), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n701), .B2(new_n705), .ZN(new_n706));
  NOR4_X1   g505(.A1(new_n667), .A2(G43gat), .A3(new_n627), .A4(new_n688), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(KEYINPUT105), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(KEYINPUT47), .ZN(new_n709));
  OR3_X1    g508(.A1(new_n706), .A2(new_n709), .A3(new_n707), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n706), .B2(new_n707), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1330gat));
  NOR3_X1   g511(.A1(new_n692), .A2(G50gat), .A3(new_n495), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n495), .B(new_n700), .C1(new_n681), .C2(new_n684), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  OAI21_X1  g516(.A(G50gat), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n701), .A2(new_n717), .A3(new_n433), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n715), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n716), .A2(new_n409), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n714), .B1(new_n721), .B2(new_n713), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(G1331gat));
  AND2_X1   g522(.A1(new_n677), .A2(new_n679), .ZN(new_n724));
  INV_X1    g523(.A(new_n582), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n686), .A2(new_n253), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n725), .A2(new_n626), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n518), .B(KEYINPUT107), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(new_n547), .ZN(G1332gat));
  NAND3_X1  g530(.A1(new_n724), .A2(new_n490), .A3(new_n727), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT49), .B(G64gat), .Z(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT108), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n733), .B(new_n737), .C1(new_n732), .C2(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1333gat));
  OAI21_X1  g538(.A(G71gat), .B1(new_n728), .B2(new_n347), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n340), .A2(G71gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n728), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n740), .B(KEYINPUT50), .C1(new_n728), .C2(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1334gat));
  NOR2_X1   g545(.A1(new_n728), .A2(new_n495), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT109), .B(G78gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1335gat));
  NOR2_X1   g548(.A1(new_n582), .A2(new_n726), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n681), .B2(new_n684), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G85gat), .B1(new_n753), .B2(new_n518), .ZN(new_n754));
  INV_X1    g553(.A(new_n253), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n582), .A2(new_n755), .A3(new_n627), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n676), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n676), .A2(KEYINPUT51), .A3(new_n756), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n652), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n595), .A3(new_n466), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n754), .A2(new_n762), .ZN(G1336gat));
  AOI21_X1  g562(.A(new_n596), .B1(new_n752), .B2(new_n490), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n596), .A3(new_n490), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n767), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT52), .B1(new_n769), .B2(new_n764), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1337gat));
  OAI21_X1  g570(.A(G99gat), .B1(new_n753), .B2(new_n347), .ZN(new_n772));
  INV_X1    g571(.A(G99gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n761), .A2(new_n773), .A3(new_n666), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1338gat));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(KEYINPUT53), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n760), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n495), .A2(G106gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n686), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(KEYINPUT53), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT110), .B(G106gat), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n752), .B2(new_n433), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n777), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n761), .A2(new_n779), .B1(new_n776), .B2(KEYINPUT53), .ZN(new_n786));
  INV_X1    g585(.A(new_n777), .ZN(new_n787));
  AOI211_X1 g586(.A(new_n495), .B(new_n751), .C1(new_n681), .C2(new_n684), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n786), .B(new_n787), .C1(new_n788), .C2(new_n783), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n785), .A2(new_n789), .ZN(G1339gat));
  NAND4_X1  g589(.A1(new_n582), .A2(new_n253), .A3(new_n627), .A4(new_n652), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n633), .A2(new_n638), .A3(new_n635), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n640), .A2(KEYINPUT54), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n645), .B1(new_n648), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n793), .A2(KEYINPUT55), .A3(new_n795), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n626), .A2(new_n798), .A3(new_n646), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n231), .A2(new_n232), .A3(new_n204), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n241), .A2(new_n232), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n203), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n248), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n244), .A2(new_n249), .A3(new_n250), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n800), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n805), .B(new_n804), .C1(new_n650), .C2(new_n651), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n646), .B(new_n799), .C1(new_n251), .C2(new_n252), .ZN(new_n809));
  INV_X1    g608(.A(new_n798), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n807), .B1(new_n811), .B2(new_n627), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n791), .B1(new_n812), .B2(new_n582), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n814), .A2(new_n340), .A3(new_n433), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n518), .A2(new_n490), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(G113gat), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n817), .A2(new_n818), .A3(new_n253), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n814), .A2(new_n729), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n345), .A2(new_n339), .A3(new_n495), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n490), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n755), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n819), .B1(new_n825), .B2(new_n818), .ZN(G1340gat));
  INV_X1    g625(.A(G120gat), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n817), .A2(new_n827), .A3(new_n652), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n686), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(new_n827), .ZN(G1341gat));
  INV_X1    g629(.A(G127gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n824), .A2(new_n831), .A3(new_n582), .ZN(new_n832));
  OAI21_X1  g631(.A(G127gat), .B1(new_n817), .B2(new_n725), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n504), .A2(new_n626), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT112), .ZN(new_n836));
  OR3_X1    g635(.A1(new_n823), .A2(G134gat), .A3(new_n836), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n838));
  OAI21_X1  g637(.A(G134gat), .B1(new_n817), .B2(new_n627), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G1343gat));
  AND2_X1   g640(.A1(new_n347), .A2(new_n816), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n433), .A2(KEYINPUT57), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n633), .A2(new_n638), .A3(new_n635), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(new_n648), .A3(new_n794), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n636), .A2(new_n794), .A3(new_n639), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n647), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT113), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n793), .A2(new_n849), .A3(new_n795), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n797), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT114), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n799), .A2(new_n646), .ZN(new_n853));
  INV_X1    g652(.A(new_n252), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n805), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n848), .A2(new_n856), .A3(new_n797), .A4(new_n850), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n852), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n626), .B1(new_n858), .B2(new_n808), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n725), .B1(new_n859), .B2(new_n807), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n843), .B1(new_n860), .B2(new_n791), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n813), .B2(new_n433), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n842), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(G141gat), .B1(new_n863), .B2(new_n253), .ZN(new_n864));
  XOR2_X1   g663(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n865));
  NAND3_X1  g664(.A1(new_n820), .A2(new_n347), .A3(new_n433), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n490), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n755), .A2(new_n351), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n864), .B(new_n865), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n863), .A2(KEYINPUT115), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n873), .B(new_n842), .C1(new_n861), .C2(new_n862), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n755), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n871), .B1(new_n876), .B2(G141gat), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n870), .B1(new_n877), .B2(new_n878), .ZN(G1344gat));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880));
  XNOR2_X1  g679(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n495), .A2(KEYINPUT57), .ZN(new_n883));
  INV_X1    g682(.A(new_n859), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n800), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n800), .A2(new_n885), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n886), .A2(new_n805), .A3(new_n804), .A4(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n582), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n791), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT57), .B1(new_n814), .B2(new_n495), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n686), .A4(new_n842), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n882), .B1(new_n893), .B2(G148gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n872), .A2(new_n686), .A3(new_n874), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n353), .A2(KEYINPUT59), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT117), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n899), .A3(new_n896), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n894), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n867), .A2(new_n353), .A3(new_n686), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n880), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n895), .A2(new_n899), .A3(new_n896), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n899), .B1(new_n895), .B2(new_n896), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT120), .B(new_n902), .C1(new_n907), .C2(new_n894), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n904), .A2(new_n908), .ZN(G1345gat));
  AOI21_X1  g708(.A(G155gat), .B1(new_n867), .B2(new_n582), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n582), .A2(G155gat), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT121), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n910), .B1(new_n875), .B2(new_n912), .ZN(G1346gat));
  AOI21_X1  g712(.A(new_n361), .B1(new_n875), .B2(new_n626), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n866), .A2(G162gat), .A3(new_n836), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n914), .A2(new_n915), .ZN(G1347gat));
  INV_X1    g715(.A(new_n729), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n504), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n815), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n253), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n814), .A2(new_n466), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n490), .A3(new_n822), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n755), .A2(new_n276), .A3(new_n278), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1348gat));
  INV_X1    g723(.A(new_n922), .ZN(new_n925));
  AOI21_X1  g724(.A(G176gat), .B1(new_n925), .B2(new_n686), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n815), .A2(G176gat), .A3(new_n686), .A4(new_n918), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n926), .A2(new_n929), .A3(new_n930), .ZN(G1349gat));
  NAND3_X1  g730(.A1(new_n925), .A2(new_n255), .A3(new_n582), .ZN(new_n932));
  OAI22_X1  g731(.A1(new_n919), .A2(new_n725), .B1(new_n259), .B2(new_n258), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n932), .A2(new_n933), .B1(KEYINPUT123), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(KEYINPUT123), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n935), .B(new_n936), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n919), .B2(new_n627), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT61), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n925), .A2(new_n256), .A3(new_n626), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1351gat));
  NOR3_X1   g740(.A1(new_n705), .A2(new_n504), .A3(new_n495), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n921), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(G197gat), .A3(new_n253), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT124), .Z(new_n945));
  AND4_X1   g744(.A1(new_n347), .A2(new_n891), .A3(new_n892), .A4(new_n918), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n755), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G197gat), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(new_n948), .ZN(G1352gat));
  INV_X1    g748(.A(new_n943), .ZN(new_n950));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n951), .A3(new_n686), .ZN(new_n952));
  XNOR2_X1  g751(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n951), .B1(new_n946), .B2(new_n686), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n956), .B(new_n957), .ZN(G1353gat));
  NAND3_X1  g757(.A1(new_n950), .A2(new_n400), .A3(new_n582), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n946), .A2(new_n582), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  OAI21_X1  g762(.A(new_n384), .B1(new_n943), .B2(new_n627), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT127), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n627), .A2(new_n384), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n946), .B2(new_n966), .ZN(G1355gat));
endmodule


