

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  BUF_X1 U322 ( .A(n500), .Z(n290) );
  XNOR2_X1 U323 ( .A(n422), .B(n421), .ZN(n524) );
  XNOR2_X1 U324 ( .A(n416), .B(KEYINPUT41), .ZN(n556) );
  XNOR2_X1 U325 ( .A(n456), .B(n455), .ZN(n525) );
  INV_X1 U326 ( .A(G92GAT), .ZN(n379) );
  XNOR2_X1 U327 ( .A(n380), .B(n379), .ZN(n381) );
  INV_X1 U328 ( .A(KEYINPUT48), .ZN(n421) );
  XNOR2_X1 U329 ( .A(n382), .B(n381), .ZN(n383) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n458) );
  XOR2_X1 U331 ( .A(n469), .B(KEYINPUT28), .Z(n527) );
  XNOR2_X1 U332 ( .A(n458), .B(KEYINPUT58), .ZN(n459) );
  XNOR2_X1 U333 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G92GAT), .B(G218GAT), .Z(n292) );
  XNOR2_X1 U335 ( .A(G36GAT), .B(G190GAT), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n292), .B(n291), .ZN(n428) );
  XOR2_X1 U337 ( .A(G99GAT), .B(G106GAT), .Z(n367) );
  XOR2_X1 U338 ( .A(G29GAT), .B(G85GAT), .Z(n334) );
  XOR2_X1 U339 ( .A(n367), .B(n334), .Z(n294) );
  XOR2_X1 U340 ( .A(G43GAT), .B(G134GAT), .Z(n445) );
  XOR2_X1 U341 ( .A(G50GAT), .B(G162GAT), .Z(n315) );
  XNOR2_X1 U342 ( .A(n445), .B(n315), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U344 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n296) );
  NAND2_X1 U345 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n303) );
  XOR2_X1 U348 ( .A(KEYINPUT75), .B(KEYINPUT64), .Z(n300) );
  XNOR2_X1 U349 ( .A(KEYINPUT66), .B(KEYINPUT74), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U351 ( .A(n301), .B(KEYINPUT10), .Z(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n428), .B(n304), .ZN(n307) );
  XOR2_X1 U354 ( .A(KEYINPUT69), .B(KEYINPUT8), .Z(n305) );
  XNOR2_X1 U355 ( .A(n305), .B(KEYINPUT7), .ZN(n358) );
  INV_X1 U356 ( .A(n358), .ZN(n306) );
  XOR2_X1 U357 ( .A(n307), .B(n306), .Z(n546) );
  XOR2_X1 U358 ( .A(KEYINPUT76), .B(n546), .Z(n476) );
  XOR2_X1 U359 ( .A(KEYINPUT89), .B(KEYINPUT92), .Z(n309) );
  XNOR2_X1 U360 ( .A(G148GAT), .B(KEYINPUT24), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U362 ( .A(n310), .B(G106GAT), .Z(n312) );
  XOR2_X1 U363 ( .A(KEYINPUT71), .B(G78GAT), .Z(n368) );
  XNOR2_X1 U364 ( .A(n368), .B(G218GAT), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n319) );
  XOR2_X1 U366 ( .A(G155GAT), .B(KEYINPUT3), .Z(n314) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n340) );
  XOR2_X1 U369 ( .A(n315), .B(n340), .Z(n317) );
  NAND2_X1 U370 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U372 ( .A(n319), .B(n318), .Z(n327) );
  XOR2_X1 U373 ( .A(KEYINPUT21), .B(G211GAT), .Z(n321) );
  XNOR2_X1 U374 ( .A(KEYINPUT90), .B(G204GAT), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U376 ( .A(G197GAT), .B(n322), .Z(n429) );
  XOR2_X1 U377 ( .A(KEYINPUT91), .B(KEYINPUT22), .Z(n324) );
  XNOR2_X1 U378 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n429), .B(n325), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n469) );
  XOR2_X1 U382 ( .A(KEYINPUT95), .B(KEYINPUT6), .Z(n329) );
  XNOR2_X1 U383 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U385 ( .A(KEYINPUT96), .B(KEYINPUT93), .Z(n331) );
  XNOR2_X1 U386 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n348) );
  XOR2_X1 U389 ( .A(G148GAT), .B(G57GAT), .Z(n378) );
  XOR2_X1 U390 ( .A(n378), .B(n334), .Z(n336) );
  XNOR2_X1 U391 ( .A(G134GAT), .B(G162GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n344) );
  XOR2_X1 U393 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n342) );
  XOR2_X1 U394 ( .A(KEYINPUT83), .B(G127GAT), .Z(n338) );
  XNOR2_X1 U395 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U397 ( .A(G113GAT), .B(n339), .Z(n452) );
  XNOR2_X1 U398 ( .A(n452), .B(n340), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U400 ( .A(n344), .B(n343), .Z(n346) );
  NAND2_X1 U401 ( .A1(G225GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U403 ( .A(n348), .B(n347), .Z(n467) );
  XOR2_X1 U404 ( .A(KEYINPUT98), .B(n467), .Z(n514) );
  INV_X1 U405 ( .A(KEYINPUT54), .ZN(n439) );
  XOR2_X1 U406 ( .A(KEYINPUT47), .B(KEYINPUT113), .Z(n412) );
  XOR2_X1 U407 ( .A(G113GAT), .B(G141GAT), .Z(n350) );
  XNOR2_X1 U408 ( .A(G169GAT), .B(G197GAT), .ZN(n349) );
  XOR2_X1 U409 ( .A(n350), .B(n349), .Z(n366) );
  XOR2_X1 U410 ( .A(G29GAT), .B(G43GAT), .Z(n352) );
  XNOR2_X1 U411 ( .A(G50GAT), .B(G36GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n355) );
  XOR2_X1 U413 ( .A(G1GAT), .B(G8GAT), .Z(n354) );
  XNOR2_X1 U414 ( .A(G22GAT), .B(G15GAT), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n397) );
  XOR2_X1 U416 ( .A(n355), .B(n397), .Z(n364) );
  XOR2_X1 U417 ( .A(KEYINPUT70), .B(KEYINPUT67), .Z(n357) );
  XNOR2_X1 U418 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n357), .B(n356), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n358), .B(KEYINPUT68), .ZN(n360) );
  NAND2_X1 U421 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n570) );
  INV_X1 U426 ( .A(n570), .ZN(n550) );
  XOR2_X1 U427 ( .A(G176GAT), .B(G64GAT), .Z(n433) );
  XOR2_X1 U428 ( .A(G71GAT), .B(KEYINPUT13), .Z(n398) );
  XOR2_X1 U429 ( .A(n433), .B(n398), .Z(n370) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U431 ( .A(n370), .B(n369), .Z(n384) );
  XOR2_X1 U432 ( .A(KEYINPUT31), .B(KEYINPUT73), .Z(n372) );
  XNOR2_X1 U433 ( .A(G120GAT), .B(G204GAT), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n375) );
  XNOR2_X1 U435 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n373), .B(KEYINPUT32), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n377) );
  AND2_X1 U438 ( .A1(G230GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n382) );
  XNOR2_X1 U440 ( .A(G85GAT), .B(n378), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n416) );
  NOR2_X1 U442 ( .A1(n550), .A2(n556), .ZN(n386) );
  XNOR2_X1 U443 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n407) );
  XOR2_X1 U445 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n388) );
  XNOR2_X1 U446 ( .A(KEYINPUT15), .B(KEYINPUT81), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n406) );
  XOR2_X1 U448 ( .A(G78GAT), .B(G155GAT), .Z(n390) );
  XNOR2_X1 U449 ( .A(G127GAT), .B(G211GAT), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U451 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n392) );
  XNOR2_X1 U452 ( .A(G183GAT), .B(G64GAT), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U454 ( .A(n394), .B(n393), .Z(n404) );
  XOR2_X1 U455 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n396) );
  XNOR2_X1 U456 ( .A(G57GAT), .B(KEYINPUT79), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n402) );
  XOR2_X1 U458 ( .A(n398), .B(n397), .Z(n400) );
  NAND2_X1 U459 ( .A1(G231GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U463 ( .A(n406), .B(n405), .Z(n560) );
  INV_X1 U464 ( .A(n560), .ZN(n576) );
  NOR2_X1 U465 ( .A1(n407), .A2(n576), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n408), .B(KEYINPUT111), .ZN(n409) );
  NOR2_X1 U467 ( .A1(n546), .A2(n409), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n410), .B(KEYINPUT112), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n420) );
  XNOR2_X1 U470 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n415) );
  XNOR2_X1 U471 ( .A(KEYINPUT36), .B(KEYINPUT104), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n413), .B(n476), .ZN(n581) );
  NOR2_X1 U473 ( .A1(n581), .A2(n560), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n418) );
  NOR2_X1 U475 ( .A1(n570), .A2(n416), .ZN(n417) );
  NAND2_X1 U476 ( .A1(n418), .A2(n417), .ZN(n419) );
  NAND2_X1 U477 ( .A1(n420), .A2(n419), .ZN(n422) );
  XOR2_X1 U478 ( .A(KEYINPUT85), .B(KEYINPUT18), .Z(n424) );
  XNOR2_X1 U479 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U481 ( .A(n425), .B(KEYINPUT86), .Z(n427) );
  XNOR2_X1 U482 ( .A(G169GAT), .B(G183GAT), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n456) );
  XOR2_X1 U484 ( .A(KEYINPUT99), .B(n428), .Z(n431) );
  XNOR2_X1 U485 ( .A(G8GAT), .B(n429), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U487 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U488 ( .A1(G226GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n456), .B(n436), .ZN(n517) );
  XNOR2_X1 U491 ( .A(KEYINPUT117), .B(n517), .ZN(n437) );
  NOR2_X1 U492 ( .A1(n524), .A2(n437), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  NOR2_X1 U494 ( .A1(n514), .A2(n440), .ZN(n568) );
  NAND2_X1 U495 ( .A1(n469), .A2(n568), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n441), .B(KEYINPUT55), .ZN(n457) );
  XOR2_X1 U497 ( .A(KEYINPUT84), .B(G71GAT), .Z(n443) );
  XNOR2_X1 U498 ( .A(G99GAT), .B(G190GAT), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U500 ( .A(n444), .B(KEYINPUT87), .Z(n447) );
  XNOR2_X1 U501 ( .A(G15GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U503 ( .A(KEYINPUT65), .B(G176GAT), .Z(n449) );
  NAND2_X1 U504 ( .A1(G227GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U506 ( .A(n451), .B(n450), .Z(n454) );
  XNOR2_X1 U507 ( .A(n452), .B(KEYINPUT20), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n457), .A2(n525), .ZN(n559) );
  NOR2_X1 U510 ( .A1(n476), .A2(n559), .ZN(n460) );
  NOR2_X1 U511 ( .A1(n416), .A2(n550), .ZN(n491) );
  NOR2_X1 U512 ( .A1(n525), .A2(n469), .ZN(n461) );
  XNOR2_X1 U513 ( .A(n461), .B(KEYINPUT26), .ZN(n567) );
  XNOR2_X1 U514 ( .A(n517), .B(KEYINPUT27), .ZN(n470) );
  NAND2_X1 U515 ( .A1(n567), .A2(n470), .ZN(n466) );
  NAND2_X1 U516 ( .A1(n525), .A2(n517), .ZN(n462) );
  NAND2_X1 U517 ( .A1(n462), .A2(n469), .ZN(n463) );
  XNOR2_X1 U518 ( .A(n463), .B(KEYINPUT100), .ZN(n464) );
  XOR2_X1 U519 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NAND2_X1 U520 ( .A1(n466), .A2(n465), .ZN(n468) );
  NAND2_X1 U521 ( .A1(n468), .A2(n467), .ZN(n474) );
  XOR2_X1 U522 ( .A(KEYINPUT88), .B(n525), .Z(n472) );
  NAND2_X1 U523 ( .A1(n470), .A2(n514), .ZN(n523) );
  NOR2_X1 U524 ( .A1(n527), .A2(n523), .ZN(n471) );
  NAND2_X1 U525 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U526 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U527 ( .A(KEYINPUT101), .B(n475), .ZN(n488) );
  INV_X1 U528 ( .A(n476), .ZN(n535) );
  NOR2_X1 U529 ( .A1(n535), .A2(n560), .ZN(n477) );
  XOR2_X1 U530 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  NOR2_X1 U531 ( .A1(n488), .A2(n478), .ZN(n502) );
  AND2_X1 U532 ( .A1(n491), .A2(n502), .ZN(n485) );
  NAND2_X1 U533 ( .A1(n514), .A2(n485), .ZN(n481) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n479), .B(KEYINPUT102), .ZN(n480) );
  XNOR2_X1 U536 ( .A(n481), .B(n480), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n517), .A2(n485), .ZN(n482) );
  XNOR2_X1 U538 ( .A(n482), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U540 ( .A1(n485), .A2(n525), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  XOR2_X1 U542 ( .A(G22GAT), .B(KEYINPUT103), .Z(n487) );
  NAND2_X1 U543 ( .A1(n485), .A2(n527), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n494) );
  NOR2_X1 U546 ( .A1(n581), .A2(n488), .ZN(n489) );
  NAND2_X1 U547 ( .A1(n560), .A2(n489), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n490), .ZN(n513) );
  NAND2_X1 U549 ( .A1(n513), .A2(n491), .ZN(n492) );
  XOR2_X1 U550 ( .A(KEYINPUT38), .B(n492), .Z(n500) );
  NAND2_X1 U551 ( .A1(n290), .A2(n514), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U553 ( .A(G29GAT), .B(n495), .Z(G1328GAT) );
  NAND2_X1 U554 ( .A1(n290), .A2(n517), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(KEYINPUT106), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n290), .A2(n525), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(KEYINPUT40), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n290), .A2(n527), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U562 ( .A1(n570), .A2(n556), .ZN(n512) );
  NAND2_X1 U563 ( .A1(n502), .A2(n512), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(KEYINPUT107), .ZN(n509) );
  NAND2_X1 U565 ( .A1(n509), .A2(n514), .ZN(n504) );
  XNOR2_X1 U566 ( .A(KEYINPUT42), .B(n504), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U568 ( .A1(n517), .A2(n509), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n506), .B(KEYINPUT108), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(n507), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n525), .A2(n509), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U574 ( .A1(n509), .A2(n527), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  XOR2_X1 U576 ( .A(G85GAT), .B(KEYINPUT109), .Z(n516) );
  AND2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n520), .A2(n514), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n520), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n525), .A2(n520), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n527), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n524), .A2(n523), .ZN(n540) );
  NAND2_X1 U588 ( .A1(n540), .A2(n525), .ZN(n526) );
  NOR2_X1 U589 ( .A1(n527), .A2(n526), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n536), .A2(n570), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n528), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  INV_X1 U593 ( .A(n556), .ZN(n529) );
  NAND2_X1 U594 ( .A1(n536), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n533) );
  NAND2_X1 U597 ( .A1(n536), .A2(n576), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n540), .A2(n567), .ZN(n547) );
  NOR2_X1 U605 ( .A1(n550), .A2(n547), .ZN(n541) );
  XOR2_X1 U606 ( .A(G141GAT), .B(n541), .Z(G1344GAT) );
  NOR2_X1 U607 ( .A1(n556), .A2(n547), .ZN(n543) );
  XNOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n544), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n560), .A2(n547), .ZN(n545) );
  XOR2_X1 U612 ( .A(G155GAT), .B(n545), .Z(G1346GAT) );
  INV_X1 U613 ( .A(n546), .ZN(n548) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U615 ( .A(G162GAT), .B(n549), .Z(G1347GAT) );
  XNOR2_X1 U616 ( .A(G169GAT), .B(KEYINPUT118), .ZN(n553) );
  NOR2_X1 U617 ( .A1(n559), .A2(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n555) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n558) );
  NOR2_X1 U623 ( .A1(n556), .A2(n559), .ZN(n557) );
  XOR2_X1 U624 ( .A(n558), .B(n557), .Z(G1349GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U626 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G183GAT), .B(n563), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n565) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT59), .B(n566), .Z(n572) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT123), .B(n569), .Z(n580) );
  INV_X1 U635 ( .A(n580), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U639 ( .A1(n577), .A2(n416), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n575), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(n582), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

