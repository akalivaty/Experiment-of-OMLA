

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581;

  XOR2_X1 U323 ( .A(n306), .B(n305), .Z(n566) );
  XNOR2_X1 U324 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U325 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n385) );
  XNOR2_X1 U326 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U327 ( .A(n386), .B(n385), .ZN(n410) );
  INV_X1 U328 ( .A(G218GAT), .ZN(n446) );
  NOR2_X1 U329 ( .A1(n553), .A2(n455), .ZN(n580) );
  XOR2_X1 U330 ( .A(KEYINPUT93), .B(n465), .Z(n542) );
  XNOR2_X1 U331 ( .A(n446), .B(KEYINPUT62), .ZN(n447) );
  XNOR2_X1 U332 ( .A(n448), .B(n447), .ZN(G1355GAT) );
  XNOR2_X1 U333 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n291) );
  XNOR2_X1 U334 ( .A(n291), .B(KEYINPUT7), .ZN(n350) );
  XNOR2_X1 U335 ( .A(G36GAT), .B(G190GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n292), .B(G218GAT), .ZN(n381) );
  XNOR2_X1 U337 ( .A(n350), .B(n381), .ZN(n306) );
  XOR2_X1 U338 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n294) );
  XOR2_X1 U339 ( .A(G50GAT), .B(G162GAT), .Z(n412) );
  XOR2_X1 U340 ( .A(G99GAT), .B(G85GAT), .Z(n315) );
  XNOR2_X1 U341 ( .A(n412), .B(n315), .ZN(n293) );
  XNOR2_X1 U342 ( .A(n294), .B(n293), .ZN(n300) );
  XOR2_X1 U343 ( .A(KEYINPUT70), .B(KEYINPUT9), .Z(n296) );
  XNOR2_X1 U344 ( .A(G106GAT), .B(G92GAT), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n296), .B(n295), .ZN(n298) );
  AND2_X1 U346 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XOR2_X1 U347 ( .A(n301), .B(KEYINPUT72), .Z(n304) );
  XNOR2_X1 U348 ( .A(G29GAT), .B(G134GAT), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n302), .B(KEYINPUT71), .ZN(n403) );
  XNOR2_X1 U350 ( .A(n403), .B(KEYINPUT10), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U352 ( .A(KEYINPUT36), .B(n566), .Z(n481) );
  XNOR2_X1 U353 ( .A(G120GAT), .B(G148GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n307), .B(G57GAT), .ZN(n393) );
  XOR2_X1 U355 ( .A(G71GAT), .B(KEYINPUT13), .Z(n332) );
  XOR2_X1 U356 ( .A(n393), .B(n332), .Z(n311) );
  XOR2_X1 U357 ( .A(G106GAT), .B(G78GAT), .Z(n411) );
  XOR2_X1 U358 ( .A(G64GAT), .B(G92GAT), .Z(n309) );
  XNOR2_X1 U359 ( .A(G176GAT), .B(G204GAT), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n376) );
  XNOR2_X1 U361 ( .A(n411), .B(n376), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n319) );
  XOR2_X1 U363 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n313) );
  XNOR2_X1 U364 ( .A(KEYINPUT69), .B(KEYINPUT33), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U366 ( .A(n315), .B(n314), .Z(n317) );
  NAND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n319), .B(n318), .ZN(n575) );
  XOR2_X1 U370 ( .A(G1GAT), .B(G8GAT), .Z(n321) );
  XNOR2_X1 U371 ( .A(G22GAT), .B(G15GAT), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n346) );
  XOR2_X1 U373 ( .A(n346), .B(KEYINPUT75), .Z(n323) );
  NAND2_X1 U374 ( .A1(G231GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n339) );
  XOR2_X1 U376 ( .A(KEYINPUT77), .B(KEYINPUT73), .Z(n325) );
  XNOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT76), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U379 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n327) );
  XNOR2_X1 U380 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n337) );
  XOR2_X1 U383 ( .A(G78GAT), .B(G211GAT), .Z(n331) );
  XNOR2_X1 U384 ( .A(G127GAT), .B(G155GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n333) );
  XOR2_X1 U386 ( .A(n333), .B(n332), .Z(n335) );
  XNOR2_X1 U387 ( .A(G183GAT), .B(G64GAT), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U390 ( .A(n339), .B(n338), .Z(n579) );
  INV_X1 U391 ( .A(n579), .ZN(n479) );
  OR2_X1 U392 ( .A1(n481), .A2(n479), .ZN(n340) );
  XNOR2_X1 U393 ( .A(KEYINPUT45), .B(n340), .ZN(n341) );
  NOR2_X1 U394 ( .A1(n575), .A2(n341), .ZN(n359) );
  XOR2_X1 U395 ( .A(KEYINPUT65), .B(G113GAT), .Z(n343) );
  XNOR2_X1 U396 ( .A(G169GAT), .B(G197GAT), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n358) );
  XOR2_X1 U398 ( .A(G50GAT), .B(G29GAT), .Z(n345) );
  XNOR2_X1 U399 ( .A(G36GAT), .B(G141GAT), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n347) );
  XOR2_X1 U401 ( .A(n347), .B(n346), .Z(n356) );
  XOR2_X1 U402 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n349) );
  XNOR2_X1 U403 ( .A(KEYINPUT66), .B(KEYINPUT68), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n354) );
  XOR2_X1 U405 ( .A(n350), .B(KEYINPUT67), .Z(n352) );
  NAND2_X1 U406 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n358), .B(n357), .ZN(n497) );
  NAND2_X1 U411 ( .A1(n359), .A2(n497), .ZN(n367) );
  XOR2_X1 U412 ( .A(KEYINPUT114), .B(KEYINPUT47), .Z(n365) );
  XOR2_X1 U413 ( .A(KEYINPUT41), .B(n575), .Z(n562) );
  INV_X1 U414 ( .A(n497), .ZN(n570) );
  AND2_X1 U415 ( .A1(n562), .A2(n570), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n360), .B(KEYINPUT46), .ZN(n361) );
  NOR2_X1 U417 ( .A1(n579), .A2(n361), .ZN(n363) );
  INV_X1 U418 ( .A(n566), .ZN(n362) );
  NAND2_X1 U419 ( .A1(n363), .A2(n362), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n366) );
  NAND2_X1 U421 ( .A1(n367), .A2(n366), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n368), .B(KEYINPUT48), .ZN(n540) );
  XOR2_X1 U423 ( .A(KEYINPUT80), .B(KEYINPUT18), .Z(n370) );
  XNOR2_X1 U424 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U426 ( .A(n371), .B(KEYINPUT81), .Z(n373) );
  XNOR2_X1 U427 ( .A(G169GAT), .B(G183GAT), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n442) );
  XOR2_X1 U429 ( .A(G8GAT), .B(KEYINPUT94), .Z(n375) );
  NAND2_X1 U430 ( .A1(G226GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U432 ( .A(n377), .B(n376), .Z(n383) );
  XOR2_X1 U433 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n379) );
  XNOR2_X1 U434 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U436 ( .A(G197GAT), .B(n380), .Z(n416) );
  XNOR2_X1 U437 ( .A(n416), .B(n381), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U439 ( .A(n442), .B(n384), .ZN(n516) );
  INV_X1 U440 ( .A(n516), .ZN(n457) );
  NAND2_X1 U441 ( .A1(n540), .A2(n457), .ZN(n386) );
  XOR2_X1 U442 ( .A(KEYINPUT92), .B(KEYINPUT89), .Z(n388) );
  XNOR2_X1 U443 ( .A(G1GAT), .B(KEYINPUT91), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n390) );
  XOR2_X1 U445 ( .A(G162GAT), .B(G85GAT), .Z(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n407) );
  XOR2_X1 U447 ( .A(KEYINPUT5), .B(KEYINPUT88), .Z(n392) );
  XNOR2_X1 U448 ( .A(KEYINPUT90), .B(KEYINPUT1), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U450 ( .A(n394), .B(n393), .Z(n401) );
  XOR2_X1 U451 ( .A(G127GAT), .B(KEYINPUT78), .Z(n396) );
  XNOR2_X1 U452 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n431) );
  XOR2_X1 U454 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n398) );
  XNOR2_X1 U455 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U457 ( .A(G141GAT), .B(n399), .Z(n426) );
  XNOR2_X1 U458 ( .A(n431), .B(n426), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U460 ( .A(n402), .B(KEYINPUT4), .Z(n405) );
  XNOR2_X1 U461 ( .A(n403), .B(KEYINPUT6), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n409) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n465) );
  NAND2_X1 U466 ( .A1(n410), .A2(n542), .ZN(n553) );
  XOR2_X1 U467 ( .A(KEYINPUT87), .B(G218GAT), .Z(n414) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U470 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U471 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U473 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n420) );
  XNOR2_X1 U474 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U476 ( .A(n422), .B(n421), .Z(n428) );
  XOR2_X1 U477 ( .A(G148GAT), .B(KEYINPUT23), .Z(n424) );
  XNOR2_X1 U478 ( .A(G22GAT), .B(G204GAT), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n554) );
  XOR2_X1 U482 ( .A(G99GAT), .B(G134GAT), .Z(n430) );
  NAND2_X1 U483 ( .A1(G227GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U485 ( .A(n432), .B(n431), .Z(n440) );
  XOR2_X1 U486 ( .A(KEYINPUT20), .B(KEYINPUT79), .Z(n434) );
  XNOR2_X1 U487 ( .A(G43GAT), .B(G190GAT), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U489 ( .A(G120GAT), .B(G71GAT), .Z(n436) );
  XNOR2_X1 U490 ( .A(G15GAT), .B(G176GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n523) );
  INV_X1 U495 ( .A(n523), .ZN(n557) );
  NAND2_X1 U496 ( .A1(n554), .A2(n557), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n443), .B(KEYINPUT96), .ZN(n444) );
  XNOR2_X1 U498 ( .A(KEYINPUT26), .B(n444), .ZN(n455) );
  INV_X1 U499 ( .A(n580), .ZN(n445) );
  NOR2_X1 U500 ( .A1(n481), .A2(n445), .ZN(n448) );
  XOR2_X1 U501 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n450) );
  XNOR2_X1 U502 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n471) );
  NOR2_X1 U504 ( .A1(n497), .A2(n575), .ZN(n484) );
  NOR2_X1 U505 ( .A1(n566), .A2(n479), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n451), .B(KEYINPUT16), .ZN(n468) );
  XOR2_X1 U507 ( .A(n554), .B(KEYINPUT28), .Z(n520) );
  XOR2_X1 U508 ( .A(n516), .B(KEYINPUT27), .Z(n454) );
  NAND2_X1 U509 ( .A1(n520), .A2(n454), .ZN(n452) );
  OR2_X1 U510 ( .A1(n542), .A2(n452), .ZN(n525) );
  XNOR2_X1 U511 ( .A(KEYINPUT95), .B(n525), .ZN(n453) );
  NAND2_X1 U512 ( .A1(n557), .A2(n453), .ZN(n467) );
  INV_X1 U513 ( .A(n454), .ZN(n456) );
  NOR2_X1 U514 ( .A1(n456), .A2(n455), .ZN(n539) );
  XNOR2_X1 U515 ( .A(n539), .B(KEYINPUT97), .ZN(n463) );
  NAND2_X1 U516 ( .A1(n457), .A2(n523), .ZN(n458) );
  XOR2_X1 U517 ( .A(KEYINPUT98), .B(n458), .Z(n459) );
  NOR2_X1 U518 ( .A1(n554), .A2(n459), .ZN(n461) );
  XOR2_X1 U519 ( .A(KEYINPUT99), .B(KEYINPUT25), .Z(n460) );
  XNOR2_X1 U520 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n478) );
  NAND2_X1 U524 ( .A1(n468), .A2(n478), .ZN(n498) );
  INV_X1 U525 ( .A(n498), .ZN(n469) );
  NAND2_X1 U526 ( .A1(n484), .A2(n469), .ZN(n476) );
  NOR2_X1 U527 ( .A1(n542), .A2(n476), .ZN(n470) );
  XOR2_X1 U528 ( .A(n471), .B(n470), .Z(G1324GAT) );
  NOR2_X1 U529 ( .A1(n516), .A2(n476), .ZN(n472) );
  XOR2_X1 U530 ( .A(G8GAT), .B(n472), .Z(G1325GAT) );
  NOR2_X1 U531 ( .A1(n557), .A2(n476), .ZN(n474) );
  XNOR2_X1 U532 ( .A(KEYINPUT35), .B(KEYINPUT102), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(n475), .ZN(G1326GAT) );
  NOR2_X1 U535 ( .A1(n520), .A2(n476), .ZN(n477) );
  XOR2_X1 U536 ( .A(G22GAT), .B(n477), .Z(G1327GAT) );
  NAND2_X1 U537 ( .A1(n479), .A2(n478), .ZN(n480) );
  NOR2_X1 U538 ( .A1(n481), .A2(n480), .ZN(n483) );
  XNOR2_X1 U539 ( .A(KEYINPUT37), .B(KEYINPUT103), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(n513) );
  NAND2_X1 U541 ( .A1(n484), .A2(n513), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(KEYINPUT38), .ZN(n491) );
  NOR2_X1 U543 ( .A1(n542), .A2(n491), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n486), .B(KEYINPUT39), .ZN(n487) );
  XNOR2_X1 U545 ( .A(G29GAT), .B(n487), .ZN(G1328GAT) );
  NOR2_X1 U546 ( .A1(n491), .A2(n516), .ZN(n488) );
  XOR2_X1 U547 ( .A(G36GAT), .B(n488), .Z(G1329GAT) );
  NOR2_X1 U548 ( .A1(n557), .A2(n491), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT40), .B(n489), .Z(n490) );
  XNOR2_X1 U550 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  XNOR2_X1 U551 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n493) );
  NOR2_X1 U552 ( .A1(n520), .A2(n491), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G50GAT), .B(n494), .ZN(G1331GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n496) );
  XNOR2_X1 U556 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n501) );
  NAND2_X1 U558 ( .A1(n497), .A2(n562), .ZN(n511) );
  NOR2_X1 U559 ( .A1(n498), .A2(n511), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(KEYINPUT107), .ZN(n506) );
  NOR2_X1 U561 ( .A1(n542), .A2(n506), .ZN(n500) );
  XOR2_X1 U562 ( .A(n501), .B(n500), .Z(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT106), .B(n502), .ZN(G1332GAT) );
  NOR2_X1 U564 ( .A1(n516), .A2(n506), .ZN(n503) );
  XOR2_X1 U565 ( .A(G64GAT), .B(n503), .Z(G1333GAT) );
  NOR2_X1 U566 ( .A1(n557), .A2(n506), .ZN(n504) );
  XOR2_X1 U567 ( .A(KEYINPUT110), .B(n504), .Z(n505) );
  XNOR2_X1 U568 ( .A(G71GAT), .B(n505), .ZN(G1334GAT) );
  NOR2_X1 U569 ( .A1(n506), .A2(n520), .ZN(n510) );
  XOR2_X1 U570 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n508) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT112), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  INV_X1 U574 ( .A(n511), .ZN(n512) );
  NAND2_X1 U575 ( .A1(n513), .A2(n512), .ZN(n519) );
  NOR2_X1 U576 ( .A1(n542), .A2(n519), .ZN(n515) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n516), .A2(n519), .ZN(n517) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n517), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n557), .A2(n519), .ZN(n518) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(n521), .Z(n522) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  XOR2_X1 U586 ( .A(G113GAT), .B(KEYINPUT115), .Z(n527) );
  NAND2_X1 U587 ( .A1(n540), .A2(n523), .ZN(n524) );
  NOR2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n534), .A2(n570), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n527), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U592 ( .A1(n534), .A2(n562), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G120GAT), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n532) );
  NAND2_X1 U596 ( .A1(n534), .A2(n579), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U600 ( .A1(n534), .A2(n566), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n538) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT118), .Z(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n551), .A2(n570), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n543), .B(KEYINPUT120), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n546) );
  NAND2_X1 U610 ( .A1(n551), .A2(n562), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT53), .Z(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n551), .A2(n579), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n549), .B(KEYINPUT122), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n566), .A2(n551), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT55), .ZN(n556) );
  NOR2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n567) );
  NAND2_X1 U622 ( .A1(n570), .A2(n567), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n560) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT124), .B(n561), .Z(n564) );
  NAND2_X1 U628 ( .A1(n567), .A2(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n567), .A2(n579), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1351GAT) );
  NAND2_X1 U635 ( .A1(n580), .A2(n570), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n577) );
  NAND2_X1 U641 ( .A1(n580), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n578), .Z(G1353GAT) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
endmodule

