//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT65), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT66), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(new_n463), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  OR2_X1    g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(G101), .A3(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n475), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NAND3_X1  g057(.A1(new_n468), .A2(G2105), .A3(new_n472), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT67), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(new_n478), .A2(G112), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n474), .A2(G136), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n486), .A2(new_n490), .ZN(G162));
  AND2_X1   g066(.A1(KEYINPUT68), .A2(G114), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT68), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2105), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n483), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n478), .A2(G138), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n472), .A2(new_n464), .A3(new_n467), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n468), .A2(KEYINPUT69), .A3(new_n472), .A4(new_n500), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(KEYINPUT4), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n476), .A2(new_n506), .A3(new_n500), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n499), .B1(new_n505), .B2(new_n507), .ZN(G164));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n509), .A2(new_n510), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n514), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n519), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n517), .B(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n513), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n528), .B(new_n530), .C1(new_n531), .C2(new_n518), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n527), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n521), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n513), .A2(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n537), .B2(new_n518), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G171));
  INV_X1    g114(.A(new_n518), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT71), .B(G43), .Z(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(G81), .B1(new_n513), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n543), .B2(new_n521), .ZN(new_n544));
  XOR2_X1   g119(.A(new_n544), .B(KEYINPUT72), .Z(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  XNOR2_X1  g125(.A(new_n517), .B(KEYINPUT74), .ZN(new_n551));
  INV_X1    g126(.A(G65), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(G78), .A2(G543), .ZN(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(KEYINPUT75), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n555), .A2(KEYINPUT75), .B1(G91), .B2(new_n540), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n513), .A2(G53), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT9), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT73), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  XNOR2_X1  g139(.A(new_n517), .B(KEYINPUT70), .ZN(new_n565));
  INV_X1    g140(.A(G74), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n521), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n513), .A2(G49), .ZN(new_n568));
  INV_X1    g143(.A(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n569), .B2(new_n518), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n567), .A2(new_n570), .ZN(G288));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  OR3_X1    g147(.A1(new_n518), .A2(KEYINPUT76), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n517), .A2(G61), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(new_n513), .B2(G48), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT76), .B1(new_n518), .B2(new_n572), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n521), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n540), .A2(G85), .B1(new_n513), .B2(G47), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(new_n540), .A2(G92), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT10), .Z(new_n585));
  INV_X1    g160(.A(G66), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n551), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g162(.A1(G79), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n513), .A2(G54), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n592), .B2(G171), .ZN(G284));
  OAI21_X1  g169(.A(new_n593), .B1(new_n592), .B2(G171), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n558), .A2(new_n561), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  XOR2_X1   g173(.A(G297), .B(KEYINPUT77), .Z(G280));
  INV_X1    g174(.A(new_n591), .ZN(new_n600));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G860), .ZN(G148));
  INV_X1    g177(.A(new_n545), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(new_n592), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n591), .A2(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n592), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n474), .A2(G135), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n478), .A2(G111), .ZN(new_n609));
  OAI21_X1  g184(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n610));
  INV_X1    g185(.A(G123), .ZN(new_n611));
  OAI221_X1 g186(.A(new_n608), .B1(new_n609), .B2(new_n610), .C1(new_n484), .C2(new_n611), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(G2096), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(G2096), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n478), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(G156));
  XOR2_X1   g194(.A(KEYINPUT15), .B(G2435), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2438), .ZN(new_n621));
  XOR2_X1   g196(.A(G2427), .B(G2430), .Z(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT79), .B(KEYINPUT14), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n621), .A2(new_n622), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT80), .Z(new_n627));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n627), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(new_n637), .A3(G14), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g216(.A1(G2072), .A2(G2078), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n442), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n641), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT18), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n643), .A2(KEYINPUT81), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(KEYINPUT81), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(new_n645), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n643), .B(KEYINPUT17), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n650), .B(new_n641), .C1(new_n651), .C2(new_n645), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n645), .A3(new_n640), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n647), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n658), .A2(new_n661), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT20), .Z(new_n665));
  AOI211_X1 g240(.A(new_n663), .B(new_n665), .C1(new_n658), .C2(new_n662), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  XNOR2_X1  g247(.A(KEYINPUT82), .B(G29), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n674), .A2(G35), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(G162), .B2(new_n674), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2090), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n485), .A2(G129), .ZN(new_n680));
  NAND3_X1  g255(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT26), .ZN(new_n682));
  AND3_X1   g257(.A1(new_n478), .A2(G105), .A3(G2104), .ZN(new_n683));
  AOI211_X1 g258(.A(new_n682), .B(new_n683), .C1(new_n474), .C2(G141), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n687), .B2(G32), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT27), .B(G1996), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G5), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G171), .B2(new_n692), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(G1961), .ZN(new_n695));
  NOR2_X1   g270(.A1(G4), .A2(G16), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n600), .B2(G16), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n695), .B1(new_n697), .B2(G1348), .ZN(new_n698));
  INV_X1    g273(.A(new_n697), .ZN(new_n699));
  INV_X1    g274(.A(G1348), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n699), .A2(new_n700), .B1(G1961), .B2(new_n694), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n702), .A2(G28), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n687), .B1(new_n702), .B2(G28), .ZN(new_n704));
  NOR2_X1   g279(.A1(KEYINPUT31), .A2(G11), .ZN(new_n705));
  AND2_X1   g280(.A1(KEYINPUT31), .A2(G11), .ZN(new_n706));
  OAI22_X1  g281(.A1(new_n703), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n692), .A2(G21), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G168), .B2(new_n692), .ZN(new_n709));
  OAI22_X1  g284(.A1(new_n612), .A2(new_n673), .B1(new_n709), .B2(G1966), .ZN(new_n710));
  AOI211_X1 g285(.A(new_n707), .B(new_n710), .C1(G1966), .C2(new_n709), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n691), .A2(new_n698), .A3(new_n701), .A4(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n545), .A2(new_n692), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n692), .B2(G19), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n679), .B(new_n712), .C1(G1341), .C2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(G34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(G34), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n718), .A2(new_n673), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n481), .B2(new_n687), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT90), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(G2084), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT92), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT87), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT25), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n474), .A2(G139), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n728), .B(new_n729), .C1(new_n478), .C2(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(G33), .B(new_n731), .S(G29), .Z(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT88), .Z(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(G2072), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(G2072), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n689), .A2(new_n690), .B1(G2084), .B2(new_n722), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n716), .B(new_n724), .C1(new_n725), .C2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n725), .B2(new_n737), .ZN(new_n739));
  MUX2_X1   g314(.A(G24), .B(G290), .S(G16), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1986), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n673), .A2(G25), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n485), .A2(G119), .ZN(new_n743));
  NOR2_X1   g318(.A1(G95), .A2(G2105), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT83), .Z(new_n745));
  INV_X1    g320(.A(G107), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n466), .B1(new_n746), .B2(G2105), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n474), .A2(G131), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n742), .B1(new_n749), .B2(new_n674), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT35), .B(G1991), .Z(new_n751));
  AOI21_X1  g326(.A(new_n741), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n692), .A2(G22), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G166), .B2(new_n692), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1971), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n692), .A2(G23), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n567), .A2(new_n570), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n692), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT33), .B(G1976), .Z(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n692), .A2(G6), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G305), .B2(G16), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT32), .B(G1981), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n760), .A2(new_n761), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n763), .A2(new_n765), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n755), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT34), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n750), .A2(new_n751), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n752), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(KEYINPUT84), .A2(KEYINPUT36), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n774), .B(new_n775), .Z(new_n776));
  NOR2_X1   g351(.A1(G164), .A2(new_n673), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G27), .B2(new_n673), .ZN(new_n778));
  INV_X1    g353(.A(G2078), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n780), .B(new_n781), .C1(new_n715), .C2(G1341), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n692), .A2(G20), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT23), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n597), .B2(new_n692), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1956), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n673), .A2(G26), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n478), .A2(G116), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n474), .A2(G140), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G128), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n484), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT85), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(G29), .ZN(new_n798));
  INV_X1    g373(.A(G2067), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n782), .A2(new_n786), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n739), .A2(new_n776), .A3(new_n801), .ZN(G150));
  INV_X1    g377(.A(G150), .ZN(G311));
  NAND2_X1  g378(.A1(new_n526), .A2(G67), .ZN(new_n804));
  NAND2_X1  g379(.A1(G80), .A2(G543), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n521), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n540), .A2(G93), .B1(new_n513), .B2(G55), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT95), .ZN(new_n810));
  INV_X1    g385(.A(new_n806), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n811), .A2(new_n812), .A3(new_n807), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n545), .B2(new_n809), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n810), .A2(new_n544), .A3(new_n813), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n544), .A2(KEYINPUT72), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n544), .A2(KEYINPUT72), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n820), .A2(new_n817), .A3(new_n821), .A4(new_n809), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n591), .A2(new_n601), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n824), .B(new_n826), .Z(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  INV_X1    g404(.A(G860), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n828), .B2(KEYINPUT39), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n816), .B1(new_n829), .B2(new_n831), .ZN(G145));
  NOR2_X1   g407(.A1(new_n731), .A2(KEYINPUT97), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT96), .Z(new_n834));
  AND2_X1   g409(.A1(new_n501), .A2(new_n502), .ZN(new_n835));
  OAI21_X1  g410(.A(KEYINPUT4), .B1(new_n501), .B2(new_n502), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n507), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n499), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n834), .A2(new_n839), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n749), .B(new_n616), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n840), .B2(new_n841), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n796), .B(new_n686), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n474), .A2(G142), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT98), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n485), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n478), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n847), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n844), .B2(new_n845), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n612), .B(G160), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G162), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n859), .B1(new_n855), .B2(new_n857), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g440(.A(new_n824), .B(new_n605), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n597), .A2(KEYINPUT99), .A3(new_n591), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(G299), .B2(new_n600), .ZN(new_n869));
  NAND2_X1  g444(.A1(G299), .A2(new_n600), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n867), .A2(KEYINPUT41), .A3(new_n869), .A4(new_n870), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n866), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n871), .B2(new_n866), .ZN(new_n876));
  XNOR2_X1  g451(.A(G290), .B(G305), .ZN(new_n877));
  XNOR2_X1  g452(.A(G288), .B(G303), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(KEYINPUT101), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT100), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT42), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n881), .A2(new_n884), .B1(new_n882), .B2(new_n880), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n592), .B1(new_n876), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n876), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(KEYINPUT102), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n814), .B2(new_n592), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n887), .B2(new_n890), .ZN(G295));
  AOI21_X1  g466(.A(new_n888), .B1(new_n887), .B2(new_n890), .ZN(G331));
  NAND2_X1  g467(.A1(new_n873), .A2(new_n874), .ZN(new_n893));
  OAI21_X1  g468(.A(G171), .B1(new_n818), .B2(new_n823), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n818), .A2(new_n823), .A3(G171), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n895), .A2(G286), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n824), .A2(G301), .ZN(new_n898));
  AOI21_X1  g473(.A(G168), .B1(new_n898), .B2(new_n894), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n893), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(G286), .B1(new_n895), .B2(new_n896), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(G168), .A3(new_n894), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n871), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n879), .B(KEYINPUT100), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n905), .A2(new_n861), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n900), .A2(new_n903), .ZN(new_n907));
  INV_X1    g482(.A(new_n904), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT43), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n861), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n873), .A2(new_n912), .A3(new_n874), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n871), .A2(KEYINPUT103), .A3(new_n872), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n913), .B(new_n914), .C1(new_n897), .C2(new_n899), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n904), .B1(new_n915), .B2(new_n903), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT44), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n917), .B1(new_n906), .B2(new_n909), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n911), .A2(new_n916), .A3(KEYINPUT43), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n923), .ZN(G397));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n925));
  XOR2_X1   g500(.A(KEYINPUT104), .B(G1384), .Z(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(G164), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n475), .A2(new_n479), .A3(G40), .A4(new_n480), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(G290), .A2(G1986), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT105), .ZN(new_n934));
  AND2_X1   g509(.A1(G290), .A2(G1986), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT106), .Z(new_n937));
  XNOR2_X1  g512(.A(new_n796), .B(G2067), .ZN(new_n938));
  INV_X1    g513(.A(G1996), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n685), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n749), .B(new_n751), .Z(new_n942));
  OAI21_X1  g517(.A(new_n932), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT125), .ZN(new_n945));
  INV_X1    g520(.A(G8), .ZN(new_n946));
  INV_X1    g521(.A(G1966), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n925), .B1(G164), .B2(G1384), .ZN(new_n948));
  NOR3_X1   g523(.A1(G164), .A2(new_n925), .A3(G1384), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT115), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n930), .B(new_n948), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G1384), .B1(new_n837), .B2(new_n838), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n950), .A3(KEYINPUT45), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n947), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G2084), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  INV_X1    g533(.A(new_n507), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n960), .B2(new_n503), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n957), .B(new_n958), .C1(new_n961), .C2(new_n499), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n963));
  AND4_X1   g538(.A1(new_n956), .A2(new_n962), .A3(new_n963), .A4(new_n930), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n946), .B1(new_n955), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(G286), .A2(G8), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT120), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT51), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n967), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(KEYINPUT51), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n966), .B2(KEYINPUT121), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT45), .B(new_n958), .C1(new_n961), .C2(new_n499), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT115), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n974), .A2(new_n930), .A3(new_n953), .A4(new_n948), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n964), .B1(new_n975), .B2(new_n947), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT121), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n976), .A2(new_n977), .A3(new_n946), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n969), .B1(new_n972), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n976), .A2(new_n967), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(G164), .A2(new_n926), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT45), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n984), .A2(new_n779), .A3(new_n930), .A4(new_n948), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT123), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(KEYINPUT123), .A3(new_n986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n839), .A2(new_n958), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n929), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n962), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT122), .B(G1961), .Z(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n986), .A2(G2078), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n991), .B(new_n996), .C1(new_n975), .C2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(G171), .B(KEYINPUT54), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n994), .B2(new_n995), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT124), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n928), .A2(new_n1003), .A3(new_n929), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT124), .B1(new_n927), .B2(new_n930), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n984), .B(new_n997), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n999), .A2(new_n1001), .B1(new_n1007), .B2(new_n991), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n982), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n963), .A2(new_n1012), .A3(new_n930), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n962), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(new_n963), .B2(new_n930), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n930), .B1(new_n952), .B2(new_n957), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT112), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(KEYINPUT113), .A3(new_n962), .A4(new_n1013), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT107), .B(G2090), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n984), .A2(new_n930), .A3(new_n948), .ZN(new_n1022));
  INV_X1    g597(.A(G1971), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n946), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G303), .A2(G8), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n1026), .B(KEYINPUT55), .Z(new_n1027));
  OAI21_X1  g602(.A(new_n1010), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1027), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1024), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1020), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1018), .A2(new_n962), .A3(new_n1013), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1032), .B2(new_n1011), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1030), .B1(new_n1033), .B2(new_n1019), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT114), .B(new_n1029), .C1(new_n1034), .C2(new_n946), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n952), .A2(new_n930), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n576), .A2(G651), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n513), .A2(G48), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n518), .A2(new_n572), .ZN(new_n1041));
  OAI21_X1  g616(.A(G1981), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1981), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n573), .A2(new_n577), .A3(new_n1043), .A4(new_n578), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1042), .A2(new_n1044), .A3(KEYINPUT49), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT111), .B1(new_n1037), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n946), .B1(new_n952), .B2(new_n930), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n1052), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n757), .A2(G1976), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT109), .B(G1976), .Z(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1036), .A2(G8), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1051), .A2(KEYINPUT110), .A3(new_n1057), .A4(new_n1055), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT52), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1054), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n993), .A2(new_n962), .A3(new_n1020), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1024), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(G8), .A3(new_n1027), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT108), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n946), .B1(new_n1024), .B2(new_n1066), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT108), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1027), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1065), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1028), .A2(new_n1035), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n945), .B1(new_n1009), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G1956), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1022), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT56), .B(G2072), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1032), .A2(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n558), .A2(new_n560), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1081));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1080), .A2(new_n1081), .B1(new_n1082), .B2(G299), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1036), .B(KEYINPUT118), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n799), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n994), .A2(new_n700), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(new_n591), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1084), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1088), .A2(KEYINPUT60), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1086), .A2(KEYINPUT60), .A3(new_n1087), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n600), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1094), .A3(new_n591), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1088), .A2(KEYINPUT119), .A3(KEYINPUT60), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1092), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1084), .A2(KEYINPUT61), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1084), .A2(KEYINPUT61), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1036), .B(new_n1103), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1077), .A2(new_n939), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n603), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1101), .A2(new_n1102), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1091), .B1(new_n1100), .B2(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1028), .A2(new_n1035), .A3(new_n1073), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n955), .A2(new_n965), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n977), .B1(new_n976), .B2(new_n946), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(new_n971), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n980), .B1(new_n1117), .B2(new_n969), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1007), .A2(new_n991), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n996), .B1(new_n975), .B2(new_n998), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n989), .B2(new_n990), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1121), .B2(new_n1000), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1113), .A2(new_n1123), .A3(KEYINPUT125), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1075), .A2(new_n1112), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n982), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n1118), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n999), .A2(G171), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1118), .B2(new_n1128), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1126), .A2(new_n1129), .A3(new_n1131), .A4(new_n1113), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n976), .A2(new_n946), .A3(G286), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1028), .A2(new_n1035), .A3(new_n1073), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1070), .A2(new_n1027), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n1065), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1138), .B(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1133), .A2(KEYINPUT63), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1136), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(G1976), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1054), .A2(new_n1146), .A3(new_n757), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1037), .B1(new_n1147), .B2(new_n1044), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1065), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1141), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1132), .A2(new_n1145), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n944), .B1(new_n1125), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n931), .B1(new_n938), .B2(new_n686), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT127), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n932), .A2(new_n939), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT46), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT47), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n934), .A2(new_n932), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT48), .Z(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n943), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n743), .A2(new_n751), .A3(new_n748), .ZN(new_n1162));
  OAI22_X1  g737(.A1(new_n941), .A2(new_n1162), .B1(G2067), .B2(new_n797), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n932), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1158), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1152), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g741(.A1(new_n921), .A2(new_n922), .ZN(new_n1168));
  NOR4_X1   g742(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1169));
  OAI21_X1  g743(.A(new_n1169), .B1(new_n863), .B2(new_n862), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n1168), .A2(new_n1170), .ZN(G308));
  OAI221_X1 g745(.A(new_n1169), .B1(new_n863), .B2(new_n862), .C1(new_n921), .C2(new_n922), .ZN(G225));
endmodule


