//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G141gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G197gat), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT11), .B(G169gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NOR3_X1   g011(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(KEYINPUT80), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  AND4_X1   g014(.A1(KEYINPUT80), .A2(new_n215), .A3(new_n208), .A4(new_n209), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n211), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G50gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G43gat), .ZN(new_n219));
  INV_X1    g018(.A(G43gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G50gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT15), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n210), .B1(new_n225), .B2(KEYINPUT15), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n220), .A2(G50gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n218), .A2(G43gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n212), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n231), .A2(new_n213), .A3(KEYINPUT81), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT81), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n208), .A3(new_n209), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(new_n212), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n226), .B(new_n230), .C1(new_n232), .C2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n224), .A2(KEYINPUT17), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G15gat), .B(G22gat), .ZN(new_n238));
  INV_X1    g037(.A(G1gat), .ZN(new_n239));
  AND3_X1   g038(.A1(new_n239), .A2(KEYINPUT83), .A3(KEYINPUT16), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT83), .B1(new_n239), .B2(KEYINPUT16), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n238), .B(KEYINPUT84), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT85), .B1(new_n238), .B2(G1gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT85), .ZN(new_n244));
  INV_X1    g043(.A(G15gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(G22gat), .ZN(new_n246));
  INV_X1    g045(.A(G22gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(G15gat), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n244), .B(new_n239), .C1(new_n246), .C2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n242), .A2(new_n243), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G8gat), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n239), .B(new_n251), .C1(new_n246), .C2(new_n248), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT83), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT16), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n253), .B1(new_n254), .B2(G1gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n239), .A2(KEYINPUT83), .A3(KEYINPUT16), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n257), .A2(new_n238), .B1(KEYINPUT84), .B2(G8gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n250), .A2(G8gat), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n237), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n224), .A2(new_n236), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT17), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT82), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT82), .ZN(new_n264));
  AOI211_X1 g063(.A(new_n264), .B(KEYINPUT17), .C1(new_n224), .C2(new_n236), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n260), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT86), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G229gat), .A2(G233gat), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n230), .A2(new_n222), .A3(new_n211), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT81), .B1(new_n231), .B2(new_n213), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n234), .A2(new_n233), .A3(new_n212), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n270), .A2(new_n273), .B1(new_n217), .B2(new_n223), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n259), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n264), .B1(new_n274), .B2(KEYINPUT17), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n261), .A2(KEYINPUT82), .A3(new_n262), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(KEYINPUT86), .A3(new_n260), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n268), .A2(new_n269), .A3(new_n276), .A4(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT18), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n269), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(new_n282), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n268), .A2(new_n276), .A3(new_n280), .A4(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT87), .B(KEYINPUT13), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(new_n284), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n259), .A2(new_n274), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(new_n275), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT88), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT88), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n292), .B(new_n288), .C1(new_n289), .C2(new_n275), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n207), .B1(new_n283), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n207), .B1(new_n291), .B2(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n286), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT89), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n283), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n297), .A2(new_n286), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n281), .A2(new_n282), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT89), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n296), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G197gat), .B(G204gat), .ZN(new_n306));
  INV_X1    g105(.A(G211gat), .ZN(new_n307));
  INV_X1    g106(.A(G218gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(KEYINPUT22), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G211gat), .B(G218gat), .Z(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G141gat), .B(G148gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  OR3_X1    g113(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT2), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n313), .A2(new_n317), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(new_n317), .B2(new_n313), .ZN(new_n323));
  XOR2_X1   g122(.A(G155gat), .B(G162gat), .Z(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n312), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n328), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n325), .B1(new_n330), .B2(new_n326), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(G22gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(G228gat), .A2(G233gat), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT77), .B1(new_n333), .B2(new_n334), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G78gat), .B(G106gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(new_n218), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n339), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n341), .A3(new_n336), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n340), .A2(new_n344), .A3(new_n342), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT25), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n350), .A2(G169gat), .A3(G176gat), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(G169gat), .B2(G176gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT66), .ZN(new_n353));
  NAND3_X1  g152(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n354), .A2(KEYINPUT67), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(KEYINPUT67), .ZN(new_n356));
  INV_X1    g155(.A(G183gat), .ZN(new_n357));
  INV_X1    g156(.A(G190gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT24), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(new_n357), .B2(new_n358), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n355), .A2(new_n356), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G169gat), .ZN(new_n363));
  INV_X1    g162(.A(G176gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n350), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n349), .B1(new_n353), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT27), .B(G183gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n358), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n370), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n371));
  OR4_X1    g170(.A1(KEYINPUT68), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT26), .B1(new_n365), .B2(KEYINPUT68), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n372), .B(new_n373), .C1(new_n363), .C2(new_n364), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n371), .B(new_n374), .C1(KEYINPUT28), .C2(new_n370), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n359), .A2(KEYINPUT65), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n359), .A2(KEYINPUT65), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n376), .A2(new_n354), .A3(new_n361), .A4(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n378), .A2(new_n349), .A3(new_n352), .A4(new_n366), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n368), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT69), .B(G113gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G120gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G127gat), .B(G134gat), .ZN(new_n384));
  INV_X1    g183(.A(G113gat), .ZN(new_n385));
  INV_X1    g184(.A(G120gat), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT1), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n388), .A2(KEYINPUT70), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n385), .B2(new_n386), .ZN(new_n390));
  INV_X1    g189(.A(new_n384), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n388), .A2(KEYINPUT70), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n381), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT64), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT34), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n400), .A2(KEYINPUT34), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n396), .A2(new_n399), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT33), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(G15gat), .B(G43gat), .Z(new_n406));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n401), .B(new_n402), .C1(new_n405), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n403), .A2(KEYINPUT32), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n402), .A2(new_n401), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n409), .B1(new_n403), .B2(new_n404), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n410), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n412), .B1(new_n410), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G226gat), .A2(G233gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n381), .A2(new_n419), .ZN(new_n420));
  OR2_X1    g219(.A1(new_n368), .A2(new_n380), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n328), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n423), .A2(new_n312), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n312), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n424), .A2(new_n429), .A3(new_n425), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(KEYINPUT30), .A3(new_n432), .ZN(new_n433));
  OR3_X1    g232(.A1(new_n426), .A2(KEYINPUT30), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n348), .A2(new_n418), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n394), .B2(new_n325), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT74), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n394), .A2(new_n437), .A3(new_n325), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(new_n438), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n440), .B1(new_n442), .B2(KEYINPUT74), .ZN(new_n443));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444));
  OR2_X1    g243(.A1(new_n325), .A2(new_n326), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(new_n395), .A3(new_n327), .ZN(new_n446));
  XOR2_X1   g245(.A(KEYINPUT73), .B(KEYINPUT5), .Z(new_n447));
  NAND4_X1  g246(.A1(new_n443), .A2(new_n444), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n394), .B(new_n325), .ZN(new_n449));
  INV_X1    g248(.A(new_n444), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n446), .A2(new_n444), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(new_n442), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G1gat), .B(G29gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT0), .ZN(new_n456));
  XNOR2_X1  g255(.A(G57gat), .B(G85gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT6), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n448), .A2(new_n458), .A3(new_n453), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT75), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(KEYINPUT75), .A3(new_n461), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n459), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT35), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n462), .A2(new_n466), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n348), .A2(new_n418), .A3(new_n435), .A4(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n436), .A2(new_n470), .B1(new_n472), .B2(new_n469), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n430), .B1(new_n426), .B2(KEYINPUT37), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n426), .A2(KEYINPUT37), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n474), .B2(KEYINPUT79), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n471), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n475), .A2(KEYINPUT79), .A3(new_n478), .A4(new_n476), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n432), .A4(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n435), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n443), .A2(new_n446), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n450), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n486), .A2(KEYINPUT39), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n486), .B(KEYINPUT39), .C1(new_n450), .C2(new_n449), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n458), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT78), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(KEYINPUT40), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n454), .A2(new_n459), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n489), .A2(new_n491), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n484), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n483), .A2(new_n495), .A3(new_n348), .ZN(new_n496));
  INV_X1    g295(.A(new_n348), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n468), .B2(new_n484), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(new_n416), .B2(new_n417), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n410), .A2(new_n415), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n411), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n410), .A2(new_n412), .A3(new_n415), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(KEYINPUT36), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n496), .A2(new_n498), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n305), .B1(new_n473), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G71gat), .B(G78gat), .ZN(new_n508));
  AND2_X1   g307(.A1(G57gat), .A2(G64gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(G57gat), .A2(G64gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n508), .B1(KEYINPUT9), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n514));
  AND2_X1   g313(.A1(G71gat), .A2(G78gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(KEYINPUT9), .ZN(new_n516));
  NAND2_X1  g315(.A1(G71gat), .A2(G78gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT9), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(KEYINPUT90), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n516), .A2(new_n511), .A3(new_n508), .A4(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT91), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n513), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT92), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G183gat), .B(G211gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n259), .B1(new_n524), .B2(new_n525), .ZN(new_n532));
  XNOR2_X1  g331(.A(G127gat), .B(G155gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n532), .B(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n531), .B(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT93), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(KEYINPUT41), .ZN(new_n540));
  XNOR2_X1  g339(.A(G134gat), .B(G162gat), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n540), .B(new_n541), .Z(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(G85gat), .A3(G92gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT94), .B1(G85gat), .B2(G92gat), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT96), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(KEYINPUT96), .A2(G99gat), .A3(G106gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(KEYINPUT8), .A3(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n554), .A2(new_n544), .A3(G85gat), .A4(G92gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n548), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n549), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n556), .B(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n559), .A2(new_n261), .B1(KEYINPUT41), .B2(new_n539), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT97), .Z(new_n561));
  XOR2_X1   g360(.A(G190gat), .B(G218gat), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n556), .A2(new_n549), .A3(new_n557), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n548), .A2(new_n553), .A3(new_n558), .A4(new_n555), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n279), .A2(new_n237), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n561), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n563), .B1(new_n561), .B2(new_n567), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n543), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n570), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(new_n542), .A3(new_n568), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n537), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G120gat), .B(G148gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT99), .ZN(new_n577));
  XOR2_X1   g376(.A(G176gat), .B(G204gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT100), .ZN(new_n581));
  NOR2_X1   g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n515), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n585), .A2(KEYINPUT91), .A3(new_n516), .A4(new_n519), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n520), .A2(new_n521), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n512), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n559), .A2(new_n588), .A3(KEYINPUT10), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n588), .B(new_n566), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n581), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n524), .A2(new_n566), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n559), .A2(new_n588), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n592), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n589), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(KEYINPUT100), .A3(new_n594), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603));
  OR3_X1    g402(.A1(new_n591), .A2(new_n603), .A3(new_n594), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n591), .B2(new_n594), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n580), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n604), .A2(new_n605), .A3(new_n580), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n593), .A2(new_n595), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT101), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n575), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n202), .B1(new_n507), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n507), .A2(new_n202), .A3(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n468), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g420(.A(KEYINPUT16), .B(G8gat), .Z(new_n622));
  INV_X1    g421(.A(new_n618), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n484), .B(new_n622), .C1(new_n623), .C2(new_n616), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n435), .B1(new_n617), .B2(new_n618), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n624), .B1(new_n625), .B2(new_n251), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT42), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT42), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(G1325gat));
  NOR2_X1   g429(.A1(new_n623), .A2(new_n616), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n505), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n500), .A2(new_n504), .A3(KEYINPUT103), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(G15gat), .B1(new_n631), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n619), .A2(new_n245), .A3(new_n418), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(G1326gat));
  XNOR2_X1  g438(.A(KEYINPUT43), .B(G22gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n619), .B2(new_n497), .ZN(new_n643));
  AOI211_X1 g442(.A(KEYINPUT104), .B(new_n348), .C1(new_n617), .C2(new_n618), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT104), .B1(new_n631), .B2(new_n348), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n619), .A2(new_n642), .A3(new_n497), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n647), .A3(new_n640), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(G1327gat));
  INV_X1    g448(.A(new_n537), .ZN(new_n650));
  INV_X1    g449(.A(new_n574), .ZN(new_n651));
  INV_X1    g450(.A(new_n614), .ZN(new_n652));
  AND4_X1   g451(.A1(new_n507), .A2(new_n650), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(new_n208), .A3(new_n468), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT45), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n473), .A2(new_n506), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n574), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n614), .B(KEYINPUT105), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n304), .A3(new_n650), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT106), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n633), .A2(new_n496), .A3(new_n498), .A4(new_n634), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n574), .B1(new_n664), .B2(new_n473), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n659), .B(new_n663), .C1(new_n665), .C2(KEYINPUT44), .ZN(new_n666));
  OAI21_X1  g465(.A(G29gat), .B1(new_n666), .B2(new_n467), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n655), .A2(new_n667), .ZN(G1328gat));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n209), .A3(new_n484), .ZN(new_n669));
  AND2_X1   g468(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n670));
  NOR2_X1   g469(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(G36gat), .B1(new_n666), .B2(new_n435), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n672), .B(new_n673), .C1(new_n670), .C2(new_n669), .ZN(G1329gat));
  INV_X1    g473(.A(new_n665), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n675), .A2(new_n657), .B1(new_n656), .B2(new_n658), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n676), .A2(new_n677), .A3(new_n635), .A4(new_n663), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT108), .B1(new_n666), .B2(new_n636), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n678), .A2(G43gat), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n653), .A2(new_n220), .A3(new_n418), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT47), .ZN(new_n682));
  OAI21_X1  g481(.A(G43gat), .B1(new_n666), .B2(new_n636), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(new_n681), .ZN(new_n684));
  OAI22_X1  g483(.A1(new_n680), .A2(new_n682), .B1(KEYINPUT47), .B2(new_n684), .ZN(G1330gat));
  OAI21_X1  g484(.A(G50gat), .B1(new_n666), .B2(new_n348), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n653), .A2(new_n218), .A3(new_n497), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT48), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n686), .A2(KEYINPUT48), .A3(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(G1331gat));
  NAND4_X1  g491(.A1(new_n660), .A2(new_n305), .A3(new_n537), .A4(new_n574), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n693), .B1(new_n664), .B2(new_n473), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n467), .B(KEYINPUT109), .Z(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g496(.A1(new_n694), .A2(new_n484), .ZN(new_n698));
  NOR2_X1   g497(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n699));
  AND2_X1   g498(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n698), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT110), .ZN(G1333gat));
  NAND2_X1  g502(.A1(new_n694), .A2(new_n635), .ZN(new_n704));
  INV_X1    g503(.A(new_n418), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(G71gat), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n704), .A2(G71gat), .B1(new_n694), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g507(.A1(new_n694), .A2(new_n497), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT111), .B(G78gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1335gat));
  NOR2_X1   g510(.A1(new_n537), .A2(new_n304), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n665), .A2(KEYINPUT51), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT51), .B1(new_n665), .B2(new_n712), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n467), .A2(G85gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n614), .A3(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n537), .A2(new_n304), .A3(new_n652), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n659), .B(new_n718), .C1(new_n665), .C2(KEYINPUT44), .ZN(new_n719));
  OAI21_X1  g518(.A(G85gat), .B1(new_n719), .B2(new_n467), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(G1336gat));
  NOR2_X1   g520(.A1(new_n435), .A2(G92gat), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n660), .B(new_n722), .C1(new_n713), .C2(new_n714), .ZN(new_n723));
  OAI21_X1  g522(.A(G92gat), .B1(new_n719), .B2(new_n435), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT52), .ZN(G1337gat));
  NOR2_X1   g525(.A1(new_n705), .A2(G99gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n715), .A2(new_n614), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G99gat), .B1(new_n719), .B2(new_n636), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1338gat));
  NOR2_X1   g529(.A1(new_n348), .A2(G106gat), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n660), .B(new_n731), .C1(new_n713), .C2(new_n714), .ZN(new_n732));
  OAI21_X1  g531(.A(G106gat), .B1(new_n719), .B2(new_n348), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g534(.A1(new_n537), .A2(new_n652), .A3(new_n305), .A4(new_n574), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT54), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n596), .A2(new_n737), .A3(new_n601), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n600), .B2(new_n594), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n599), .A2(new_n595), .A3(new_n589), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n580), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT55), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n574), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n610), .A2(new_n611), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n738), .A2(new_n741), .A3(KEYINPUT55), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT112), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n738), .A2(new_n741), .A3(new_n747), .A4(KEYINPUT55), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n744), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n299), .B1(new_n283), .B2(new_n298), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n301), .A2(KEYINPUT89), .A3(new_n302), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n268), .A2(new_n276), .A3(new_n280), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n289), .A2(new_n275), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n752), .A2(new_n269), .B1(new_n753), .B2(new_n288), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n750), .A2(new_n751), .B1(new_n206), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n743), .A2(new_n749), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n742), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n749), .A2(new_n304), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n613), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n607), .A2(new_n608), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n755), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n651), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n751), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n742), .B1(new_n766), .B2(new_n296), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n767), .A2(new_n749), .B1(new_n614), .B2(new_n755), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT113), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n757), .B1(new_n765), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n736), .B1(new_n770), .B2(new_n537), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(new_n695), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n418), .A3(new_n348), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n484), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n305), .A2(new_n382), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n467), .A2(new_n484), .ZN(new_n777));
  AND4_X1   g576(.A1(new_n418), .A2(new_n771), .A3(new_n348), .A4(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G113gat), .B1(new_n779), .B2(new_n305), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(KEYINPUT114), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(KEYINPUT114), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n776), .B1(new_n781), .B2(new_n782), .ZN(G1340gat));
  NAND2_X1  g582(.A1(new_n614), .A2(new_n386), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT115), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n774), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G120gat), .B1(new_n779), .B2(new_n661), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1341gat));
  AND3_X1   g587(.A1(new_n778), .A2(G127gat), .A3(new_n537), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n484), .A3(new_n650), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n790), .A2(KEYINPUT116), .ZN(new_n791));
  AOI21_X1  g590(.A(G127gat), .B1(new_n790), .B2(KEYINPUT116), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(G1342gat));
  NAND2_X1  g592(.A1(new_n435), .A2(new_n651), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n773), .A2(G134gat), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT56), .ZN(new_n796));
  OAI21_X1  g595(.A(G134gat), .B1(new_n779), .B2(new_n574), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT117), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(G1343gat));
  INV_X1    g598(.A(G141gat), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n635), .A2(new_n348), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n772), .A2(new_n801), .A3(new_n435), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n802), .B2(new_n305), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n636), .A2(new_n777), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n305), .A2(new_n800), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n651), .B1(new_n759), .B2(new_n762), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n650), .B1(new_n807), .B2(new_n757), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n736), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n348), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT118), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT57), .B1(new_n771), .B2(new_n497), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n805), .B(new_n806), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT119), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n803), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n816), .A2(KEYINPUT119), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n818), .B(new_n819), .ZN(G1344gat));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n348), .B1(new_n808), .B2(new_n736), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n821), .B1(new_n822), .B2(KEYINPUT57), .ZN(new_n823));
  INV_X1    g622(.A(new_n736), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n756), .B1(new_n768), .B2(new_n651), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n825), .B2(new_n650), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT120), .B(new_n810), .C1(new_n826), .C2(new_n348), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n771), .A2(new_n811), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(new_n614), .A3(new_n805), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n832));
  INV_X1    g631(.A(G148gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n614), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n813), .A2(new_n814), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n804), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n833), .B1(new_n836), .B2(new_n614), .ZN(new_n837));
  OAI221_X1 g636(.A(new_n832), .B1(new_n802), .B2(new_n834), .C1(new_n837), .C2(KEYINPUT59), .ZN(G1345gat));
  NOR3_X1   g637(.A1(new_n802), .A2(KEYINPUT121), .A3(new_n650), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n839), .A2(G155gat), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT121), .B1(new_n802), .B2(new_n650), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n537), .A2(G155gat), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n840), .A2(new_n841), .B1(new_n836), .B2(new_n842), .ZN(G1346gat));
  NAND2_X1  g642(.A1(new_n836), .A2(new_n651), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(G162gat), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n772), .A2(new_n801), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n794), .A2(G162gat), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(G1347gat));
  AND2_X1   g647(.A1(new_n771), .A2(new_n467), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n497), .A2(new_n705), .A3(new_n435), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n851), .A2(G169gat), .A3(new_n305), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT122), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n771), .A2(new_n348), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n695), .A2(new_n705), .A3(new_n435), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G169gat), .B1(new_n856), .B2(new_n305), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n853), .A2(new_n857), .ZN(G1348gat));
  OAI21_X1  g657(.A(G176gat), .B1(new_n856), .B2(new_n661), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n614), .A2(new_n364), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n851), .B2(new_n860), .ZN(G1349gat));
  OAI21_X1  g660(.A(G183gat), .B1(new_n856), .B2(new_n650), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n537), .A2(new_n369), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n851), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g664(.A1(new_n854), .A2(new_n651), .A3(new_n855), .ZN(new_n866));
  XNOR2_X1  g665(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n866), .A2(G190gat), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n866), .B2(G190gat), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n651), .A2(new_n358), .ZN(new_n870));
  OAI22_X1  g669(.A1(new_n868), .A2(new_n869), .B1(new_n851), .B2(new_n870), .ZN(G1351gat));
  NOR3_X1   g670(.A1(new_n635), .A2(new_n435), .A3(new_n348), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n849), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(G197gat), .A3(new_n305), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT124), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n874), .B(new_n875), .ZN(new_n876));
  OR3_X1    g675(.A1(new_n635), .A2(new_n435), .A3(new_n695), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n830), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n305), .ZN(new_n880));
  OAI21_X1  g679(.A(G197gat), .B1(new_n880), .B2(KEYINPUT125), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n880), .A2(KEYINPUT125), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n876), .B1(new_n881), .B2(new_n882), .ZN(G1352gat));
  OR3_X1    g682(.A1(new_n873), .A2(G204gat), .A3(new_n652), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(KEYINPUT126), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n885), .A2(KEYINPUT126), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(G204gat), .B1(new_n879), .B2(new_n661), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n888), .B(new_n889), .C1(new_n886), .C2(new_n884), .ZN(G1353gat));
  INV_X1    g689(.A(new_n873), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n307), .A3(new_n537), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n823), .A2(new_n827), .B1(new_n771), .B2(new_n811), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(new_n650), .A3(new_n877), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n307), .B1(new_n894), .B2(KEYINPUT127), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n877), .B1(new_n828), .B2(new_n829), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT127), .B1(new_n896), .B2(new_n537), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT63), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n830), .A2(KEYINPUT127), .A3(new_n537), .A4(new_n878), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G211gat), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(new_n897), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n892), .B1(new_n899), .B2(new_n903), .ZN(G1354gat));
  OAI21_X1  g703(.A(G218gat), .B1(new_n879), .B2(new_n574), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n891), .A2(new_n308), .A3(new_n651), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1355gat));
endmodule


