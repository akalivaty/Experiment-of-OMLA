//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1226, new_n1227, new_n1228, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n214), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT64), .Z(new_n223));
  AOI22_X1  g0023(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G87), .ZN(new_n227));
  INV_X1    g0027(.A(G250), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  INV_X1    g0031(.A(G238), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n230), .B1(new_n202), .B2(new_n231), .C1(new_n203), .C2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n210), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT1), .Z(new_n235));
  NAND2_X1  g0035(.A1(new_n223), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n231), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n256));
  AND3_X1   g0056(.A1(new_n254), .A2(KEYINPUT66), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT66), .B1(new_n254), .B2(new_n256), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G226), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(new_n254), .A3(G274), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n254), .B1(new_n267), .B2(new_n225), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G222), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n269), .B1(new_n270), .B2(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  OR2_X1    g0072(.A1(KEYINPUT67), .A2(G223), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT67), .A2(G223), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n268), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n260), .A2(new_n264), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G179), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT69), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(G20), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n218), .A2(KEYINPUT69), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n282), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n290), .A2(new_n291), .A3(new_n217), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n290), .B2(new_n217), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G13), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n295), .A2(new_n218), .A3(G1), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n289), .A2(new_n294), .B1(new_n201), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n294), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(G1), .B2(new_n218), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n297), .B1(new_n299), .B2(new_n201), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n280), .B(new_n300), .C1(G169), .C2(new_n278), .ZN(new_n301));
  INV_X1    g0101(.A(G200), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n276), .A2(new_n264), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n260), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(G190), .B2(new_n278), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n300), .A2(KEYINPUT9), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n297), .B(new_n308), .C1(new_n299), .C2(new_n201), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n306), .B1(new_n305), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n301), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT16), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT7), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n269), .B2(G20), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n218), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n203), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n202), .A2(new_n203), .ZN(new_n321));
  NOR2_X1   g0121(.A1(G58), .A2(G68), .ZN(new_n322));
  OAI21_X1  g0122(.A(G20), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n281), .A2(G159), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n316), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT7), .B1(new_n267), .B2(new_n218), .ZN(new_n327));
  NOR4_X1   g0127(.A1(new_n265), .A2(new_n266), .A3(new_n317), .A4(G20), .ZN(new_n328));
  OAI21_X1  g0128(.A(G68), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n325), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(KEYINPUT16), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n326), .A2(new_n331), .A3(new_n294), .ZN(new_n332));
  INV_X1    g0132(.A(new_n288), .ZN(new_n333));
  INV_X1    g0133(.A(new_n296), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n294), .B1(new_n255), .B2(G20), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n333), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n254), .A2(new_n256), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n264), .B1(new_n231), .B2(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(G226), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT75), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n284), .A2(new_n227), .ZN(new_n342));
  INV_X1    g0142(.A(G223), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(G1698), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n269), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT75), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n269), .A2(new_n346), .A3(G226), .A4(G1698), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n341), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n254), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n339), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(G200), .ZN(new_n351));
  AOI211_X1 g0151(.A(G190), .B(new_n339), .C1(new_n348), .C2(new_n349), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n332), .B(new_n337), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT17), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n335), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n299), .B2(new_n288), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n329), .A2(new_n330), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n298), .B1(new_n358), .B2(new_n316), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n357), .B1(new_n359), .B2(new_n331), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n350), .A2(new_n279), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(G169), .B2(new_n350), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT18), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n332), .A2(new_n337), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n348), .A2(new_n349), .ZN(new_n365));
  INV_X1    g0165(.A(new_n339), .ZN(new_n366));
  AOI21_X1  g0166(.A(G169), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI211_X1 g0167(.A(G179), .B(new_n339), .C1(new_n348), .C2(new_n349), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT18), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n364), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n363), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n355), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n336), .A2(G77), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT70), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n288), .B(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n281), .ZN(new_n378));
  INV_X1    g0178(.A(new_n287), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT15), .B(G87), .Z(new_n380));
  AOI22_X1  g0180(.A1(new_n379), .A2(new_n380), .B1(G20), .B2(G77), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n298), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n334), .A2(G77), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n375), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G169), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G238), .A2(G1698), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n269), .B(new_n386), .C1(new_n231), .C2(G1698), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(new_n349), .C1(G107), .C2(new_n269), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n264), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n257), .A2(new_n258), .A3(new_n226), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n390), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n392), .A2(new_n279), .A3(new_n388), .A4(new_n264), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n384), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G200), .B1(new_n389), .B2(new_n390), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n392), .A2(G190), .A3(new_n388), .A4(new_n264), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n384), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(new_n399), .A3(KEYINPUT71), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n396), .A2(new_n399), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT71), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n315), .A2(new_n373), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n287), .A2(new_n225), .B1(new_n218), .B2(G68), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n405), .A2(KEYINPUT74), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n405), .A2(KEYINPUT74), .B1(G50), .B2(new_n281), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n298), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT11), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n296), .A2(new_n203), .ZN(new_n410));
  XOR2_X1   g0210(.A(new_n410), .B(KEYINPUT12), .Z(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(G68), .B2(new_n336), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n408), .A2(KEYINPUT11), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT14), .ZN(new_n417));
  OAI211_X1 g0217(.A(G226), .B(new_n272), .C1(new_n265), .C2(new_n266), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT72), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G97), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT73), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT73), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(G33), .A3(G97), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n269), .A2(G232), .A3(G1698), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n420), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n418), .A2(new_n419), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n349), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  INV_X1    g0230(.A(new_n264), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n259), .B2(G238), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n430), .B1(new_n429), .B2(new_n432), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n417), .B(G169), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n429), .A2(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT13), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n435), .B1(new_n279), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n417), .B1(new_n439), .B2(G169), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n416), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(G200), .ZN(new_n443));
  INV_X1    g0243(.A(G190), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n415), .B(new_n443), .C1(new_n444), .C2(new_n439), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n404), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n295), .A2(G1), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n448), .A2(G20), .B1(new_n255), .B2(G33), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n292), .B2(new_n293), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT77), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT77), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n449), .B(new_n452), .C1(new_n292), .C2(new_n293), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(G97), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n296), .A2(new_n206), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n207), .B1(new_n318), .B2(new_n319), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT6), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G97), .A2(G107), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n208), .A2(KEYINPUT76), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(KEYINPUT76), .ZN(new_n460));
  AND2_X1   g0260(.A1(G97), .A2(G107), .ZN(new_n461));
  NOR2_X1   g0261(.A1(G97), .A2(G107), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n464));
  AND4_X1   g0264(.A1(G20), .A2(new_n459), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n225), .A2(G20), .A3(G33), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n456), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n454), .B(new_n455), .C1(new_n467), .C2(new_n298), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  OR2_X1    g0269(.A1(KEYINPUT3), .A2(G33), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT3), .A2(G33), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n226), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT78), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(KEYINPUT4), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n469), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(G250), .B1(new_n265), .B2(new_n266), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n272), .B1(new_n477), .B2(new_n475), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(G244), .B1(new_n265), .B2(new_n266), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT78), .B1(new_n480), .B2(G1698), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n254), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n262), .A2(G1), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G41), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(G274), .A3(new_n254), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n254), .ZN(new_n491));
  INV_X1    g0291(.A(G257), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n385), .B1(new_n483), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n228), .B1(new_n470), .B2(new_n471), .ZN(new_n495));
  OAI21_X1  g0295(.A(G1698), .B1(new_n495), .B2(new_n474), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n480), .A2(new_n474), .B1(G33), .B2(G283), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n473), .B1(new_n472), .B2(new_n272), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n496), .B(new_n497), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n493), .B1(new_n500), .B2(new_n349), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n279), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n468), .A2(new_n494), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(new_n349), .ZN(new_n504));
  INV_X1    g0304(.A(new_n493), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT80), .B1(new_n506), .B2(new_n444), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT80), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n501), .A2(new_n508), .A3(G190), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT79), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n501), .B2(new_n302), .ZN(new_n512));
  OAI211_X1 g0312(.A(KEYINPUT79), .B(G200), .C1(new_n483), .C2(new_n493), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n468), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n503), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n451), .A2(G107), .A3(new_n453), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n296), .B(new_n207), .C1(new_n517), .C2(KEYINPUT25), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(KEYINPUT25), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n218), .B(G87), .C1(new_n265), .C2(new_n266), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT22), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT22), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n269), .A2(new_n525), .A3(new_n218), .A4(G87), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT24), .ZN(new_n528));
  INV_X1    g0328(.A(G116), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n284), .A2(new_n529), .A3(G20), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT84), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n218), .B2(G107), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT23), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n531), .B(new_n534), .C1(new_n218), .C2(G107), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n530), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n527), .A2(new_n528), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n528), .B1(new_n527), .B2(new_n536), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n294), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G257), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n541), .B(new_n542), .C1(new_n477), .C2(G1698), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n349), .ZN(new_n544));
  INV_X1    g0344(.A(new_n491), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G264), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n546), .A3(new_n489), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(G190), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n349), .A2(new_n543), .B1(new_n545), .B2(G264), .ZN(new_n549));
  AOI21_X1  g0349(.A(G200), .B1(new_n549), .B2(new_n489), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n522), .B(new_n540), .C1(new_n548), .C2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n334), .A2(new_n380), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n285), .A2(G97), .A3(new_n286), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT82), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n422), .A2(new_n424), .A3(KEYINPUT19), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n218), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n227), .A2(new_n206), .A3(new_n207), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n269), .A2(new_n218), .A3(G68), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT82), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n553), .A2(new_n562), .A3(new_n554), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n556), .A2(new_n560), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n552), .B1(new_n564), .B2(new_n294), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n451), .A2(new_n380), .A3(new_n453), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n226), .A2(G1698), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G238), .B2(G1698), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n569), .A2(new_n267), .B1(new_n284), .B2(new_n529), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n349), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n228), .B1(new_n255), .B2(G45), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n254), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT81), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n254), .A3(KEYINPUT81), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n254), .A2(G274), .A3(new_n484), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n571), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(G179), .ZN(new_n580));
  INV_X1    g0380(.A(G274), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n349), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n570), .A2(new_n349), .B1(new_n582), .B2(new_n484), .ZN(new_n583));
  AOI21_X1  g0383(.A(G169), .B1(new_n583), .B2(new_n577), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n567), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n284), .A2(new_n529), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G238), .A2(G1698), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n226), .B2(G1698), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n587), .B1(new_n589), .B2(new_n269), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n578), .B1(new_n590), .B2(new_n254), .ZN(new_n591));
  INV_X1    g0391(.A(new_n576), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT81), .B1(new_n572), .B2(new_n254), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n302), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n583), .A2(new_n444), .A3(new_n577), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n451), .A2(G87), .A3(new_n453), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n565), .A3(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n551), .A2(new_n586), .A3(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n449), .B(G116), .C1(new_n292), .C2(new_n293), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n296), .A2(new_n529), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n290), .A2(new_n217), .B1(G20), .B2(new_n529), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n469), .B(new_n218), .C1(G33), .C2(new_n206), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT20), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n603), .A2(KEYINPUT20), .A3(new_n604), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n601), .B(new_n602), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n272), .A2(G257), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G264), .A2(G1698), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n608), .B(new_n609), .C1(new_n265), .C2(new_n266), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n610), .B(new_n349), .C1(G303), .C2(new_n269), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n490), .A2(G270), .A3(new_n254), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n489), .A3(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n613), .A2(KEYINPUT21), .A3(G169), .ZN(new_n614));
  AND4_X1   g0414(.A1(G179), .A2(new_n611), .A3(new_n489), .A4(new_n612), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n607), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n607), .A2(G169), .A3(new_n613), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT83), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n618), .B1(new_n617), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n616), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n547), .A2(new_n385), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n549), .A2(new_n279), .A3(new_n489), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n527), .A2(new_n536), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT24), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n298), .B1(new_n626), .B2(new_n537), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n623), .B(new_n624), .C1(new_n627), .C2(new_n521), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n613), .A2(new_n444), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n607), .B(new_n630), .C1(G200), .C2(new_n613), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n622), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n447), .A2(new_n515), .A3(new_n600), .A4(new_n632), .ZN(G372));
  OAI211_X1 g0433(.A(new_n628), .B(new_n616), .C1(new_n621), .C2(new_n620), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n514), .A2(new_n510), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n468), .A2(new_n502), .A3(new_n494), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n600), .A2(new_n634), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n564), .A2(new_n294), .ZN(new_n639));
  INV_X1    g0439(.A(new_n552), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n639), .A2(new_n640), .A3(new_n566), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n579), .A2(new_n385), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(G179), .B2(new_n579), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n599), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n638), .B1(new_n644), .B2(new_n636), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n503), .A2(KEYINPUT26), .A3(new_n586), .A4(new_n599), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n637), .A2(new_n647), .A3(new_n586), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n447), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n301), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n364), .A2(new_n369), .A3(new_n370), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n370), .B1(new_n364), .B2(new_n369), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n440), .A2(new_n441), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(new_n416), .B1(new_n445), .B2(new_n395), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n653), .B1(new_n655), .B2(new_n355), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n305), .A2(new_n310), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT10), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n311), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n650), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n649), .A2(new_n660), .ZN(G369));
  INV_X1    g0461(.A(KEYINPUT86), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n448), .A2(new_n218), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(new_n607), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n622), .A2(new_n662), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n662), .B1(new_n622), .B2(new_n669), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n631), .A2(new_n669), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n670), .A2(new_n671), .B1(new_n622), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G330), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n668), .B1(new_n627), .B2(new_n521), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n551), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n628), .ZN(new_n677));
  INV_X1    g0477(.A(new_n668), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n629), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n622), .A2(new_n678), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n684), .B1(new_n629), .B2(new_n678), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n682), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n211), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n559), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n215), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  INV_X1    g0493(.A(new_n586), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n645), .B2(new_n646), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n668), .B1(new_n695), .B2(new_n637), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT29), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n613), .A2(new_n279), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(KEYINPUT88), .B2(new_n579), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n579), .A2(KEYINPUT88), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n702), .A2(new_n506), .A3(new_n547), .A4(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(KEYINPUT87), .A2(KEYINPUT30), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n591), .A2(new_n594), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(new_n615), .A3(new_n549), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n705), .B1(new_n707), .B2(new_n506), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n706), .A2(new_n549), .ZN(new_n709));
  INV_X1    g0509(.A(new_n705), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n501), .A3(new_n615), .A4(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n704), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT31), .B1(new_n712), .B2(new_n668), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n632), .A2(new_n515), .A3(new_n600), .A4(new_n678), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n700), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n699), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n693), .B1(new_n720), .B2(G1), .ZN(G364));
  NOR2_X1   g0521(.A1(new_n295), .A2(G20), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G45), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n689), .A2(G1), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n674), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n673), .A2(G330), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n673), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n724), .B(KEYINPUT89), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n218), .A2(G190), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G179), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G159), .ZN(new_n738));
  OR3_X1    g0538(.A1(new_n737), .A2(KEYINPUT32), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n218), .A2(G179), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n444), .A3(G200), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G107), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G87), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT32), .B1(new_n737), .B2(new_n738), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n739), .A2(new_n743), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n279), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n735), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n218), .A2(new_n279), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n444), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n269), .B1(new_n750), .B2(new_n225), .C1(new_n754), .C2(new_n201), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n749), .A2(G20), .A3(G190), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT91), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n748), .B(new_n755), .C1(G58), .C2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n751), .A2(new_n444), .A3(G200), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n218), .B1(new_n736), .B2(G190), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n203), .B1(new_n761), .B2(new_n206), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT92), .ZN(new_n763));
  INV_X1    g0563(.A(G326), .ZN(new_n764));
  INV_X1    g0564(.A(G294), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n754), .A2(new_n764), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  INV_X1    g0567(.A(G303), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n767), .A2(new_n741), .B1(new_n744), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G322), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n267), .B1(new_n756), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  INV_X1    g0573(.A(G329), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n750), .A2(new_n773), .B1(new_n737), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT33), .B(G317), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT93), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n760), .B1(new_n777), .B2(KEYINPUT93), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n772), .B(new_n775), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n759), .A2(new_n763), .B1(new_n770), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n217), .B1(G20), .B2(new_n385), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n730), .A2(new_n782), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n687), .A2(new_n267), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n786), .A2(G355), .B1(new_n529), .B2(new_n687), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n687), .A2(new_n269), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT90), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(G45), .B2(new_n215), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n251), .A2(new_n262), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n734), .B(new_n784), .C1(new_n785), .C2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n727), .B1(new_n732), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  AND2_X1   g0595(.A1(new_n391), .A2(new_n393), .ZN(new_n796));
  INV_X1    g0596(.A(new_n383), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n378), .A2(new_n381), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n374), .B(new_n797), .C1(new_n798), .C2(new_n298), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n796), .A2(KEYINPUT95), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT95), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n384), .B2(new_n394), .ZN(new_n802));
  AND3_X1   g0602(.A1(new_n800), .A2(new_n802), .A3(new_n399), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n648), .A2(new_n678), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n799), .A2(new_n668), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n803), .A2(new_n805), .B1(new_n395), .B2(new_n668), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n804), .B1(new_n696), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n718), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT96), .Z(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n808), .A2(new_n718), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT97), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n812), .A2(KEYINPUT97), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n811), .A2(new_n724), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n782), .A2(new_n728), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n734), .B1(new_n225), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n760), .ZN(new_n818));
  INV_X1    g0618(.A(new_n750), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(G150), .B1(new_n819), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  INV_X1    g0621(.A(G143), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n754), .B2(new_n821), .C1(new_n757), .C2(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT34), .Z(new_n824));
  NAND2_X1  g0624(.A1(new_n742), .A2(G68), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n825), .B(new_n269), .C1(new_n826), .C2(new_n737), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n744), .A2(new_n201), .B1(new_n761), .B2(new_n202), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n824), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n756), .A2(new_n765), .B1(new_n761), .B2(new_n206), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT94), .Z(new_n831));
  OAI221_X1 g0631(.A(new_n267), .B1(new_n737), .B2(new_n773), .C1(new_n529), .C2(new_n750), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n227), .A2(new_n741), .B1(new_n744), .B2(new_n207), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n754), .A2(new_n768), .B1(new_n767), .B2(new_n760), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n831), .A2(new_n832), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n829), .A2(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n817), .B1(new_n783), .B2(new_n836), .C1(new_n807), .C2(new_n729), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n815), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G384));
  INV_X1    g0639(.A(KEYINPUT40), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT38), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n360), .A2(new_n666), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n360), .B(new_n354), .C1(new_n352), .C2(new_n351), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n353), .A2(KEYINPUT17), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n843), .B1(new_n653), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n666), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n364), .B1(new_n369), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n849), .A2(new_n850), .A3(new_n353), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n849), .B2(new_n353), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n841), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT98), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n842), .B1(new_n355), .B2(new_n372), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n849), .A2(new_n353), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n849), .A2(new_n850), .A3(new_n353), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n856), .A2(KEYINPUT38), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n854), .A2(new_n855), .A3(new_n861), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n856), .A2(new_n860), .A3(KEYINPUT98), .A4(KEYINPUT38), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n415), .A2(new_n678), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n442), .A2(new_n445), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n654), .A2(new_n864), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n806), .B1(new_n716), .B2(new_n715), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n862), .A2(new_n863), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n849), .A2(KEYINPUT99), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n857), .A2(new_n871), .A3(KEYINPUT37), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT100), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n849), .B(new_n353), .C1(KEYINPUT99), .C2(new_n850), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n875), .A2(new_n876), .A3(new_n847), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n861), .B1(new_n877), .B2(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n715), .A2(new_n716), .ZN(new_n879));
  AND4_X1   g0679(.A1(KEYINPUT40), .A2(new_n879), .A3(new_n868), .A4(new_n807), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n840), .A2(new_n870), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n447), .A2(new_n879), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT101), .ZN(new_n884));
  OAI21_X1  g0684(.A(G330), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n882), .B2(new_n884), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n654), .A2(new_n416), .A3(new_n678), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n888), .B(new_n861), .C1(new_n877), .C2(KEYINPUT38), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n862), .A2(KEYINPUT39), .A3(new_n863), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n668), .B1(new_n800), .B2(new_n802), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n804), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n868), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n862), .A2(new_n863), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n895), .A2(new_n896), .B1(new_n653), .B2(new_n848), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n697), .A2(new_n447), .A3(new_n698), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n660), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n898), .B(new_n900), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n886), .A2(new_n901), .B1(new_n255), .B2(new_n722), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n901), .B2(new_n886), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n459), .A2(new_n463), .A3(new_n464), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT35), .ZN(new_n905));
  OAI211_X1 g0705(.A(G116), .B(new_n219), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n905), .B2(new_n904), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT36), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n216), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n201), .A2(G68), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n255), .B(G13), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  OR3_X1    g0711(.A1(new_n903), .A2(new_n908), .A3(new_n911), .ZN(G367));
  AOI21_X1  g0712(.A(new_n678), .B1(new_n565), .B2(new_n598), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT102), .Z(new_n914));
  OR2_X1    g0714(.A1(new_n914), .A2(new_n644), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n694), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n730), .ZN(new_n918));
  INV_X1    g0718(.A(new_n380), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n785), .B1(new_n211), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n789), .B2(new_n244), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n269), .B1(new_n741), .B2(new_n225), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT108), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n750), .A2(new_n201), .B1(new_n737), .B2(new_n821), .ZN(new_n924));
  INV_X1    g0724(.A(new_n756), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(G150), .B2(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n753), .A2(G143), .B1(new_n745), .B2(G58), .ZN(new_n927));
  INV_X1    g0727(.A(new_n761), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n818), .A2(G159), .B1(new_n928), .B2(G68), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n923), .A2(new_n926), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT46), .B1(new_n745), .B2(G116), .ZN(new_n931));
  XNOR2_X1  g0731(.A(KEYINPUT107), .B(G317), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n737), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n267), .B1(new_n750), .B2(new_n767), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n768), .B2(new_n757), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n745), .A2(KEYINPUT46), .A3(G116), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT106), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n753), .A2(G311), .B1(new_n742), .B2(G97), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n818), .A2(G294), .B1(new_n928), .B2(G107), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n930), .B1(new_n936), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT47), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n734), .B(new_n921), .C1(new_n945), .C2(new_n782), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n918), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n688), .B(KEYINPUT41), .Z(new_n948));
  INV_X1    g0748(.A(new_n680), .ZN(new_n949));
  INV_X1    g0749(.A(new_n683), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT104), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(new_n673), .A3(G330), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n949), .A2(new_n950), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n674), .A2(KEYINPUT104), .A3(new_n951), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n953), .B2(new_n955), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n719), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n468), .A2(new_n668), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n515), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n503), .A2(new_n668), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n685), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT45), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT44), .B1(new_n685), .B2(new_n963), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n685), .A2(KEYINPUT44), .A3(new_n963), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n966), .A2(new_n682), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n964), .B(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n967), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n681), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n959), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n948), .B1(new_n973), .B2(new_n720), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n723), .A2(G1), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT105), .Z(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n963), .A2(new_n684), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n515), .A2(new_n629), .A3(new_n960), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n668), .B1(new_n981), .B2(new_n636), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n979), .B2(KEYINPUT42), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n917), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n917), .A2(new_n985), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n980), .A2(new_n983), .A3(new_n985), .A4(new_n917), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n963), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n990), .A2(new_n682), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n990), .B1(new_n682), .B2(new_n991), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n992), .B1(KEYINPUT103), .B2(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(KEYINPUT103), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n947), .B1(new_n978), .B2(new_n996), .ZN(G387));
  INV_X1    g0797(.A(new_n958), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n977), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT109), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n818), .A2(G311), .B1(new_n819), .B2(G303), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n754), .B2(new_n771), .C1(new_n757), .C2(new_n932), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT48), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n745), .A2(G294), .B1(new_n928), .B2(G283), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT49), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n267), .B1(new_n737), .B2(new_n764), .C1(new_n529), .C2(new_n741), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n756), .A2(new_n201), .B1(new_n750), .B2(new_n203), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n737), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n267), .B(new_n1013), .C1(G150), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n928), .A2(new_n380), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G159), .A2(new_n753), .B1(new_n818), .B2(new_n333), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n745), .A2(G77), .B1(new_n742), .B2(G97), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n783), .B1(new_n1012), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n241), .A2(G45), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n377), .A2(new_n201), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT50), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n690), .B(new_n262), .C1(new_n203), .C2(new_n225), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n789), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n786), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1025), .B1(G107), .B2(new_n211), .C1(new_n690), .C2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n734), .B(new_n1020), .C1(new_n785), .C2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n949), .B2(new_n731), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT110), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n959), .A2(new_n689), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n720), .B2(new_n998), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1000), .A2(new_n1030), .A3(new_n1032), .ZN(G393));
  NAND3_X1  g0833(.A1(new_n972), .A2(new_n969), .A3(KEYINPUT111), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT111), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n681), .C1(new_n970), .C2(new_n971), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n688), .B(new_n973), .C1(new_n1037), .C2(new_n959), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n789), .A2(new_n248), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n785), .B1(new_n206), .B2(new_n211), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n743), .B(new_n267), .C1(new_n771), .C2(new_n737), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n818), .A2(G303), .B1(new_n819), .B2(G294), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n529), .B2(new_n761), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT113), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1041), .B(new_n1044), .C1(G283), .C2(new_n745), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n753), .A2(G317), .B1(new_n925), .B2(G311), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT112), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT52), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n753), .A2(G150), .B1(new_n925), .B2(G159), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT51), .Z(new_n1050));
  OAI221_X1 g0850(.A(new_n269), .B1(new_n737), .B2(new_n822), .C1(new_n227), .C2(new_n741), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n928), .A2(G77), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n201), .B2(new_n760), .C1(new_n203), .C2(new_n744), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(new_n377), .C2(new_n819), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1045), .A2(new_n1048), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n733), .B1(new_n1039), .B2(new_n1040), .C1(new_n1055), .C2(new_n783), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n730), .B2(new_n991), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n1037), .B2(new_n977), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1038), .A2(new_n1058), .ZN(G390));
  INV_X1    g0859(.A(KEYINPUT114), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n800), .A2(new_n802), .A3(new_n399), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n668), .B(new_n1061), .C1(new_n695), .C2(new_n637), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1060), .B1(new_n1062), .B2(new_n892), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n804), .A2(new_n893), .A3(KEYINPUT114), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n868), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n887), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n872), .A2(new_n874), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(KEYINPUT100), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n856), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n841), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1066), .B1(new_n1071), .B2(new_n861), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1065), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n892), .B1(new_n696), .B2(new_n803), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n868), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n887), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n889), .A3(new_n890), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n717), .A2(new_n807), .A3(new_n868), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1073), .A2(new_n1079), .A3(new_n1077), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(KEYINPUT116), .B1(new_n1083), .B2(new_n976), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1073), .A2(new_n1079), .A3(new_n1077), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1079), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT116), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n1088), .A3(new_n977), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n889), .A2(new_n728), .A3(new_n890), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n816), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n733), .B1(new_n333), .B2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n742), .A2(G50), .B1(new_n928), .B2(G159), .ZN(new_n1093));
  INV_X1    g0893(.A(G128), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1093), .B1(new_n821), .B2(new_n760), .C1(new_n1094), .C2(new_n754), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT54), .B(G143), .ZN(new_n1096));
  INV_X1    g0896(.A(G125), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n750), .A2(new_n1096), .B1(new_n737), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n267), .B1(new_n925), .B2(G132), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n1101));
  INV_X1    g0901(.A(G150), .ZN(new_n1102));
  OR3_X1    g0902(.A1(new_n744), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1101), .B1(new_n744), .B2(new_n1102), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1099), .A2(new_n1100), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1052), .B1(new_n207), .B2(new_n760), .C1(new_n754), .C2(new_n767), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n925), .A2(G116), .B1(new_n1014), .B2(G294), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n269), .B1(new_n819), .B2(G97), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1107), .A2(new_n746), .A3(new_n825), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1095), .A2(new_n1105), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1092), .B1(new_n1110), .B2(new_n782), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1084), .A2(new_n1089), .B1(new_n1090), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n447), .A2(new_n717), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n899), .A2(new_n660), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1075), .B1(new_n718), .B2(new_n806), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1079), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n894), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n1115), .A3(new_n1079), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1114), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n689), .B1(new_n1083), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT115), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n1087), .B2(new_n1120), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1081), .A2(new_n1120), .A3(new_n1123), .A4(new_n1082), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1122), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1112), .A2(new_n1127), .ZN(G378));
  OR2_X1    g0928(.A1(new_n891), .A2(new_n897), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n300), .A2(new_n848), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n314), .A2(KEYINPUT121), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT121), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n659), .A2(new_n1132), .A3(new_n301), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1131), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1130), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n1134), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1130), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1131), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n881), .B2(G330), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n870), .A2(new_n840), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n878), .A2(new_n880), .ZN(new_n1147));
  AND4_X1   g0947(.A1(G330), .A2(new_n1146), .A3(new_n1147), .A4(new_n1144), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1129), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1146), .A2(new_n1147), .A3(G330), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1144), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n881), .A2(G330), .A3(new_n1144), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n1153), .A3(new_n898), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1149), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n977), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n753), .A2(G125), .B1(G150), .B2(new_n928), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT119), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n756), .A2(new_n1094), .B1(new_n750), .B2(new_n821), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1096), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1159), .B1(new_n745), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1158), .B(new_n1161), .C1(new_n826), .C2(new_n760), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  AOI211_X1 g0963(.A(G33), .B(G41), .C1(new_n1014), .C2(G124), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n738), .C2(new_n741), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n925), .A2(G107), .B1(new_n1014), .B2(G283), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n919), .B2(new_n750), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n261), .B(new_n267), .C1(new_n744), .C2(new_n225), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT118), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n760), .A2(new_n206), .B1(new_n761), .B2(new_n203), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n754), .A2(new_n529), .B1(new_n741), .B2(new_n202), .ZN(new_n1173));
  OR4_X1    g0973(.A1(new_n1169), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT58), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n201), .B1(new_n265), .B2(G41), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n782), .B1(new_n1167), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT120), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n724), .B1(new_n201), .B2(new_n816), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n1144), .C2(new_n729), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1156), .A2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1114), .B(KEYINPUT122), .Z(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1186), .B2(new_n1155), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1185), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1081), .A2(new_n1120), .A3(new_n1082), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT115), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1188), .B1(new_n1190), .B2(new_n1125), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT123), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1149), .A2(new_n1192), .A3(new_n1154), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1152), .A2(new_n1153), .A3(new_n898), .A4(KEYINPUT123), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(KEYINPUT57), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n688), .B1(new_n1191), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1184), .B1(new_n1187), .B2(new_n1196), .ZN(G375));
  AND2_X1   g0997(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(new_n976), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G116), .A2(new_n818), .B1(new_n745), .B2(G97), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n765), .B2(new_n754), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n267), .B1(new_n737), .B2(new_n768), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n756), .A2(new_n767), .B1(new_n750), .B2(new_n207), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1016), .B1(new_n225), .B2(new_n741), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n269), .B1(new_n737), .B2(new_n1094), .C1(new_n1102), .C2(new_n750), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n818), .A2(new_n1160), .B1(new_n928), .B2(G50), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n202), .B2(new_n741), .C1(new_n738), .C2(new_n744), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1206), .B(new_n1208), .C1(G137), .C2(new_n758), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n753), .A2(G132), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT124), .Z(new_n1211));
  AOI21_X1  g1011(.A(new_n1205), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n733), .B1(G68), .B2(new_n1091), .C1(new_n1212), .C2(new_n783), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1075), .B2(new_n728), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1199), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1198), .A2(new_n1114), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n948), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1217), .A3(new_n1121), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1218), .ZN(G381));
  OR2_X1    g1019(.A1(G393), .A2(G396), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1220), .A2(G384), .A3(G390), .A4(G381), .ZN(new_n1221));
  INV_X1    g1021(.A(G387), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1112), .A2(new_n1127), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n1224), .A2(G375), .ZN(G407));
  NAND2_X1  g1025(.A1(new_n667), .A2(G213), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1223), .A2(new_n1227), .ZN(new_n1228));
  OAI211_X1 g1028(.A(G407), .B(G213), .C1(G375), .C2(new_n1228), .ZN(G409));
  NAND3_X1  g1029(.A1(G387), .A2(new_n1038), .A3(new_n1058), .ZN(new_n1230));
  OAI211_X1 g1030(.A(G390), .B(new_n947), .C1(new_n978), .C2(new_n996), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G393), .A2(G396), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1220), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT126), .B1(new_n1222), .B2(G390), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1232), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(KEYINPUT126), .A3(new_n1231), .A4(new_n1230), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(G378), .B(new_n1184), .C1(new_n1187), .C2(new_n1196), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1155), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1191), .A2(new_n948), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1193), .A2(new_n977), .A3(new_n1194), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1183), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1223), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1227), .B1(new_n1240), .B2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1198), .A2(KEYINPUT60), .A3(new_n1114), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(new_n688), .A3(new_n1121), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT60), .B1(new_n1198), .B2(new_n1114), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1215), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1250), .A2(new_n838), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n838), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1246), .A2(KEYINPUT125), .A3(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT125), .B1(new_n1246), .B2(new_n1254), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1255), .A2(new_n1256), .A3(KEYINPUT62), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1240), .A2(new_n1245), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1226), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1227), .A2(G2897), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1253), .B(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT62), .B1(new_n1259), .B2(new_n1253), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1239), .B1(new_n1257), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1246), .A2(KEYINPUT63), .A3(new_n1254), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1262), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1265), .A2(new_n1270), .ZN(G405));
  NAND2_X1  g1071(.A1(G375), .A2(new_n1223), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1253), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(G375), .A2(new_n1223), .A3(new_n1254), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1239), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1240), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1277), .A2(KEYINPUT127), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1268), .A2(new_n1274), .A3(new_n1273), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1276), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1278), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(G402));
endmodule


