//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G22gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(G228gat), .A2(G233gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G141gat), .B(G148gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n209), .B(new_n212), .C1(new_n213), .C2(KEYINPUT2), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(G148gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n209), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n214), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT74), .B(G197gat), .Z(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G204gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT74), .B(G197gat), .ZN(new_n226));
  INV_X1    g025(.A(G204gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(G211gat), .B(G218gat), .Z(new_n233));
  INV_X1    g032(.A(KEYINPUT76), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT75), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n230), .B1(new_n225), .B2(new_n228), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n234), .B1(new_n238), .B2(KEYINPUT75), .ZN(new_n239));
  INV_X1    g038(.A(new_n233), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n236), .B(new_n237), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n223), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n236), .B1(new_n239), .B2(new_n240), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n214), .A2(new_n242), .A3(new_n222), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n237), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n208), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT29), .B1(new_n232), .B2(new_n240), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n238), .A2(new_n233), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT3), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT83), .B1(new_n251), .B2(new_n223), .ZN(new_n252));
  INV_X1    g051(.A(new_n250), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(new_n233), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n242), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT83), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n214), .A2(new_n222), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n208), .B1(new_n244), .B2(new_n246), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n252), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n248), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n262), .B1(new_n248), .B2(new_n260), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n207), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n260), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n261), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n248), .A2(new_n260), .A3(new_n262), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(new_n206), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT64), .Z(new_n272));
  INV_X1    g071(.A(G127gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(G134gat), .ZN(new_n274));
  INV_X1    g073(.A(G134gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(G127gat), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT70), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G113gat), .ZN(new_n278));
  INV_X1    g077(.A(G120gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(G113gat), .B2(G120gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(G127gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n273), .A2(G134gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n277), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n289), .B(new_n286), .C1(new_n280), .C2(new_n282), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n294), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(KEYINPUT23), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n307));
  INV_X1    g106(.A(G169gat), .ZN(new_n308));
  INV_X1    g107(.A(G176gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n305), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n299), .A2(new_n304), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n299), .A2(KEYINPUT68), .A3(new_n304), .A4(new_n311), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n294), .A2(new_n296), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT65), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n294), .A2(new_n318), .A3(new_n296), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n300), .B1(KEYINPUT23), .B2(new_n306), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n300), .A2(KEYINPUT23), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n314), .A2(new_n315), .B1(new_n323), .B2(new_n305), .ZN(new_n324));
  INV_X1    g123(.A(G183gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT27), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT27), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G183gat), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT28), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT27), .B(G183gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT28), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n329), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(new_n334), .A3(new_n293), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT26), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n302), .A2(new_n336), .A3(new_n303), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT69), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n300), .B1(new_n336), .B2(new_n306), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n337), .B2(new_n338), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n335), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n291), .B1(new_n324), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n314), .A2(new_n315), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n305), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n291), .ZN(new_n347));
  INV_X1    g146(.A(new_n342), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n272), .B1(new_n343), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(KEYINPUT73), .A2(KEYINPUT34), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n353));
  NOR2_X1   g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT32), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n343), .A2(new_n349), .A3(new_n272), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT71), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n343), .A2(new_n349), .A3(new_n359), .A4(new_n272), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n356), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G71gat), .B(G99gat), .Z(new_n362));
  XNOR2_X1  g161(.A(G15gat), .B(G43gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(KEYINPUT72), .A3(KEYINPUT33), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT72), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n358), .A2(new_n360), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(KEYINPUT32), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n358), .A2(new_n360), .A3(new_n364), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n364), .A2(KEYINPUT33), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI221_X4 g170(.A(new_n355), .B1(new_n361), .B2(new_n365), .C1(new_n368), .C2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n355), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n371), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n361), .A2(new_n365), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n202), .B(new_n270), .C1(new_n372), .C2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(KEYINPUT78), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  AND2_X1   g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT77), .B1(new_n346), .B2(new_n348), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n324), .A2(new_n384), .A3(new_n342), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n382), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n382), .A2(KEYINPUT29), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n324), .B2(new_n342), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n244), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n384), .B1(new_n324), .B2(new_n342), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n346), .A2(KEYINPUT77), .A3(new_n348), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n391), .A3(new_n387), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n346), .A2(new_n382), .A3(new_n348), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n392), .A2(new_n244), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n381), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n244), .A3(new_n393), .ZN(new_n396));
  INV_X1    g195(.A(new_n381), .ZN(new_n397));
  INV_X1    g196(.A(new_n388), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n390), .A2(new_n391), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(new_n382), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n396), .B(new_n397), .C1(new_n400), .C2(new_n244), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(KEYINPUT30), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n389), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT30), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n397), .A4(new_n396), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G1gat), .B(G29gat), .Z(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G57gat), .B(G85gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n288), .A2(KEYINPUT79), .A3(new_n290), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT79), .B1(new_n288), .B2(new_n290), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n245), .B(new_n412), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n223), .A2(new_n291), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n223), .A2(new_n291), .A3(KEYINPUT4), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n415), .A2(new_n416), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n257), .B1(new_n413), .B2(new_n414), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n416), .B1(new_n422), .B2(new_n417), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n223), .A2(new_n291), .A3(KEYINPUT4), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT4), .B1(new_n223), .B2(new_n291), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n428), .A2(KEYINPUT5), .A3(new_n416), .A4(new_n415), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n411), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n425), .A2(new_n411), .A3(new_n429), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n425), .A2(KEYINPUT6), .A3(new_n411), .A4(new_n429), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT86), .B1(new_n406), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n438));
  AOI221_X4 g237(.A(new_n438), .B1(new_n434), .B2(new_n435), .C1(new_n402), .C2(new_n405), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n377), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n265), .A2(new_n269), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n374), .A2(new_n375), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n355), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n374), .A2(new_n373), .A3(new_n375), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n433), .A2(new_n432), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT81), .B1(new_n446), .B2(new_n430), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n431), .A2(new_n448), .A3(new_n432), .A4(new_n433), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n449), .A3(new_n435), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n406), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n202), .B1(new_n445), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n441), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n443), .A2(KEYINPUT36), .A3(new_n444), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT36), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n372), .B2(new_n376), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n433), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n416), .B1(new_n428), .B2(new_n415), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT39), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n411), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n416), .ZN(new_n463));
  INV_X1    g262(.A(new_n415), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n419), .A2(new_n420), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n422), .A2(new_n416), .A3(new_n417), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(KEYINPUT39), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n459), .B1(new_n469), .B2(KEYINPUT40), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n462), .A2(new_n468), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT40), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT84), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n474));
  AOI211_X1 g273(.A(new_n474), .B(KEYINPUT40), .C1(new_n462), .C2(new_n468), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n470), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n270), .B1(new_n406), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT37), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n396), .B(new_n479), .C1(new_n400), .C2(new_n244), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n381), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT38), .ZN(new_n482));
  INV_X1    g281(.A(new_n244), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n392), .A2(new_n483), .A3(new_n393), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT37), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n483), .B1(new_n386), .B2(new_n388), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n401), .B(new_n435), .C1(new_n446), .C2(new_n430), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n478), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n435), .ZN(new_n491));
  INV_X1    g290(.A(new_n446), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(new_n431), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n484), .B(KEYINPUT37), .C1(new_n400), .C2(new_n483), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n480), .A2(new_n494), .A3(new_n482), .A4(new_n381), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n493), .A2(new_n495), .A3(KEYINPUT85), .A4(new_n401), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n479), .B1(new_n403), .B2(new_n396), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT38), .B1(new_n498), .B2(new_n481), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n477), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI22_X1  g299(.A1(new_n440), .A2(new_n453), .B1(new_n458), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(KEYINPUT90), .B(KEYINPUT17), .Z(new_n503));
  INV_X1    g302(.A(G43gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n204), .ZN(new_n505));
  NAND2_X1  g304(.A1(G43gat), .A2(G50gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(KEYINPUT87), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G29gat), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT14), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(G29gat), .B2(G36gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT88), .ZN(new_n517));
  NAND2_X1  g316(.A1(G29gat), .A2(G36gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT88), .B1(new_n514), .B2(new_n516), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n507), .B(new_n511), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n506), .ZN(new_n522));
  NOR2_X1   g321(.A1(G43gat), .A2(G50gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n510), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n507), .A3(KEYINPUT15), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n508), .A3(new_n506), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n514), .A2(new_n516), .A3(new_n518), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n521), .A2(KEYINPUT89), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT89), .B1(new_n521), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n503), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT16), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(G1gat), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(G1gat), .B2(new_n532), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(G8gat), .Z(new_n536));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT17), .A3(new_n528), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n531), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT91), .Z(new_n540));
  INV_X1    g339(.A(new_n536), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n521), .A2(new_n528), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n521), .A2(KEYINPUT89), .A3(new_n528), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n538), .A2(new_n540), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT18), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n538), .A2(KEYINPUT18), .A3(new_n540), .A4(new_n547), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n544), .A3(new_n545), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n540), .B(KEYINPUT13), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n550), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G197gat), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT11), .B(G169gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT12), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n548), .A2(new_n549), .B1(new_n553), .B2(new_n555), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(new_n562), .A3(new_n551), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OR2_X1    g366(.A1(G71gat), .A2(G78gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(G71gat), .A2(G78gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G64gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G57gat), .ZN(new_n572));
  INV_X1    g371(.A(G57gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(G64gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n570), .B1(KEYINPUT9), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT92), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(new_n571), .B2(G57gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(KEYINPUT92), .A3(G64gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(new_n572), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n569), .B1(new_n568), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT93), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n580), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n576), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT21), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  AND2_X1   g390(.A1(new_n591), .A2(new_n273), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n273), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n536), .B(new_n588), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n536), .A2(new_n588), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n273), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT94), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G155gat), .ZN(new_n601));
  XOR2_X1   g400(.A(G183gat), .B(G211gat), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n594), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n603), .B1(new_n594), .B2(new_n598), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G85gat), .A2(G92gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT7), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT7), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(G85gat), .A3(G92gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G99gat), .B(G106gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  INV_X1    g412(.A(G85gat), .ZN(new_n614));
  INV_X1    g413(.A(G92gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(KEYINPUT8), .A2(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n612), .B1(new_n611), .B2(new_n616), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n546), .A2(new_n619), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n619), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n531), .A2(new_n537), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(KEYINPUT96), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT95), .Z(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(KEYINPUT96), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT97), .ZN(new_n635));
  INV_X1    g434(.A(new_n632), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n624), .A2(new_n627), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n635), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n636), .B1(new_n624), .B2(new_n627), .ZN(new_n640));
  AOI211_X1 g439(.A(new_n626), .B(new_n632), .C1(new_n621), .C2(new_n623), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n606), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n584), .A2(new_n586), .ZN(new_n646));
  INV_X1    g445(.A(new_n576), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n646), .A2(KEYINPUT10), .A3(new_n619), .A4(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n587), .A2(KEYINPUT99), .A3(KEYINPUT10), .A4(new_n619), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n646), .A2(new_n647), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n622), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n587), .A2(new_n619), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT98), .B(KEYINPUT10), .Z(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G230gat), .A2(G233gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(G176gat), .B(G204gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n661), .B(new_n662), .Z(new_n663));
  AND2_X1   g462(.A1(new_n654), .A2(new_n655), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n660), .B(new_n663), .C1(new_n659), .C2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n663), .ZN(new_n666));
  INV_X1    g465(.A(new_n659), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n652), .B2(new_n657), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n664), .A2(new_n659), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n645), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n502), .A2(new_n567), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n450), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT100), .B(G1gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1324gat));
  INV_X1    g477(.A(new_n406), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n683), .A2(KEYINPUT101), .A3(KEYINPUT42), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n680), .B2(G8gat), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(new_n683), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT101), .B1(new_n683), .B2(KEYINPUT42), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n684), .B1(new_n687), .B2(new_n688), .ZN(G1325gat));
  INV_X1    g488(.A(G15gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n372), .A2(new_n376), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n674), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n455), .A2(new_n457), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n674), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n696), .B2(new_n690), .ZN(G1326gat));
  NAND2_X1  g496(.A1(new_n674), .A2(new_n441), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NOR2_X1   g499(.A1(new_n502), .A2(new_n567), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n606), .A2(new_n672), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n643), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n701), .A2(new_n512), .A3(new_n675), .A4(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(KEYINPUT103), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n488), .A2(new_n478), .A3(new_n489), .ZN(new_n710));
  INV_X1    g509(.A(new_n489), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT85), .B1(new_n711), .B2(new_n495), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n499), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n477), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n406), .A2(new_n436), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n438), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n406), .A2(KEYINPUT86), .A3(new_n436), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n445), .A2(new_n718), .A3(new_n202), .A4(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n270), .B1(new_n372), .B2(new_n376), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT35), .B1(new_n721), .B2(new_n451), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  AOI211_X1 g522(.A(new_n643), .B(new_n708), .C1(new_n716), .C2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n501), .B2(new_n644), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n702), .A2(new_n567), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n727), .A2(new_n450), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n706), .B1(new_n512), .B2(new_n730), .ZN(G1328gat));
  NOR2_X1   g530(.A1(new_n727), .A2(new_n729), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n679), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(KEYINPUT104), .A3(new_n679), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(G36gat), .A3(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n701), .A2(new_n513), .A3(new_n679), .A4(new_n703), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT46), .Z(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1329gat));
  OAI211_X1 g539(.A(new_n695), .B(new_n728), .C1(new_n724), .C2(new_n726), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n504), .B1(new_n741), .B2(KEYINPUT107), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(KEYINPUT107), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n564), .A2(new_n566), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n691), .A2(G43gat), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n501), .A2(new_n744), .A3(new_n703), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT106), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n741), .A2(G43gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n747), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(G1330gat));
  AND4_X1   g553(.A1(new_n204), .A2(new_n701), .A3(new_n441), .A4(new_n703), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n441), .B(new_n728), .C1(new_n724), .C2(new_n726), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT109), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G50gat), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n758), .A2(KEYINPUT109), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n758), .A2(new_n763), .A3(G50gat), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n758), .B2(G50gat), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n764), .A2(new_n765), .A3(new_n755), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n762), .B1(new_n766), .B2(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g566(.A1(new_n501), .A2(new_n567), .A3(new_n645), .A4(new_n671), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n675), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT110), .B(G57gat), .Z(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1332gat));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n679), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT49), .B(G64gat), .Z(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n772), .B2(new_n774), .ZN(G1333gat));
  NAND2_X1  g574(.A1(new_n768), .A2(new_n695), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n691), .A2(G71gat), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n776), .A2(G71gat), .B1(new_n768), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g578(.A1(new_n768), .A2(new_n441), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g580(.A(new_n643), .B1(new_n716), .B2(new_n723), .ZN(new_n782));
  INV_X1    g581(.A(new_n606), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(new_n744), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n782), .A2(KEYINPUT51), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT51), .B1(new_n782), .B2(new_n784), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n787), .A2(new_n614), .A3(new_n675), .A4(new_n671), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n501), .B(new_n644), .C1(KEYINPUT103), .C2(new_n707), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n782), .B2(new_n725), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n783), .A2(new_n744), .A3(new_n672), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n792), .A2(new_n675), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n788), .B1(new_n793), .B2(new_n614), .ZN(G1336gat));
  NOR3_X1   g593(.A1(new_n406), .A2(G92gat), .A3(new_n672), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n790), .A2(new_n679), .A3(new_n791), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n799), .A2(G92gat), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n795), .B(KEYINPUT111), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n787), .A2(new_n801), .B1(new_n799), .B2(G92gat), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n798), .A2(new_n800), .B1(new_n802), .B2(new_n797), .ZN(G1337gat));
  NAND2_X1  g602(.A1(new_n792), .A2(new_n695), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G99gat), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n691), .A2(G99gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n787), .A2(new_n671), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1338gat));
  OAI211_X1 g607(.A(new_n441), .B(new_n791), .C1(new_n724), .C2(new_n726), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n809), .A2(G106gat), .B1(KEYINPUT112), .B2(KEYINPUT53), .ZN(new_n810));
  OR2_X1    g609(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n270), .A2(G106gat), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n671), .B(new_n812), .C1(new_n785), .C2(new_n786), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n811), .B1(new_n810), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(G1339gat));
  NAND3_X1  g615(.A1(new_n652), .A2(new_n667), .A3(new_n657), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT113), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n652), .A2(new_n657), .A3(new_n819), .A4(new_n667), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n818), .A2(new_n660), .A3(KEYINPUT54), .A4(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n663), .B1(new_n668), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n823), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n744), .A2(new_n665), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n540), .B1(new_n538), .B2(new_n547), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n829), .A2(KEYINPUT114), .B1(new_n553), .B2(new_n555), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n831), .B(new_n540), .C1(new_n538), .C2(new_n547), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n561), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n566), .A3(new_n671), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n644), .B1(new_n828), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n826), .A2(new_n665), .A3(new_n827), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n833), .A2(new_n638), .A3(new_n642), .A4(new_n566), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n606), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n645), .A2(new_n567), .A3(new_n672), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n721), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n675), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n406), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(new_n278), .A3(new_n567), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n842), .B(KEYINPUT115), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n406), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n744), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(new_n278), .ZN(G1340gat));
  NOR3_X1   g647(.A1(new_n843), .A2(new_n279), .A3(new_n672), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n671), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n279), .ZN(G1341gat));
  NAND3_X1  g650(.A1(new_n846), .A2(new_n273), .A3(new_n783), .ZN(new_n852));
  OAI21_X1  g651(.A(G127gat), .B1(new_n843), .B2(new_n606), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1342gat));
  NOR2_X1   g653(.A1(new_n679), .A2(new_n643), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n845), .A2(new_n275), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n275), .B1(new_n842), .B2(new_n855), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT116), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n860), .A3(new_n275), .A4(new_n855), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n857), .A2(new_n859), .A3(new_n861), .ZN(G1343gat));
  AOI21_X1  g661(.A(new_n270), .B1(new_n839), .B2(new_n840), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n679), .A2(new_n450), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n694), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n215), .A3(new_n744), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n836), .A2(KEYINPUT117), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n826), .A2(new_n871), .A3(new_n665), .A4(new_n827), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n744), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n644), .B1(new_n873), .B2(new_n834), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n606), .B1(new_n874), .B2(new_n838), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n840), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n869), .B1(new_n876), .B2(new_n441), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n863), .A2(new_n869), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n866), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n877), .A2(new_n879), .A3(new_n567), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n868), .B1(new_n880), .B2(new_n215), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT58), .ZN(G1344gat));
  NAND4_X1  g681(.A1(new_n863), .A2(new_n866), .A3(new_n217), .A4(new_n671), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT118), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n865), .A2(KEYINPUT119), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n865), .A2(KEYINPUT119), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n671), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n834), .B1(new_n836), .B2(new_n567), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n838), .B1(new_n888), .B2(new_n643), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n840), .B1(new_n889), .B2(new_n783), .ZN(new_n890));
  AND4_X1   g689(.A1(KEYINPUT120), .A2(new_n890), .A3(KEYINPUT57), .A4(new_n441), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT120), .B1(new_n863), .B2(KEYINPUT57), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n840), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n567), .B1(new_n836), .B2(KEYINPUT117), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n833), .A2(new_n566), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n895), .A2(new_n872), .B1(new_n671), .B2(new_n896), .ZN(new_n897));
  OAI22_X1  g696(.A1(new_n897), .A2(new_n644), .B1(new_n836), .B2(new_n837), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n894), .B1(new_n898), .B2(new_n606), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n869), .B1(new_n899), .B2(new_n270), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n887), .B1(new_n893), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n884), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n865), .B1(new_n863), .B2(new_n869), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n899), .A2(new_n270), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n904), .B(new_n671), .C1(new_n905), .C2(new_n869), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT59), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT121), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n890), .A2(KEYINPUT57), .A3(new_n441), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n863), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT57), .B1(new_n876), .B2(new_n441), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT59), .B(G148gat), .C1(new_n915), .C2(new_n887), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n877), .A2(new_n879), .A3(new_n672), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n217), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n916), .A2(new_n919), .A3(new_n920), .A4(new_n884), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n908), .A2(new_n921), .ZN(G1345gat));
  OAI21_X1  g721(.A(new_n904), .B1(new_n905), .B2(new_n869), .ZN(new_n923));
  OAI21_X1  g722(.A(G155gat), .B1(new_n923), .B2(new_n606), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n867), .A2(new_n210), .A3(new_n783), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1346gat));
  OAI21_X1  g725(.A(G162gat), .B1(new_n923), .B2(new_n643), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n867), .A2(new_n211), .A3(new_n644), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1347gat));
  NOR2_X1   g728(.A1(new_n675), .A2(new_n406), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n841), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n308), .A3(new_n744), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n692), .A2(new_n930), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(KEYINPUT122), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(KEYINPUT122), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n934), .A2(new_n935), .A3(new_n441), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n890), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n744), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT123), .B1(new_n939), .B2(G169gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n932), .B1(new_n940), .B2(new_n941), .ZN(G1348gat));
  AOI21_X1  g741(.A(G176gat), .B1(new_n931), .B2(new_n671), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT124), .Z(new_n944));
  NOR3_X1   g743(.A1(new_n937), .A2(new_n309), .A3(new_n672), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n944), .A2(new_n945), .ZN(G1349gat));
  OAI21_X1  g745(.A(G183gat), .B1(new_n937), .B2(new_n606), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n332), .A3(new_n783), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g749(.A1(new_n931), .A2(new_n329), .A3(new_n644), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n938), .A2(new_n644), .ZN(new_n952));
  XNOR2_X1  g751(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n952), .A2(G190gat), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n952), .B2(G190gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(G1351gat));
  AND2_X1   g755(.A1(new_n694), .A2(new_n930), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n957), .B1(new_n913), .B2(new_n914), .ZN(new_n958));
  INV_X1    g757(.A(G197gat), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n958), .A2(new_n959), .A3(new_n567), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n694), .A2(new_n441), .A3(new_n930), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n890), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n744), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n960), .A2(new_n964), .ZN(G1352gat));
  OAI21_X1  g764(.A(G204gat), .B1(new_n958), .B2(new_n672), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n963), .A2(new_n227), .A3(new_n671), .ZN(new_n967));
  AND2_X1   g766(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n968));
  NOR2_X1   g767(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n966), .B(new_n970), .C1(new_n968), .C2(new_n967), .ZN(G1353gat));
  OR3_X1    g770(.A1(new_n962), .A2(G211gat), .A3(new_n606), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n783), .B(new_n957), .C1(new_n913), .C2(new_n914), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  OAI211_X1 g775(.A(new_n644), .B(new_n957), .C1(new_n913), .C2(new_n914), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(G218gat), .ZN(new_n978));
  OR3_X1    g777(.A1(new_n962), .A2(G218gat), .A3(new_n643), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n978), .A2(KEYINPUT127), .A3(new_n979), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1355gat));
endmodule


