//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT30), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G128), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT64), .A2(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT64), .A2(G143), .ZN(new_n192));
  AOI21_X1  g006(.A(G146), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT65), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT65), .A2(G146), .ZN(new_n195));
  AOI21_X1  g009(.A(G143), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n190), .B1(new_n193), .B2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(G143), .A3(new_n195), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n191), .A2(G146), .A3(new_n192), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT69), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI211_X1 g019(.A(KEYINPUT66), .B(new_n204), .C1(new_n205), .C2(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(KEYINPUT68), .A3(G137), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT68), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G134), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT11), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G134), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(KEYINPUT11), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n203), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n210), .A2(new_n207), .ZN(new_n218));
  OAI22_X1  g032(.A1(KEYINPUT66), .A2(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n204), .A2(KEYINPUT66), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n218), .A2(new_n221), .A3(KEYINPUT69), .A4(new_n206), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n217), .A2(new_n222), .A3(G131), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT67), .B(G131), .Z(new_n224));
  NAND4_X1  g038(.A1(new_n218), .A2(new_n221), .A3(new_n224), .A4(new_n206), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n202), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT70), .B1(new_n209), .B2(G134), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n214), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n209), .A2(KEYINPUT70), .A3(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(G131), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n198), .A2(new_n199), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n198), .A2(new_n199), .A3(KEYINPUT71), .A4(new_n233), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G128), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT64), .A2(G143), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT64), .A2(G143), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT65), .A2(G146), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT65), .A2(G146), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n240), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n231), .B1(new_n238), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n188), .B1(new_n226), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT72), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT76), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT2), .A2(G113), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AND3_X1   g070(.A1(KEYINPUT73), .A2(KEYINPUT2), .A3(G113), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT73), .B1(KEYINPUT2), .B2(G113), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(G116), .B(G119), .Z(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n260), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT74), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT2), .A2(G113), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(KEYINPUT73), .A2(KEYINPUT2), .A3(G113), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT74), .A3(new_n256), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n263), .B1(new_n265), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n262), .B1(new_n272), .B2(KEYINPUT75), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n274));
  AOI211_X1 g088(.A(new_n274), .B(new_n263), .C1(new_n265), .C2(new_n271), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n254), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT74), .B1(new_n270), .B2(new_n256), .ZN(new_n277));
  AOI211_X1 g091(.A(new_n264), .B(new_n255), .C1(new_n268), .C2(new_n269), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n260), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n274), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n272), .A2(KEYINPUT75), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT76), .A4(new_n262), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n284), .B(new_n188), .C1(new_n226), .C2(new_n251), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n238), .A2(new_n250), .ZN(new_n286));
  INV_X1    g100(.A(new_n231), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT77), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n189), .B1(new_n244), .B2(new_n248), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n197), .A2(KEYINPUT77), .A3(new_n201), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n225), .ZN(new_n295));
  INV_X1    g109(.A(G131), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n218), .A2(new_n221), .A3(new_n206), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n296), .B1(new_n297), .B2(new_n203), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n298), .B2(new_n222), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n288), .B(KEYINPUT30), .C1(new_n294), .C2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n253), .A2(new_n283), .A3(new_n285), .A4(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n290), .A2(new_n291), .A3(new_n289), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT77), .B1(new_n197), .B2(new_n201), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n223), .A2(new_n225), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n306), .A2(new_n307), .B1(new_n286), .B2(new_n287), .ZN(new_n308));
  AOI22_X1  g122(.A1(KEYINPUT72), .A2(new_n252), .B1(new_n308), .B2(KEYINPUT30), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n309), .A2(KEYINPUT78), .A3(new_n283), .A4(new_n285), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n276), .A2(new_n312), .A3(new_n282), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(new_n276), .B2(new_n282), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n236), .A2(new_n237), .B1(new_n240), .B2(new_n249), .ZN(new_n315));
  OAI22_X1  g129(.A1(new_n299), .A2(new_n294), .B1(new_n315), .B2(new_n231), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT80), .B(KEYINPUT27), .ZN(new_n318));
  INV_X1    g132(.A(G237), .ZN(new_n319));
  INV_X1    g133(.A(G953), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(G210), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n318), .B(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G101), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n311), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT31), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT31), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n311), .A2(new_n328), .A3(new_n325), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n324), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n273), .A2(new_n254), .A3(new_n275), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n261), .B1(new_n279), .B2(new_n274), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT76), .B1(new_n333), .B2(new_n281), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT79), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n316), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n276), .A2(new_n312), .A3(new_n282), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n288), .B(KEYINPUT81), .C1(new_n294), .C2(new_n299), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n335), .A2(new_n337), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n340), .A2(KEYINPUT82), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT82), .B1(new_n340), .B2(new_n341), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n226), .A2(new_n251), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(new_n276), .B2(new_n282), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT28), .B1(new_n317), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n331), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n187), .B1(new_n330), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT32), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI211_X1 g165(.A(new_n317), .B(new_n331), .C1(new_n303), .C2(new_n310), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n353));
  AOI21_X1  g167(.A(G902), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n308), .B1(new_n335), .B2(new_n338), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT28), .B1(new_n317), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n353), .B1(new_n344), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n340), .A2(new_n341), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n340), .A2(KEYINPUT82), .A3(new_n341), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n360), .A2(new_n353), .A3(new_n347), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n331), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n354), .B1(new_n357), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G472), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n360), .A2(new_n361), .A3(new_n347), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n324), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n327), .A3(new_n329), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n351), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G214), .B1(G237), .B2(G902), .ZN(new_n371));
  NAND2_X1  g185(.A1(G234), .A2(G237), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(G952), .A3(new_n320), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(G902), .A3(G953), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT21), .B(G898), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT6), .ZN(new_n380));
  INV_X1    g194(.A(G101), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n382), .A2(KEYINPUT3), .A3(G107), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  AND2_X1   g198(.A1(KEYINPUT88), .A2(G104), .ZN(new_n385));
  NOR2_X1   g199(.A1(KEYINPUT88), .A2(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n383), .B1(new_n387), .B2(KEYINPUT3), .ZN(new_n388));
  OR2_X1    g202(.A1(KEYINPUT88), .A2(G104), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT88), .A2(G104), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(G107), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n381), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n392), .A2(KEYINPUT4), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT89), .ZN(new_n394));
  INV_X1    g208(.A(new_n383), .ZN(new_n395));
  AOI21_X1  g209(.A(G107), .B1(new_n389), .B2(new_n390), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n391), .A2(new_n381), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n394), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n391), .A2(new_n381), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n388), .A3(KEYINPUT89), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n392), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n393), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n283), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n382), .A2(G107), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n381), .B1(new_n387), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n398), .A2(new_n394), .A3(new_n399), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT89), .B1(new_n401), .B2(new_n388), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G113), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT92), .B(KEYINPUT5), .Z(new_n414));
  INV_X1    g228(.A(G116), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G119), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n413), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n260), .B2(new_n414), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n262), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n412), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n406), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G110), .B(G122), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n380), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n420), .B1(new_n283), .B2(new_n405), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n426), .A2(KEYINPUT93), .A3(new_n423), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT93), .B1(new_n426), .B2(new_n423), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n422), .A2(new_n380), .A3(new_n424), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n202), .A2(G125), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n431), .A2(KEYINPUT94), .ZN(new_n432));
  INV_X1    g246(.A(G125), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n315), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(KEYINPUT94), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT95), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n436), .A2(KEYINPUT95), .ZN(new_n439));
  INV_X1    g253(.A(G224), .ZN(new_n440));
  OAI22_X1  g254(.A1(new_n438), .A2(new_n439), .B1(new_n440), .B2(G953), .ZN(new_n441));
  INV_X1    g255(.A(new_n439), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n440), .A2(G953), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n443), .A3(new_n437), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n429), .A2(new_n430), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G210), .B1(G237), .B2(G902), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n406), .A2(new_n421), .A3(new_n423), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT93), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n426), .A2(KEYINPUT93), .A3(new_n423), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT7), .B1(new_n440), .B2(G953), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n436), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n408), .B1(new_n400), .B2(new_n402), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n456), .A2(new_n417), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n455), .B1(new_n261), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n423), .B(KEYINPUT8), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n458), .B(new_n459), .C1(new_n455), .C2(new_n419), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n436), .A2(new_n453), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n454), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n452), .B2(new_n462), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n446), .A2(new_n447), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n447), .B1(new_n446), .B2(new_n463), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n371), .B(new_n379), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G110), .B(G140), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n320), .A2(G227), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n412), .A2(new_n315), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n198), .A2(new_n199), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n232), .B1(new_n244), .B2(KEYINPUT1), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n238), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n455), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n307), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT12), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(KEYINPUT12), .A3(new_n307), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT10), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n315), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n476), .A2(new_n483), .B1(new_n484), .B2(new_n455), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n405), .A2(new_n306), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n307), .B(KEYINPUT90), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n470), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT12), .B1(new_n477), .B2(new_n307), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n479), .B(new_n299), .C1(new_n471), .C2(new_n476), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n488), .B(new_n470), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n469), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n469), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n299), .B1(new_n485), .B2(new_n486), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(G469), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G469), .ZN(new_n501));
  INV_X1    g315(.A(G902), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n469), .B1(new_n504), .B2(new_n497), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n488), .B(new_n495), .C1(new_n490), .C2(new_n491), .ZN(new_n506));
  AOI21_X1  g320(.A(G902), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n503), .B1(new_n507), .B2(new_n501), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n500), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G478), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT9), .B(G234), .ZN(new_n513));
  INV_X1    g327(.A(G217), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n513), .A2(new_n514), .A3(G953), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n245), .A2(G128), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT101), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n242), .A2(new_n243), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n518), .B1(new_n519), .B2(G128), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n518), .A3(G128), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT13), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n517), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n522), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(new_n520), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT13), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n205), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n517), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n205), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G116), .B(G122), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n532), .A2(new_n384), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n384), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n531), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT14), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n415), .A2(KEYINPUT14), .A3(G122), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G107), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n534), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G134), .B1(new_n527), .B2(new_n517), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n531), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n516), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n544), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n546), .B(new_n515), .C1(new_n529), .C2(new_n536), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n512), .B1(new_n548), .B2(new_n502), .ZN(new_n549));
  AOI211_X1 g363(.A(G902), .B(new_n511), .C1(new_n545), .C2(new_n547), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT100), .ZN(new_n552));
  INV_X1    g366(.A(G140), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G125), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n433), .A2(G140), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT84), .ZN(new_n556));
  OR3_X1    g370(.A1(new_n433), .A2(KEYINPUT84), .A3(G140), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT16), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n554), .A2(KEYINPUT16), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(G146), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT16), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n556), .B2(new_n557), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n564), .A2(new_n241), .A3(new_n560), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT99), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n319), .A2(new_n320), .A3(G214), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n191), .A3(new_n192), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT96), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT96), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n519), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  INV_X1    g385(.A(new_n567), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G143), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n224), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n568), .A2(KEYINPUT96), .B1(new_n572), .B2(G143), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n224), .A3(new_n571), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n574), .A2(KEYINPUT17), .A3(new_n575), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n559), .A2(G146), .A3(new_n561), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n241), .B1(new_n564), .B2(new_n560), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n566), .A2(new_n580), .A3(new_n581), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(KEYINPUT18), .A2(G131), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n574), .B(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n246), .A2(new_n247), .ZN(new_n589));
  XNOR2_X1  g403(.A(G125), .B(G140), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n558), .B2(new_n241), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(G113), .B(G122), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT98), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(new_n382), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n552), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n586), .A2(new_n593), .A3(KEYINPUT100), .A4(new_n597), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n599), .A2(new_n600), .B1(new_n594), .B2(new_n598), .ZN(new_n601));
  OAI21_X1  g415(.A(G475), .B1(new_n601), .B2(G902), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT20), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n599), .A2(new_n600), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n558), .A2(KEYINPUT19), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n590), .A2(KEYINPUT19), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n589), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n582), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT97), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n576), .A2(new_n579), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n608), .A2(new_n612), .A3(new_n582), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n597), .B1(new_n614), .B2(new_n593), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n604), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(G475), .A2(G902), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n603), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n615), .B1(new_n599), .B2(new_n600), .ZN(new_n620));
  INV_X1    g434(.A(new_n618), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n620), .A2(KEYINPUT20), .A3(new_n621), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n551), .B(new_n602), .C1(new_n619), .C2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(G221), .B1(new_n513), .B2(G902), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n509), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n466), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(G110), .ZN(new_n628));
  INV_X1    g442(.A(G119), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(G128), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n232), .A2(KEYINPUT23), .A3(G119), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n629), .A2(G128), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(KEYINPUT23), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n628), .B1(new_n633), .B2(KEYINPUT83), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(KEYINPUT83), .B2(new_n633), .ZN(new_n635));
  INV_X1    g449(.A(new_n632), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n630), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT24), .B(G110), .ZN(new_n638));
  OAI221_X1 g452(.A(new_n635), .B1(new_n637), .B2(new_n638), .C1(new_n562), .C2(new_n565), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n320), .A2(G221), .A3(G234), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT22), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G137), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n637), .A2(new_n638), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n643), .B1(new_n633), .B2(G110), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n582), .A2(new_n591), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n639), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT86), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT86), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n639), .A2(new_n648), .A3(new_n642), .A4(new_n645), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n639), .A2(new_n645), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT85), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n642), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n647), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n514), .B1(G234), .B2(new_n502), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(G902), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT87), .B1(new_n654), .B2(G902), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n659), .A2(KEYINPUT25), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(KEYINPUT25), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n656), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n370), .A2(new_n627), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G101), .ZN(G3));
  OR2_X1    g481(.A1(new_n619), .A2(new_n622), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n602), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT33), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n548), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n545), .A2(KEYINPUT33), .A3(new_n547), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n671), .A2(G478), .A3(new_n502), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n548), .A2(new_n502), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n510), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n673), .A2(new_n678), .A3(new_n675), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n669), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n466), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n368), .A2(new_n502), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n683), .A2(G472), .B1(new_n187), .B2(new_n368), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(KEYINPUT91), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n495), .B1(new_n686), .B2(new_n492), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n501), .A3(new_n498), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n505), .A2(new_n506), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n501), .A3(new_n502), .ZN(new_n690));
  INV_X1    g504(.A(new_n503), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n625), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n693), .A2(new_n664), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n682), .A2(new_n684), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT34), .B(G104), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G6));
  INV_X1    g512(.A(new_n551), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n668), .A2(new_n699), .A3(new_n602), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n466), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n684), .A3(new_n695), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT35), .B(G107), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G9));
  NOR2_X1   g518(.A1(new_n652), .A2(KEYINPUT36), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n650), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n657), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n662), .B2(new_n663), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n627), .A2(new_n684), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT103), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT37), .B(G110), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G12));
  NOR2_X1   g526(.A1(new_n464), .A2(new_n465), .ZN(new_n713));
  INV_X1    g527(.A(new_n371), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n370), .A2(new_n715), .A3(new_n708), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n373), .B(KEYINPUT104), .Z(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(G900), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n718), .B1(new_n719), .B2(new_n376), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n700), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n693), .A2(new_n694), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G128), .ZN(G30));
  XOR2_X1   g539(.A(new_n720), .B(KEYINPUT39), .Z(new_n726));
  NAND2_X1  g540(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT40), .ZN(new_n728));
  INV_X1    g542(.A(new_n669), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n728), .A2(new_n714), .A3(new_n551), .A4(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n708), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n368), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT32), .B1(new_n368), .B2(new_n187), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n311), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n331), .B1(new_n735), .B2(new_n317), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n317), .A2(new_n355), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n502), .B1(new_n739), .B2(new_n331), .ZN(new_n740));
  OAI21_X1  g554(.A(G472), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n446), .A2(new_n463), .ZN(new_n743));
  INV_X1    g557(.A(new_n447), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n446), .A2(new_n447), .A3(new_n463), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT38), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n730), .A2(new_n731), .A3(new_n742), .A4(new_n748), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(new_n519), .Z(G45));
  INV_X1    g564(.A(new_n720), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n669), .A2(new_n680), .A3(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n752), .A2(new_n694), .A3(new_n693), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n716), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G146), .ZN(G48));
  NOR2_X1   g569(.A1(new_n507), .A2(new_n501), .ZN(new_n756));
  AOI211_X1 g570(.A(G469), .B(G902), .C1(new_n505), .C2(new_n506), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n625), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n664), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n370), .A2(new_n682), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT105), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n370), .A2(new_n682), .A3(new_n760), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT41), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G113), .ZN(G15));
  NAND3_X1  g581(.A1(new_n370), .A2(new_n701), .A3(new_n760), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT106), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n370), .A2(new_n701), .A3(new_n760), .A4(KEYINPUT106), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G116), .ZN(G18));
  NAND2_X1  g587(.A1(new_n708), .A2(new_n624), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n774), .B1(new_n734), .B2(new_n365), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n747), .A2(new_n371), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(new_n759), .A3(new_n378), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G119), .ZN(G21));
  AOI21_X1  g593(.A(new_n331), .B1(new_n344), .B2(new_n356), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n187), .B1(new_n330), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n327), .A2(new_n329), .ZN(new_n782));
  AOI21_X1  g596(.A(G902), .B1(new_n782), .B2(new_n367), .ZN(new_n783));
  INV_X1    g597(.A(G472), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n665), .B(new_n781), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n551), .B1(new_n668), .B2(new_n602), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n756), .A2(new_n757), .A3(new_n378), .A4(new_n694), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n747), .A2(new_n786), .A3(new_n787), .A4(new_n371), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(G122), .Z(G24));
  NOR2_X1   g604(.A1(new_n783), .A2(new_n784), .ZN(new_n791));
  INV_X1    g605(.A(new_n781), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n791), .A2(new_n731), .A3(new_n752), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n776), .A2(new_n759), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G125), .ZN(G27));
  AOI21_X1  g610(.A(new_n664), .B1(new_n734), .B2(new_n365), .ZN(new_n797));
  INV_X1    g611(.A(new_n752), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT107), .B1(new_n688), .B2(new_n692), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT107), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n500), .A2(new_n800), .A3(new_n508), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n694), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n747), .A2(new_n714), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT108), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n804), .B1(new_n802), .B2(new_n803), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n797), .B(new_n798), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT42), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n799), .A2(new_n801), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n625), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n713), .A2(new_n371), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT108), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT42), .A3(new_n797), .A4(new_n798), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G131), .ZN(G33));
  OAI211_X1 g632(.A(new_n797), .B(new_n721), .C1(new_n805), .C2(new_n806), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G134), .ZN(G36));
  NAND3_X1  g634(.A1(new_n729), .A2(KEYINPUT43), .A3(new_n680), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT110), .Z(new_n822));
  INV_X1    g636(.A(KEYINPUT109), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n669), .B1(new_n823), .B2(new_n680), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n823), .B2(new_n680), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT43), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n731), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n684), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(KEYINPUT44), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT44), .B1(new_n828), .B2(new_n829), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n803), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n822), .A2(new_n827), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n829), .A3(new_n708), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT44), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(KEYINPUT111), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT112), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n830), .A2(new_n803), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(KEYINPUT111), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n831), .A2(new_n832), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n499), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT45), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n687), .B2(new_n498), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n847), .A3(G469), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT46), .B1(new_n848), .B2(new_n691), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n757), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(KEYINPUT46), .A3(new_n691), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n694), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n726), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n839), .A2(new_n844), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT113), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(new_n209), .ZN(G39));
  XNOR2_X1  g671(.A(new_n852), .B(KEYINPUT47), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n370), .A2(new_n812), .A3(new_n665), .A4(new_n752), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(G140), .ZN(G42));
  XOR2_X1   g675(.A(new_n758), .B(KEYINPUT49), .Z(new_n862));
  NOR2_X1   g676(.A1(new_n694), .A2(new_n714), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n729), .A2(new_n665), .A3(new_n680), .A4(new_n863), .ZN(new_n864));
  OR4_X1    g678(.A1(new_n742), .A2(new_n748), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n834), .A2(new_n718), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT116), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n834), .A2(new_n868), .A3(new_n718), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n812), .A2(new_n759), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n797), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n871), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n867), .B2(new_n869), .ZN(new_n876));
  XOR2_X1   g690(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n797), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n871), .A2(new_n665), .A3(new_n374), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(new_n742), .ZN(new_n880));
  OAI211_X1 g694(.A(G952), .B(new_n320), .C1(new_n880), .C2(new_n681), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n785), .B1(new_n867), .B2(new_n869), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(new_n882), .B2(new_n794), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n874), .A2(new_n878), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT119), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n748), .A2(new_n371), .A3(new_n759), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT50), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n882), .A2(KEYINPUT50), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n880), .A2(new_n669), .A3(new_n680), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n791), .A2(new_n731), .A3(new_n792), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n876), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n882), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n756), .A2(new_n757), .A3(new_n625), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n858), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n897), .A2(new_n812), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n886), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n882), .B(new_n803), .C1(new_n902), .C2(new_n899), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n858), .A2(KEYINPUT117), .A3(new_n898), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n905), .A2(KEYINPUT51), .A3(new_n892), .A4(new_n895), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n885), .A2(new_n901), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n466), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n681), .A2(new_n700), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n684), .A2(new_n908), .A3(new_n909), .A4(new_n695), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n666), .A2(new_n709), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n793), .B1(new_n805), .B2(new_n806), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n775), .A2(new_n722), .A3(new_n751), .A4(new_n803), .ZN(new_n913));
  AND4_X1   g727(.A1(new_n819), .A2(new_n911), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n789), .B1(new_n775), .B2(new_n777), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n765), .A2(new_n772), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n916), .A3(new_n817), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT114), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n715), .A2(new_n786), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n920), .A2(new_n720), .A3(new_n811), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n731), .A3(new_n742), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n716), .B1(new_n723), .B2(new_n753), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n923), .A3(new_n795), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT52), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT52), .A4(new_n795), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n914), .A2(new_n916), .A3(KEYINPUT114), .A4(new_n817), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n919), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT53), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT54), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n911), .A2(new_n819), .A3(new_n912), .A4(new_n913), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n809), .B2(new_n816), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT114), .B1(new_n937), .B2(new_n916), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n929), .A2(new_n928), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n933), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n917), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n941), .A2(KEYINPUT53), .A3(new_n928), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n935), .B1(KEYINPUT54), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n907), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(G952), .A2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n865), .B1(new_n945), .B2(new_n946), .ZN(G75));
  NOR2_X1   g761(.A1(new_n320), .A2(G952), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(G210), .A2(G902), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n940), .B2(new_n942), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n429), .A2(new_n430), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(new_n445), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT120), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT55), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n955), .A2(KEYINPUT56), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n949), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT56), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT121), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n951), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n931), .B1(new_n926), .B2(new_n927), .ZN(new_n961));
  AOI22_X1  g775(.A1(new_n930), .A2(new_n933), .B1(new_n941), .B2(new_n961), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n962), .A2(KEYINPUT121), .A3(new_n950), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n955), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT122), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT122), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n955), .C1(new_n960), .C2(new_n963), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n957), .B1(new_n965), .B2(new_n967), .ZN(G51));
  XNOR2_X1  g782(.A(new_n962), .B(KEYINPUT54), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n503), .B(KEYINPUT57), .Z(new_n970));
  OAI21_X1  g784(.A(new_n689), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OR3_X1    g785(.A1(new_n962), .A2(new_n502), .A3(new_n848), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n948), .B1(new_n971), .B2(new_n972), .ZN(G54));
  NOR2_X1   g787(.A1(new_n962), .A2(new_n502), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(KEYINPUT58), .A3(G475), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n975), .A2(new_n620), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n620), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n948), .ZN(G60));
  NAND2_X1  g792(.A1(new_n671), .A2(new_n672), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT123), .Z(new_n980));
  XNOR2_X1  g794(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n981));
  NAND2_X1  g795(.A1(G478), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n980), .B1(new_n944), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n980), .A2(new_n983), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n949), .B1(new_n969), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(G63));
  NAND2_X1  g801(.A1(G217), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT60), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n943), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n948), .B1(new_n991), .B2(new_n654), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n993));
  AOI21_X1  g807(.A(KEYINPUT61), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n943), .A2(new_n706), .A3(new_n990), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n992), .B(new_n995), .C1(new_n993), .C2(KEYINPUT61), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(G66));
  NAND2_X1  g813(.A1(new_n916), .A2(new_n911), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n320), .ZN(new_n1001));
  OAI21_X1  g815(.A(G953), .B1(new_n377), .B2(new_n440), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT126), .Z(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n952), .B1(G898), .B2(new_n320), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(G69));
  NAND2_X1  g820(.A1(new_n923), .A2(new_n795), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT127), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n749), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1012));
  INV_X1    g826(.A(new_n909), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1013), .A2(new_n727), .A3(new_n812), .ZN(new_n1014));
  AOI22_X1  g828(.A1(new_n858), .A2(new_n859), .B1(new_n797), .B2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n855), .A2(new_n1011), .A3(new_n1012), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n320), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n309), .A2(new_n285), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1018), .B(new_n607), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1019), .B1(G900), .B2(G953), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n854), .A2(new_n797), .A3(new_n715), .A4(new_n786), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n860), .A2(new_n819), .A3(new_n1022), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n855), .A2(new_n1023), .A3(new_n817), .A4(new_n1009), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1021), .B1(new_n1024), .B2(G953), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n320), .B1(G227), .B2(G900), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1027), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1020), .A2(new_n1029), .A3(new_n1025), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1028), .A2(new_n1030), .ZN(G72));
  NAND2_X1  g845(.A1(G472), .A2(G902), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n1032), .B(KEYINPUT63), .Z(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(new_n1024), .B2(new_n1000), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n948), .B1(new_n1034), .B2(new_n352), .ZN(new_n1035));
  INV_X1    g849(.A(new_n352), .ZN(new_n1036));
  AND3_X1   g850(.A1(new_n736), .A2(new_n1036), .A3(new_n1033), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1037), .B1(new_n934), .B2(new_n932), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1033), .B1(new_n1016), .B2(new_n1000), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(new_n737), .ZN(new_n1040));
  AND3_X1   g854(.A1(new_n1035), .A2(new_n1038), .A3(new_n1040), .ZN(G57));
endmodule


