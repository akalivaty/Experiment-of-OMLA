//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n644,
    new_n645, new_n646, new_n649, new_n651, new_n652, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT69), .B1(new_n460), .B2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G101), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT68), .B1(new_n470), .B2(G137), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI211_X1 g048(.A(G137), .B(new_n460), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n465), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT67), .B1(new_n472), .B2(new_n473), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n468), .A2(new_n479), .A3(new_n469), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n478), .A2(new_n480), .A3(G125), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n460), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n477), .A2(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n468), .A2(new_n469), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT70), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n460), .B1(new_n468), .B2(new_n469), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT71), .Z(new_n493));
  NAND2_X1  g068(.A1(new_n470), .A2(G136), .ZN(new_n494));
  NOR2_X1   g069(.A1(G100), .A2(G2105), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT72), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(new_n460), .B2(G112), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n493), .B(new_n494), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  XOR2_X1   g073(.A(new_n498), .B(KEYINPUT73), .Z(G162));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n478), .A2(new_n480), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n460), .A2(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT74), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(G102), .A2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(G114), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G2105), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n508), .A2(new_n510), .A3(new_n511), .A4(G2104), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NOR3_X1   g088(.A1(new_n503), .A2(new_n500), .A3(G2105), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n488), .A2(G126), .B1(new_n485), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n504), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(G164));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT75), .B1(new_n519), .B2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n520), .A2(new_n523), .B1(KEYINPUT6), .B2(new_n519), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(KEYINPUT5), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT76), .A3(G543), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(new_n529), .B1(KEYINPUT5), .B2(new_n526), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n524), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G50), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n518), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n530), .A2(G62), .ZN(new_n535));
  NAND2_X1  g110(.A1(G75), .A2(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n519), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(KEYINPUT77), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n535), .A2(new_n536), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n524), .A2(new_n530), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G88), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n524), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G50), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n540), .A2(new_n542), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n538), .A2(new_n546), .ZN(G166));
  AND2_X1   g122(.A1(G63), .A2(G651), .ZN(new_n548));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT7), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n549), .A2(KEYINPUT7), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n530), .A2(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n524), .A2(new_n530), .A3(G89), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n524), .A2(G51), .A3(G543), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n552), .A2(new_n553), .A3(new_n554), .A4(KEYINPUT78), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(G168));
  INV_X1    g134(.A(G90), .ZN(new_n560));
  INV_X1    g135(.A(G52), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n560), .A2(new_n531), .B1(new_n532), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n519), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n562), .A2(new_n564), .ZN(G171));
  INV_X1    g140(.A(G81), .ZN(new_n566));
  INV_X1    g141(.A(G43), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n566), .A2(new_n531), .B1(new_n532), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n519), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT79), .ZN(G153));
  NAND4_X1  g148(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT8), .ZN(new_n576));
  NAND4_X1  g151(.A1(G319), .A2(G483), .A3(G661), .A4(new_n576), .ZN(G188));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n526), .A2(KEYINPUT5), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n528), .A2(KEYINPUT76), .A3(G543), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT76), .B1(new_n528), .B2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G65), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(G651), .A2(new_n584), .B1(new_n541), .B2(G91), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT9), .ZN(new_n587));
  INV_X1    g162(.A(G53), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n586), .B(new_n587), .C1(new_n532), .C2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n588), .B1(KEYINPUT80), .B2(KEYINPUT9), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n543), .B(new_n590), .C1(KEYINPUT80), .C2(KEYINPUT9), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n585), .A2(new_n589), .A3(new_n591), .ZN(G299));
  INV_X1    g167(.A(G171), .ZN(G301));
  INV_X1    g168(.A(G168), .ZN(G286));
  INV_X1    g169(.A(G166), .ZN(G303));
  NAND2_X1  g170(.A1(new_n541), .A2(G87), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n543), .A2(G49), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G288));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n600));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g177(.A(G61), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n530), .A2(KEYINPUT81), .A3(G61), .ZN(new_n606));
  AOI211_X1 g181(.A(new_n600), .B(new_n519), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n604), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n608), .A2(new_n606), .A3(new_n601), .ZN(new_n609));
  AOI21_X1  g184(.A(KEYINPUT82), .B1(new_n609), .B2(G651), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n524), .A2(G48), .A3(G543), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n524), .A2(new_n530), .A3(G86), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n611), .A2(new_n612), .A3(new_n615), .ZN(G305));
  NAND2_X1  g191(.A1(G72), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G60), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n582), .B2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n519), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(new_n619), .ZN(new_n622));
  AOI22_X1  g197(.A1(G47), .A2(new_n543), .B1(new_n541), .B2(G85), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(G290));
  NAND2_X1  g199(.A1(G301), .A2(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n543), .A2(KEYINPUT86), .ZN(new_n626));
  INV_X1    g201(.A(G54), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n532), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(G79), .A2(G543), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT87), .B(G66), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n582), .B2(new_n631), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n626), .A2(new_n629), .B1(new_n632), .B2(G651), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT85), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n541), .A2(new_n634), .A3(G92), .ZN(new_n635));
  INV_X1    g210(.A(G92), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT85), .B1(new_n531), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n635), .A2(KEYINPUT10), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(KEYINPUT10), .B1(new_n635), .B2(new_n637), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n625), .B1(new_n641), .B2(G868), .ZN(G284));
  OAI21_X1  g217(.A(new_n625), .B1(new_n641), .B2(G868), .ZN(G321));
  INV_X1    g218(.A(G868), .ZN(new_n644));
  NOR2_X1   g219(.A1(G286), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G299), .B(KEYINPUT88), .Z(new_n646));
  AOI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(new_n644), .ZN(G297));
  XOR2_X1   g222(.A(G297), .B(KEYINPUT89), .Z(G280));
  INV_X1    g223(.A(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n641), .B1(new_n649), .B2(G860), .ZN(G148));
  NAND2_X1  g225(.A1(new_n641), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G868), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(G868), .B2(new_n571), .ZN(G323));
  XNOR2_X1  g228(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g229(.A1(new_n478), .A2(new_n480), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n461), .B(new_n462), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT12), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT13), .ZN(new_n659));
  INV_X1    g234(.A(G2100), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n491), .A2(G123), .ZN(new_n663));
  OAI21_X1  g238(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n664));
  INV_X1    g239(.A(G111), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n664), .B1(new_n665), .B2(G2105), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(G135), .B2(new_n470), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(G2096), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n661), .A2(new_n662), .A3(new_n669), .ZN(G156));
  INV_X1    g245(.A(KEYINPUT14), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2427), .B(G2438), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2430), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT15), .B(G2435), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n674), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2451), .B(G2454), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT16), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1341), .B(G1348), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n676), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2443), .B(G2446), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(new_n684), .A3(G14), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT90), .ZN(G401));
  XOR2_X1   g261(.A(G2072), .B(G2078), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT91), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT17), .ZN(new_n689));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  XNOR2_X1  g265(.A(G2084), .B(G2090), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n688), .B2(new_n690), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n689), .B2(new_n690), .ZN(new_n694));
  INV_X1    g269(.A(new_n690), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(new_n691), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT18), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n692), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G2096), .B(G2100), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G227));
  XOR2_X1   g276(.A(G1971), .B(G1976), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT19), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1956), .B(G2474), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1961), .B(G1966), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n708));
  XOR2_X1   g283(.A(new_n707), .B(new_n708), .Z(new_n709));
  AND2_X1   g284(.A1(new_n704), .A2(new_n705), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT93), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n703), .A2(new_n710), .A3(new_n706), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1991), .B(G1996), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(G1981), .B(G1986), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(G229));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G23), .ZN(new_n723));
  INV_X1    g298(.A(G288), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n722), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT33), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1976), .ZN(new_n727));
  MUX2_X1   g302(.A(G6), .B(G305), .S(G16), .Z(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT32), .B(G1981), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n722), .A2(G22), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G166), .B2(new_n722), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G1971), .Z(new_n734));
  NAND4_X1  g309(.A1(new_n727), .A2(new_n730), .A3(new_n731), .A4(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT34), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT34), .ZN(new_n737));
  INV_X1    g312(.A(G24), .ZN(new_n738));
  OR3_X1    g313(.A1(new_n738), .A2(KEYINPUT95), .A3(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT95), .B1(new_n738), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G290), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n722), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G1986), .Z(new_n743));
  INV_X1    g318(.A(G29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G25), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n491), .A2(G119), .ZN(new_n746));
  OAI21_X1  g321(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n747));
  INV_X1    g322(.A(G107), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G2105), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G131), .B2(new_n470), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n745), .B1(new_n752), .B2(new_n744), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT35), .B(G1991), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT94), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n753), .B(new_n755), .ZN(new_n756));
  AND3_X1   g331(.A1(new_n743), .A2(KEYINPUT96), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n736), .A2(new_n737), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NOR2_X1   g336(.A1(G29), .A2(G35), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G162), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT29), .B(G2090), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G16), .A2(G21), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G168), .B2(G16), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT103), .B(G1966), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT30), .B(G28), .ZN(new_n771));
  OR2_X1    g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  NAND2_X1  g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n771), .A2(new_n744), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G164), .A2(new_n744), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G27), .B2(new_n744), .ZN(new_n776));
  INV_X1    g351(.A(G2078), .ZN(new_n777));
  OAI221_X1 g352(.A(new_n774), .B1(new_n744), .B2(new_n668), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT98), .B(KEYINPUT28), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n744), .A2(G26), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n491), .A2(G128), .ZN(new_n782));
  OAI21_X1  g357(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n783));
  INV_X1    g358(.A(G116), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G2105), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G140), .B2(new_n470), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n781), .B1(new_n787), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT99), .B(G2067), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G16), .A2(G19), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n571), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT97), .B(G1341), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n722), .A2(G5), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G171), .B2(new_n722), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G1961), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n790), .A2(new_n794), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  AOI211_X1 g374(.A(new_n778), .B(new_n799), .C1(new_n777), .C2(new_n776), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n655), .A2(G127), .ZN(new_n801));
  NAND2_X1  g376(.A1(G115), .A2(G2104), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n460), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT25), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n470), .A2(G139), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n803), .B2(new_n804), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n806), .A2(new_n814), .A3(new_n744), .ZN(new_n815));
  INV_X1    g390(.A(G33), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n744), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(G2072), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n744), .A2(G32), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT102), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n656), .A2(G105), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT101), .ZN(new_n822));
  NAND3_X1  g397(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT26), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  AOI22_X1  g401(.A1(G141), .A2(new_n470), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n487), .A2(new_n490), .ZN(new_n828));
  INV_X1    g403(.A(G129), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n820), .B1(new_n822), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n821), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n491), .A2(G129), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n833), .A2(KEYINPUT102), .A3(new_n834), .A4(new_n827), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n819), .B1(new_n837), .B2(new_n744), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT27), .B(G1996), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n818), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n838), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n842), .A2(new_n839), .B1(G2072), .B2(new_n817), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n722), .A2(G20), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT23), .ZN(new_n845));
  INV_X1    g420(.A(G299), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n722), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G1956), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT24), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n744), .B1(new_n849), .B2(G34), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n849), .B2(G34), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G160), .B2(G29), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(G2084), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(G2084), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(G1961), .B2(new_n797), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n848), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n800), .A2(new_n841), .A3(new_n843), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n763), .A2(new_n764), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n722), .A2(G4), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n641), .B2(new_n722), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G1348), .ZN(new_n861));
  NOR4_X1   g436(.A1(new_n770), .A2(new_n857), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n760), .A2(new_n761), .A3(new_n862), .ZN(G150));
  INV_X1    g438(.A(G150), .ZN(G311));
  XNOR2_X1  g439(.A(KEYINPUT105), .B(G860), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n641), .A2(G559), .ZN(new_n867));
  XOR2_X1   g442(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  AOI22_X1  g444(.A1(G55), .A2(new_n543), .B1(new_n541), .B2(G93), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n519), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n571), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n869), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n866), .B1(new_n875), .B2(KEYINPUT39), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(KEYINPUT39), .B2(new_n875), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n872), .A2(new_n866), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT37), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(G145));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  INV_X1    g458(.A(G118), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n883), .B1(new_n884), .B2(G2105), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(G142), .B2(new_n470), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n491), .A2(G130), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n888), .A2(KEYINPUT106), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(KEYINPUT106), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n806), .A2(new_n814), .A3(new_n787), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n782), .A2(new_n786), .ZN(new_n893));
  INV_X1    g468(.A(new_n813), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n801), .A2(new_n802), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(G2105), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n896), .B2(KEYINPUT100), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n893), .B1(new_n897), .B2(new_n805), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n891), .B1(new_n892), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n888), .B(KEYINPUT106), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n886), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n787), .B1(new_n806), .B2(new_n814), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n897), .A2(new_n805), .A3(new_n893), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n836), .B(new_n516), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n836), .B(G164), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n904), .A3(new_n899), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n751), .B(KEYINPUT107), .Z(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(new_n658), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n907), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n911), .B1(new_n907), .B2(new_n909), .ZN(new_n915));
  OAI21_X1  g490(.A(G160), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n907), .A2(new_n909), .ZN(new_n917));
  INV_X1    g492(.A(new_n911), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G160), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n919), .A2(new_n913), .A3(new_n920), .A4(new_n912), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(G162), .B(new_n668), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n882), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n923), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n925), .B1(new_n916), .B2(new_n921), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n881), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n922), .A2(new_n923), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n921), .A3(new_n916), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT40), .A4(new_n882), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n927), .A2(new_n930), .ZN(G395));
  NAND2_X1  g506(.A1(new_n641), .A2(new_n846), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  OAI21_X1  g508(.A(G299), .B1(new_n639), .B2(new_n640), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT109), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n873), .B(new_n651), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n932), .A2(new_n934), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n942), .B1(new_n944), .B2(new_n939), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n946));
  NOR2_X1   g521(.A1(G305), .A2(new_n741), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(G166), .B(G288), .ZN(new_n949));
  NAND2_X1  g524(.A1(G305), .A2(new_n741), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n948), .B2(new_n950), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n946), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n946), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n872), .A2(new_n644), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(G295));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n958), .ZN(G331));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  NOR2_X1   g537(.A1(G286), .A2(G301), .ZN(new_n963));
  NOR2_X1   g538(.A1(G168), .A2(G171), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n873), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n568), .A2(new_n570), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n872), .B(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n964), .B2(new_n963), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n943), .A2(KEYINPUT41), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n940), .B1(new_n971), .B2(new_n935), .ZN(new_n972));
  INV_X1    g547(.A(new_n941), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n970), .A2(new_n943), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G37), .B1(new_n977), .B2(new_n953), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n951), .A2(new_n952), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n974), .A2(new_n979), .A3(new_n976), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n962), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n970), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n938), .B2(new_n941), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n983), .A2(new_n953), .A3(new_n975), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n971), .A2(new_n935), .B1(new_n966), .B2(new_n969), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n975), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n882), .B1(new_n986), .B2(new_n979), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n984), .A2(new_n987), .A3(KEYINPUT43), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n961), .B1(new_n981), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n983), .A2(new_n975), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT43), .B1(new_n991), .B2(new_n979), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n961), .B1(new_n992), .B2(new_n978), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT43), .B1(new_n984), .B2(new_n987), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n953), .B1(new_n983), .B2(new_n975), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n996), .A2(new_n980), .A3(new_n962), .A4(new_n882), .ZN(new_n997));
  AND4_X1   g572(.A1(new_n990), .A2(new_n994), .A3(KEYINPUT44), .A4(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n989), .B1(new_n995), .B2(new_n998), .ZN(G397));
  NAND3_X1  g574(.A1(new_n470), .A2(KEYINPUT68), .A3(G137), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n474), .A2(new_n475), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n1000), .A2(new_n1001), .B1(new_n656), .B2(G101), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n481), .A2(new_n482), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1002), .B(G40), .C1(new_n1003), .C2(new_n460), .ZN(new_n1004));
  INV_X1    g579(.A(G1384), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n502), .A2(new_n503), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n488), .A2(G126), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n485), .A2(new_n514), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n513), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1005), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n724), .A2(G1976), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT52), .ZN(new_n1016));
  INV_X1    g591(.A(G1976), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(G288), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1013), .A2(new_n1014), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  INV_X1    g597(.A(new_n612), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT116), .B(G86), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n541), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1022), .B1(new_n611), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n609), .A2(G651), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n600), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n609), .A2(KEYINPUT82), .A3(G651), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1023), .A2(G1981), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n615), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n611), .A2(KEYINPUT115), .A3(new_n615), .A4(new_n1030), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1026), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1013), .B1(new_n1035), .B2(KEYINPUT49), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1026), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1037), .A2(KEYINPUT49), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1021), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1010), .A2(KEYINPUT50), .ZN(new_n1041));
  INV_X1    g616(.A(G40), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n477), .A2(new_n483), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n516), .A2(new_n1044), .A3(new_n1005), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT114), .B1(new_n1046), .B2(G2090), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1044), .B1(new_n516), .B2(new_n1005), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(new_n1004), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n1050));
  INV_X1    g625(.A(G2090), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1045), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1010), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n516), .A2(KEYINPUT45), .A3(new_n1005), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1043), .A3(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT113), .B(G1971), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1047), .A2(new_n1052), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n538), .A2(new_n546), .A3(G8), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(G8), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1046), .A2(KEYINPUT117), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1049), .A2(new_n1065), .A3(new_n1045), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(new_n1066), .A3(new_n1051), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1012), .B1(new_n1067), .B2(new_n1058), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1063), .B1(new_n1068), .B2(new_n1062), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1053), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1005), .B(new_n1070), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n513), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1384), .B1(new_n1072), .B2(new_n504), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1043), .B(new_n1071), .C1(new_n1073), .C2(KEYINPUT45), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n768), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT118), .B(G2084), .Z(new_n1076));
  NAND4_X1  g651(.A1(new_n1041), .A2(new_n1043), .A3(new_n1045), .A4(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1012), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G168), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1040), .A2(new_n1069), .A3(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT119), .B1(new_n1080), .B2(KEYINPUT63), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT63), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1035), .A2(KEYINPUT49), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n1013), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1062), .ZN(new_n1089));
  AOI21_X1  g664(.A(G2090), .B1(new_n1046), .B2(KEYINPUT117), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1090), .A2(new_n1066), .B1(new_n1057), .B2(new_n1056), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1089), .B1(new_n1091), .B2(new_n1012), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1088), .A2(new_n1021), .A3(new_n1063), .A4(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1082), .B(new_n1083), .C1(new_n1093), .C2(new_n1079), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1059), .A2(G8), .A3(new_n1062), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1095), .A2(new_n1083), .A3(new_n1079), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1013), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1020), .B1(new_n1098), .B2(new_n1087), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1059), .A2(G8), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1096), .B(new_n1099), .C1(new_n1062), .C2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1081), .A2(new_n1094), .A3(new_n1101), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT120), .B(G1956), .Z(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1046), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n591), .A2(new_n589), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n584), .A2(G651), .ZN(new_n1108));
  INV_X1    g683(.A(G91), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(new_n531), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1106), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n585), .A2(KEYINPUT57), .A3(new_n589), .A4(new_n591), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1054), .A2(new_n1043), .A3(new_n1055), .A4(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1105), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G1348), .ZN(new_n1117));
  INV_X1    g692(.A(G2067), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1046), .A2(new_n1117), .B1(new_n1011), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n641), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1113), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1103), .B1(new_n1049), .B2(new_n1045), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1115), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1116), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1996), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1054), .A2(new_n1129), .A3(new_n1043), .A4(new_n1055), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT58), .B(G1341), .Z(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1128), .B1(new_n1133), .B2(new_n571), .ZN(new_n1134));
  AOI211_X1 g709(.A(new_n967), .B(new_n1127), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1113), .B1(new_n1105), .B2(new_n1115), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT61), .B1(new_n1116), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1105), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1125), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1136), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1119), .A2(KEYINPUT60), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT122), .B1(new_n1119), .B2(KEYINPUT60), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(new_n1120), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1011), .A2(new_n1118), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n516), .A2(new_n1044), .A3(new_n1005), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1147), .A2(new_n1048), .A3(new_n1004), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT60), .B(new_n1146), .C1(new_n1148), .C2(G1348), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1119), .A2(KEYINPUT122), .A3(KEYINPUT60), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n641), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1145), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1126), .B1(new_n1142), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1056), .A2(G2078), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT53), .ZN(new_n1158));
  INV_X1    g733(.A(G1961), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1157), .A2(new_n1158), .B1(new_n1159), .B2(new_n1046), .ZN(new_n1160));
  XOR2_X1   g735(.A(G171), .B(KEYINPUT54), .Z(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(KEYINPUT53), .B2(new_n1156), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1046), .A2(new_n1159), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n1164));
  OAI221_X1 g739(.A(new_n1163), .B1(new_n1074), .B2(new_n1164), .C1(new_n1156), .C2(KEYINPUT53), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1160), .A2(new_n1162), .B1(new_n1165), .B2(new_n1161), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT51), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT123), .B1(G168), .B2(new_n1012), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n557), .A2(new_n1169), .A3(G8), .A4(new_n558), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1167), .B1(new_n1078), .B2(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1148), .A2(new_n1076), .B1(new_n768), .B2(new_n1074), .ZN(new_n1174));
  OAI211_X1 g749(.A(KEYINPUT51), .B(new_n1173), .C1(new_n1174), .C2(new_n1012), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1171), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1172), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1166), .A2(new_n1178), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1155), .A2(new_n1093), .A3(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(G288), .A2(G1976), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1088), .A2(new_n1181), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1182));
  OAI22_X1  g757(.A1(new_n1182), .A2(new_n1097), .B1(new_n1040), .B2(new_n1063), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n1185));
  AOI21_X1  g760(.A(KEYINPUT124), .B1(new_n1178), .B2(KEYINPUT62), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1178), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1067), .A2(new_n1058), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1062), .B1(new_n1190), .B2(G8), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1191), .A2(new_n1095), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1172), .A2(new_n1175), .A3(new_n1193), .A4(new_n1177), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1165), .A2(G171), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1099), .A2(new_n1192), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1185), .B1(new_n1189), .B2(new_n1197), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1178), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1199), .A2(new_n1186), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1200), .A2(KEYINPUT125), .A3(new_n1196), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1102), .B(new_n1184), .C1(new_n1198), .C2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1054), .A2(new_n1004), .ZN(new_n1203));
  XOR2_X1   g778(.A(new_n1203), .B(KEYINPUT112), .Z(new_n1204));
  NAND2_X1  g779(.A1(new_n893), .A2(new_n1118), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n787), .A2(G2067), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1207), .B1(new_n836), .B2(G1996), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1204), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n837), .A2(new_n1129), .A3(new_n1203), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n751), .B(new_n755), .ZN(new_n1211));
  OAI211_X1 g786(.A(new_n1209), .B(new_n1210), .C1(new_n1204), .C2(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g787(.A(G290), .B(G1986), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1212), .B1(new_n1203), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1202), .A2(new_n1214), .ZN(new_n1215));
  NAND4_X1  g790(.A1(new_n1209), .A2(new_n755), .A3(new_n752), .A4(new_n1210), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1204), .B1(new_n1216), .B2(new_n1205), .ZN(new_n1217));
  AND2_X1   g792(.A1(new_n1217), .A2(KEYINPUT126), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1217), .A2(KEYINPUT126), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1203), .A2(new_n1129), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n1220), .B(KEYINPUT46), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1207), .A2(new_n836), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1221), .B1(new_n1204), .B2(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n1223), .B(KEYINPUT47), .ZN(new_n1224));
  NOR4_X1   g799(.A1(G290), .A2(new_n1054), .A3(G1986), .A4(new_n1004), .ZN(new_n1225));
  XOR2_X1   g800(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1226));
  XNOR2_X1  g801(.A(new_n1225), .B(new_n1226), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1224), .B1(new_n1212), .B2(new_n1227), .ZN(new_n1228));
  NOR3_X1   g803(.A1(new_n1218), .A2(new_n1219), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1215), .A2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g805(.A1(new_n928), .A2(new_n882), .A3(new_n929), .ZN(new_n1232));
  INV_X1    g806(.A(G319), .ZN(new_n1233));
  NOR3_X1   g807(.A1(G401), .A2(new_n1233), .A3(G227), .ZN(new_n1234));
  AND2_X1   g808(.A1(new_n720), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g809(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g810(.A1(new_n981), .A2(new_n988), .ZN(new_n1237));
  NOR2_X1   g811(.A1(new_n1236), .A2(new_n1237), .ZN(G308));
  OAI211_X1 g812(.A(new_n1232), .B(new_n1235), .C1(new_n981), .C2(new_n988), .ZN(G225));
endmodule


