//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1253, new_n1254, new_n1255;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  OR2_X1    g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n460), .B(new_n461), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G137), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n465), .A2(G136), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n459), .A2(G114), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OR2_X1    g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n484), .A2(new_n486), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n483), .A2(new_n487), .B1(new_n474), .B2(G126), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n459), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n468), .A2(new_n493), .A3(G138), .A4(new_n459), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT71), .B1(new_n498), .B2(G543), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT5), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n499), .A2(new_n502), .B1(new_n498), .B2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n503), .A2(G62), .ZN(new_n504));
  AND2_X1   g079(.A1(G75), .A2(G543), .ZN(new_n505));
  OAI211_X1 g080(.A(KEYINPUT72), .B(G651), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n505), .B1(new_n503), .B2(G62), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n511), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT70), .A3(G651), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n512), .A2(new_n514), .B1(KEYINPUT6), .B2(new_n509), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n503), .A2(new_n515), .A3(G88), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(G50), .A3(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n506), .A2(new_n510), .A3(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND2_X1  g095(.A1(new_n503), .A2(new_n515), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n515), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n503), .A2(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n523), .A2(new_n526), .A3(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(new_n522), .A2(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OAI221_X1 g110(.A(new_n533), .B1(new_n534), .B2(new_n524), .C1(new_n509), .C2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  AOI22_X1  g112(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n509), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n521), .A2(new_n540), .B1(new_n524), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  INV_X1    g123(.A(G65), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n499), .A2(new_n502), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n498), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT73), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n503), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n549), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g131(.A1(G78), .A2(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n524), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n515), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n560), .A2(new_n562), .B1(G91), .B2(new_n522), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n558), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND3_X1  g140(.A1(new_n503), .A2(new_n515), .A3(G87), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n515), .A2(G49), .A3(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G74), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n509), .B1(new_n552), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(KEYINPUT74), .ZN(new_n572));
  OAI211_X1 g147(.A(KEYINPUT74), .B(G651), .C1(new_n503), .C2(G74), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n569), .B1(new_n572), .B2(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(new_n503), .A2(G61), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n503), .A2(KEYINPUT75), .A3(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n521), .A2(new_n583), .B1(new_n524), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n509), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n521), .A2(new_n590), .B1(new_n524), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT76), .Z(new_n596));
  NAND2_X1  g171(.A1(new_n553), .A2(new_n555), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n509), .ZN(new_n599));
  XNOR2_X1  g174(.A(KEYINPUT77), .B(KEYINPUT10), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n522), .A2(G92), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n600), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n521), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n601), .A2(new_n604), .B1(G54), .B2(new_n525), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n596), .B1(G868), .B2(new_n607), .ZN(G284));
  OAI21_X1  g183(.A(new_n596), .B1(G868), .B2(new_n607), .ZN(G321));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(G299), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n610), .B2(G168), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(new_n610), .B2(G168), .ZN(G280));
  XNOR2_X1  g188(.A(KEYINPUT78), .B(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(G860), .B2(new_n614), .ZN(G148));
  OAI21_X1  g190(.A(KEYINPUT80), .B1(new_n543), .B2(G868), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n599), .A2(new_n605), .A3(new_n614), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  MUX2_X1   g197(.A(KEYINPUT80), .B(new_n616), .S(new_n622), .Z(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g199(.A1(new_n459), .A2(G2104), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n468), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n465), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n474), .A2(G123), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n631), .A3(new_n637), .ZN(G156));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n644), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n652), .A3(G14), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g230(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT81), .A4(G14), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT82), .ZN(new_n659));
  NOR2_X1   g234(.A1(G2072), .A2(G2078), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n442), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n661), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(KEYINPUT17), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n662), .C1(new_n659), .C2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n662), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n659), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n689), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n676), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(new_n676), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n694), .A2(new_n690), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n693), .A2(new_n696), .A3(new_n698), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(KEYINPUT95), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G21), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G168), .B2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G1966), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT92), .ZN(new_n712));
  NOR2_X1   g287(.A1(G5), .A2(G16), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT93), .Z(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G301), .B2(new_n705), .ZN(new_n715));
  INV_X1    g290(.A(G1961), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT94), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n709), .A2(new_n710), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT31), .B(G11), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT30), .B(G28), .Z(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n636), .A2(new_n723), .ZN(new_n724));
  OAI221_X1 g299(.A(new_n721), .B1(G29), .B2(new_n722), .C1(new_n724), .C2(KEYINPUT91), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(KEYINPUT91), .B2(new_n724), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n719), .A2(new_n720), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n704), .B1(new_n712), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT92), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n711), .B(new_n729), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n720), .A2(new_n726), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n730), .A2(new_n731), .A3(KEYINPUT95), .A4(new_n719), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n723), .A2(G33), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n468), .A2(G127), .ZN(new_n734));
  NAND2_X1  g309(.A1(G115), .A2(G2104), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n459), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n465), .A2(G139), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT25), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n736), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n733), .B1(new_n741), .B2(new_n723), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2072), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n723), .A2(G32), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT26), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G129), .B2(new_n474), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n465), .A2(G141), .B1(G105), .B2(new_n625), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n744), .B1(new_n750), .B2(new_n723), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT27), .B(G1996), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n743), .B(new_n753), .C1(new_n716), .C2(new_n715), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n705), .A2(G19), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n543), .B2(new_n705), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1341), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n723), .A2(G26), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT28), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n474), .A2(G128), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT89), .ZN(new_n761));
  OAI21_X1  g336(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n762));
  INV_X1    g337(.A(G116), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(G2105), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n465), .B2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n759), .B1(new_n766), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2067), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n723), .A2(G35), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n723), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT29), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G2090), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n757), .A2(new_n769), .A3(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G34), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n775), .A2(KEYINPUT24), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(KEYINPUT24), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n723), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G160), .B2(new_n723), .ZN(new_n779));
  INV_X1    g354(.A(G2084), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(G164), .A2(G29), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G27), .B2(G29), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT96), .B(G2078), .Z(new_n784));
  OAI21_X1  g359(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n783), .B2(new_n784), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n754), .A2(new_n774), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G4), .A2(G16), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n607), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT88), .B(G1348), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n772), .A2(G2090), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT97), .Z(new_n793));
  NOR3_X1   g368(.A1(new_n787), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n705), .A2(G20), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT23), .Z(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G299), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT98), .ZN(new_n798));
  INV_X1    g373(.A(G1956), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n728), .A2(new_n732), .A3(new_n794), .A4(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT86), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n582), .A2(G16), .A3(new_n586), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G6), .B2(G16), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT32), .B(G1981), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n804), .A2(new_n806), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n807), .A2(KEYINPUT85), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(G166), .A2(G16), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G16), .B2(G22), .ZN(new_n812));
  INV_X1    g387(.A(G1971), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n811), .B(G1971), .C1(G16), .C2(G22), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n705), .A2(G23), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n571), .A2(KEYINPUT74), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n568), .B1(new_n817), .B2(new_n573), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n816), .B1(new_n818), .B2(new_n705), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT33), .B(G1976), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n819), .A2(new_n821), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n814), .A2(new_n815), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(KEYINPUT85), .B1(new_n807), .B2(new_n808), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n810), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT34), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n802), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n723), .A2(G25), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n465), .A2(G131), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT83), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n832));
  INV_X1    g407(.A(G107), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(G2105), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G119), .B2(new_n474), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT84), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n829), .B1(new_n837), .B2(new_n723), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT35), .B(G1991), .Z(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n705), .A2(G24), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n593), .B2(new_n705), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(G1986), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(G1986), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n841), .A2(new_n842), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n826), .B2(new_n827), .ZN(new_n848));
  INV_X1    g423(.A(new_n824), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(new_n809), .ZN(new_n850));
  OAI211_X1 g425(.A(KEYINPUT86), .B(KEYINPUT34), .C1(new_n850), .C2(new_n825), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n828), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n801), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n828), .A2(new_n848), .A3(new_n851), .A4(new_n854), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT99), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n852), .A2(new_n856), .ZN(new_n860));
  INV_X1    g435(.A(new_n801), .ZN(new_n861));
  AND4_X1   g436(.A1(KEYINPUT99), .A2(new_n860), .A3(new_n861), .A4(new_n858), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n859), .A2(new_n862), .ZN(G311));
  NAND2_X1  g438(.A1(new_n857), .A2(new_n858), .ZN(G150));
  AOI22_X1  g439(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(new_n509), .ZN(new_n866));
  INV_X1    g441(.A(G93), .ZN(new_n867));
  INV_X1    g442(.A(G55), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n521), .A2(new_n867), .B1(new_n524), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G860), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT37), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n607), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT38), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n866), .A2(new_n869), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n543), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n543), .A2(new_n875), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n874), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(G860), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n883), .A2(KEYINPUT100), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT100), .B1(new_n883), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n872), .B1(new_n885), .B2(new_n886), .ZN(G145));
  XNOR2_X1  g462(.A(KEYINPUT102), .B(G37), .ZN(new_n888));
  INV_X1    g463(.A(new_n627), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n836), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n831), .A2(new_n627), .A3(new_n835), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n741), .B(new_n749), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n766), .A2(new_n496), .ZN(new_n897));
  NAND3_X1  g472(.A1(G164), .A2(new_n761), .A3(new_n765), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n474), .A2(G130), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(KEYINPUT101), .Z(new_n901));
  OAI21_X1  g476(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n902));
  INV_X1    g477(.A(G118), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(G2105), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n465), .A2(G142), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n901), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n899), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n899), .A2(new_n907), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n896), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n636), .B(new_n478), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(G160), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n894), .A2(new_n908), .A3(new_n909), .A4(new_n895), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n911), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n888), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT103), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n919), .B(new_n888), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n923));
  XNOR2_X1  g498(.A(G305), .B(new_n593), .ZN(new_n924));
  XNOR2_X1  g499(.A(G303), .B(G288), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n927));
  XNOR2_X1  g502(.A(G305), .B(G290), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(new_n925), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n923), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n606), .A2(G299), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n599), .A2(new_n558), .A3(new_n563), .A4(new_n605), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n619), .A2(new_n620), .A3(new_n879), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n879), .B1(new_n619), .B2(new_n620), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n940), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n938), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT41), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n934), .A2(new_n944), .A3(new_n935), .ZN(new_n945));
  XOR2_X1   g520(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n934), .B2(new_n935), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n941), .B1(new_n943), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n933), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n932), .B(new_n941), .C1(new_n943), .C2(new_n948), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n931), .A2(new_n927), .A3(new_n923), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(G868), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n875), .A2(G868), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(G295));
  AOI21_X1  g533(.A(new_n952), .B1(new_n933), .B2(new_n949), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n610), .B1(new_n959), .B2(new_n951), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT106), .B1(new_n960), .B2(new_n956), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n955), .A2(new_n962), .A3(new_n957), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(G331));
  NAND2_X1  g539(.A1(new_n879), .A2(G301), .ZN(new_n965));
  OAI21_X1  g540(.A(G171), .B1(new_n877), .B2(new_n878), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(G168), .A3(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n877), .A2(G171), .A3(new_n878), .ZN(new_n968));
  INV_X1    g543(.A(new_n543), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n870), .ZN(new_n970));
  AOI21_X1  g545(.A(G301), .B1(new_n970), .B2(new_n876), .ZN(new_n971));
  OAI21_X1  g546(.A(G286), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n937), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n967), .B(new_n972), .C1(new_n945), .C2(new_n947), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n926), .ZN(new_n977));
  INV_X1    g552(.A(G37), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(new_n975), .A3(new_n929), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n936), .A2(new_n946), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n936), .A2(new_n944), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n974), .B1(new_n984), .B2(new_n973), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n926), .ZN(new_n986));
  AND4_X1   g561(.A1(KEYINPUT43), .A2(new_n986), .A3(new_n888), .A4(new_n979), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT44), .B1(new_n981), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n986), .A2(new_n989), .A3(new_n888), .A4(new_n979), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n980), .B2(new_n989), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n988), .A2(new_n993), .ZN(G397));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n492), .A2(new_n494), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n483), .A2(new_n487), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n474), .A2(G126), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n995), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n469), .A2(new_n470), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G2105), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1004), .A2(G40), .A3(new_n466), .A4(new_n462), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT108), .ZN(new_n1007));
  INV_X1    g582(.A(G1996), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n1009), .B(KEYINPUT107), .Z(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n750), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n766), .B(G2067), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n750), .A2(new_n1008), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1007), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1015), .A2(new_n837), .A3(new_n839), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n766), .A2(G2067), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1007), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1007), .B1(new_n749), .B2(new_n1012), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1010), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1010), .A2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT47), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n836), .B(new_n840), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1007), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G290), .A2(G1986), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n1006), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT48), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1015), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1018), .A2(new_n1024), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  INV_X1    g607(.A(G40), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n467), .A2(new_n471), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n488), .B2(new_n495), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(G1976), .B(new_n569), .C1(new_n572), .C2(new_n574), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(G288), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT112), .B1(new_n1042), .B2(KEYINPUT52), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n1044), .B(new_n1045), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1041), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n576), .A2(new_n577), .B1(G73), .B2(G543), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n509), .B1(new_n1048), .B2(new_n579), .ZN(new_n1049));
  OAI21_X1  g624(.A(G1981), .B1(new_n1049), .B2(new_n585), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n582), .A2(new_n1051), .A3(new_n586), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1052), .A3(KEYINPUT49), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT113), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1050), .A2(new_n1052), .A3(new_n1055), .A4(KEYINPUT49), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT49), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1036), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1047), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1005), .B1(new_n1000), .B2(KEYINPUT50), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1035), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT110), .B(G2090), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1034), .B1(new_n1035), .B2(KEYINPUT45), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1001), .B(G1384), .C1(new_n488), .C2(new_n495), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n813), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1032), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G303), .A2(G8), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1070), .A2(KEYINPUT111), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT111), .B1(new_n1070), .B2(new_n1075), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n710), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1080), .A2(new_n780), .A3(new_n1034), .A4(new_n1064), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1032), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT63), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(G168), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1035), .A2(KEYINPUT114), .A3(new_n1063), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT114), .B1(new_n1035), .B2(new_n1063), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1062), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1065), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1069), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G8), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1075), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1084), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1061), .B1(new_n1078), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1044), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1042), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1096), .A2(new_n1097), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1005), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1035), .A2(KEYINPUT45), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1966), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1034), .B1(new_n1035), .B2(new_n1063), .ZN(new_n1103));
  AOI211_X1 g678(.A(KEYINPUT50), .B(G1384), .C1(new_n488), .C2(new_n495), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1103), .A2(G2084), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(G8), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(G286), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1095), .A2(new_n1098), .A3(new_n1099), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT63), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n818), .A2(new_n1039), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1052), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1036), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1094), .A2(new_n1109), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n1115));
  OAI21_X1  g690(.A(G286), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1079), .A2(new_n1081), .A3(G168), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(G8), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1106), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(KEYINPUT51), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1117), .A2(G8), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT51), .B1(new_n1082), .B2(KEYINPUT122), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1115), .B1(new_n1126), .B2(KEYINPUT62), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  AOI211_X1 g703(.A(KEYINPUT124), .B(new_n1128), .C1(new_n1121), .C2(new_n1125), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(G1971), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT114), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1064), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1103), .B1(new_n1133), .B2(new_n1085), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1131), .B1(new_n1065), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1092), .B1(new_n1135), .B2(new_n1032), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1095), .A2(new_n1136), .A3(new_n1098), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n1078), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1067), .A2(G2078), .A3(new_n1068), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1080), .A2(new_n1034), .A3(new_n1064), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1139), .A2(KEYINPUT53), .B1(new_n1140), .B2(new_n716), .ZN(new_n1141));
  INV_X1    g716(.A(G2078), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1002), .A2(new_n1142), .A3(new_n1101), .A4(new_n1034), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(G301), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1121), .A2(new_n1128), .A3(new_n1125), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1138), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1114), .B1(new_n1130), .B2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(KEYINPUT56), .B(G2072), .Z(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT116), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1100), .A2(new_n1101), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1134), .B2(G1956), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT115), .B1(new_n560), .B2(new_n562), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(KEYINPUT57), .ZN(new_n1155));
  NAND2_X1  g730(.A1(G299), .A2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n558), .B(new_n563), .C1(new_n1154), .C2(KEYINPUT57), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT117), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT117), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1153), .A2(new_n1161), .A3(new_n1158), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1000), .A2(new_n1005), .A3(G2067), .ZN(new_n1164));
  INV_X1    g739(.A(G1348), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1140), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n606), .ZN(new_n1167));
  OAI22_X1  g742(.A1(new_n1163), .A2(new_n1167), .B1(new_n1158), .B2(new_n1153), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1165), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1164), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT60), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n606), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n1166), .B2(KEYINPUT60), .ZN(new_n1175));
  AND4_X1   g750(.A1(new_n1174), .A2(new_n1169), .A3(new_n1170), .A4(KEYINPUT60), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1173), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n607), .B1(new_n1166), .B2(KEYINPUT60), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT121), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1166), .A2(new_n1174), .A3(KEYINPUT60), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1088), .A2(new_n799), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1185), .B1(new_n1186), .B2(new_n1152), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1183), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT120), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT120), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1186), .A2(new_n1190), .A3(new_n1185), .A4(new_n1152), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1189), .A2(KEYINPUT61), .A3(new_n1191), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1182), .B(new_n1188), .C1(new_n1163), .C2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1002), .A2(new_n1008), .A3(new_n1101), .A4(new_n1034), .ZN(new_n1194));
  XOR2_X1   g769(.A(KEYINPUT58), .B(G1341), .Z(new_n1195));
  OAI21_X1  g770(.A(new_n1195), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1194), .A2(KEYINPUT118), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(KEYINPUT118), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n543), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(KEYINPUT119), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT119), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1201), .B(new_n543), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1200), .A2(KEYINPUT59), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT59), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1199), .A2(KEYINPUT119), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1168), .B1(new_n1193), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1140), .A2(new_n716), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1100), .A2(KEYINPUT53), .A3(new_n1142), .A4(new_n1101), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1145), .ZN(new_n1211));
  OAI21_X1  g786(.A(G171), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1141), .A2(G301), .A3(new_n1145), .ZN(new_n1213));
  AOI21_X1  g788(.A(KEYINPUT54), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1214), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1212), .A2(new_n1213), .A3(KEYINPUT54), .ZN(new_n1216));
  NAND4_X1  g791(.A1(new_n1215), .A2(new_n1138), .A3(KEYINPUT123), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT123), .ZN(new_n1218));
  INV_X1    g793(.A(KEYINPUT54), .ZN(new_n1219));
  AND4_X1   g794(.A1(G301), .A2(new_n1145), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1219), .B1(new_n1146), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1124), .B1(new_n1123), .B2(new_n1116), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1122), .B1(new_n1120), .B2(KEYINPUT51), .ZN(new_n1223));
  OAI211_X1 g798(.A(new_n1221), .B(new_n1216), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  INV_X1    g799(.A(new_n1077), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1070), .A2(KEYINPUT111), .A3(new_n1075), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1227), .A2(new_n1061), .A3(new_n1136), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1218), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n1207), .A2(new_n1217), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1149), .A2(new_n1230), .ZN(new_n1231));
  AND2_X1   g806(.A1(G290), .A2(G1986), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1006), .B1(new_n1232), .B2(new_n1027), .ZN(new_n1233));
  NAND4_X1  g808(.A1(new_n1011), .A2(new_n1233), .A3(new_n1014), .A4(new_n1026), .ZN(new_n1234));
  XNOR2_X1  g809(.A(new_n1234), .B(KEYINPUT109), .ZN(new_n1235));
  INV_X1    g810(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g811(.A(KEYINPUT125), .B1(new_n1231), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g812(.A(KEYINPUT125), .ZN(new_n1238));
  AOI211_X1 g813(.A(new_n1238), .B(new_n1235), .C1(new_n1149), .C2(new_n1230), .ZN(new_n1239));
  OAI21_X1  g814(.A(new_n1031), .B1(new_n1237), .B2(new_n1239), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1242));
  NAND3_X1  g816(.A1(new_n673), .A2(G319), .A3(new_n674), .ZN(new_n1243));
  AOI21_X1  g817(.A(new_n1243), .B1(new_n655), .B2(new_n656), .ZN(new_n1244));
  NAND2_X1  g818(.A1(new_n702), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g819(.A(KEYINPUT126), .ZN(new_n1246));
  NAND2_X1  g820(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g821(.A1(new_n702), .A2(KEYINPUT126), .A3(new_n1244), .ZN(new_n1248));
  AOI22_X1  g822(.A1(new_n1247), .A2(new_n1248), .B1(new_n918), .B2(new_n920), .ZN(new_n1249));
  AND3_X1   g823(.A1(new_n991), .A2(new_n1242), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g824(.A(new_n1242), .B1(new_n991), .B2(new_n1249), .ZN(new_n1251));
  NOR2_X1   g825(.A1(new_n1250), .A2(new_n1251), .ZN(G308));
  NAND2_X1  g826(.A1(new_n991), .A2(new_n1249), .ZN(new_n1253));
  NAND2_X1  g827(.A1(new_n1253), .A2(KEYINPUT127), .ZN(new_n1254));
  NAND3_X1  g828(.A1(new_n991), .A2(new_n1249), .A3(new_n1242), .ZN(new_n1255));
  NAND2_X1  g829(.A1(new_n1254), .A2(new_n1255), .ZN(G225));
endmodule


