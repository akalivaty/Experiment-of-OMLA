//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n563, new_n564, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G101), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n467), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  XNOR2_X1  g057(.A(new_n470), .B(KEYINPUT69), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT70), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n483), .A2(new_n473), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n489), .B1(new_n491), .B2(G136), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n466), .A2(new_n469), .A3(new_n467), .A4(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n473), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n473), .A2(G138), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n470), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(new_n467), .A3(new_n476), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(G164));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT71), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n507), .A2(new_n508), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(G543), .B1(new_n506), .B2(new_n505), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(G651), .B1(new_n524), .B2(G50), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n518), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n514), .A2(G51), .A3(G543), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n510), .A2(G89), .A3(new_n516), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND2_X1  g110(.A1(new_n517), .A2(G90), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n520), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n524), .A2(G52), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n536), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n546), .B1(new_n511), .B2(new_n512), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g125(.A(KEYINPUT72), .B(new_n548), .C1(new_n520), .C2(new_n546), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n550), .A2(G651), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n524), .A2(G43), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n510), .A2(G81), .A3(new_n516), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT73), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n552), .A2(new_n554), .A3(new_n557), .A4(new_n553), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  OAI21_X1  g140(.A(G65), .B1(new_n507), .B2(new_n508), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT75), .B1(new_n568), .B2(G651), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  INV_X1    g145(.A(G651), .ZN(new_n571));
  AOI211_X1 g146(.A(new_n570), .B(new_n571), .C1(new_n566), .C2(new_n567), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n510), .A2(G91), .A3(new_n516), .ZN(new_n574));
  NAND2_X1  g149(.A1(KEYINPUT74), .A2(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n523), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  INV_X1    g152(.A(new_n575), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n514), .A2(new_n577), .A3(G543), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n573), .A2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G74), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n571), .B1(new_n520), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(G49), .B2(new_n524), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n510), .A2(G87), .A3(new_n516), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n517), .A2(G86), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n520), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(new_n524), .B2(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G305));
  NAND3_X1  g168(.A1(new_n510), .A2(G85), .A3(new_n516), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n524), .A2(G47), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n594), .A2(KEYINPUT78), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(KEYINPUT78), .B1(new_n594), .B2(new_n595), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n598));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n520), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n571), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g178(.A(KEYINPUT76), .B(new_n599), .C1(new_n520), .C2(new_n600), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n598), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n600), .B1(new_n511), .B2(new_n512), .ZN(new_n606));
  INV_X1    g181(.A(new_n599), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AND4_X1   g183(.A1(new_n598), .A2(new_n608), .A3(G651), .A4(new_n604), .ZN(new_n609));
  OAI22_X1  g184(.A1(new_n596), .A2(new_n597), .B1(new_n605), .B2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT79), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n510), .A2(G92), .A3(new_n516), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n510), .A2(KEYINPUT10), .A3(G92), .A4(new_n516), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n524), .A2(G54), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT80), .B(G66), .Z(new_n619));
  AOI22_X1  g194(.A1(new_n619), .A2(new_n513), .B1(G79), .B2(G543), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n620), .B2(new_n571), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT81), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n612), .B1(new_n624), .B2(G868), .ZN(G321));
  XOR2_X1   g200(.A(G321), .B(KEYINPUT82), .Z(G284));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n573), .A2(new_n581), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G280));
  XOR2_X1   g204(.A(G280), .B(KEYINPUT83), .Z(G297));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n559), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n621), .B1(new_n615), .B2(new_n616), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT81), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n636), .A2(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n634), .B1(new_n637), .B2(new_n633), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n491), .A2(G135), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n484), .A2(G123), .ZN(new_n641));
  OR2_X1    g216(.A1(G99), .A2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n642), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT85), .B(G2096), .Z(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n465), .A2(new_n468), .A3(G2105), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n647), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2100), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n644), .A2(new_n645), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n646), .A2(new_n651), .A3(new_n652), .ZN(G156));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n657), .B(new_n663), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(G14), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n667), .B2(new_n665), .ZN(G401));
  XOR2_X1   g244(.A(G2067), .B(G2678), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT86), .ZN(new_n671));
  NOR2_X1   g246(.A1(G2072), .A2(G2078), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n443), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT18), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n671), .A2(new_n673), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n673), .B(KEYINPUT17), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n678), .B(new_n675), .C1(new_n671), .C2(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n671), .A2(new_n679), .A3(new_n674), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2096), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n690), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n692), .B(new_n694), .C1(new_n687), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(G229));
  XNOR2_X1  g277(.A(KEYINPUT32), .B(G1981), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n588), .A2(G16), .A3(new_n592), .ZN(new_n705));
  OR2_X1    g280(.A1(G6), .A2(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(KEYINPUT88), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(KEYINPUT88), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n710), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n712), .A2(new_n703), .A3(new_n708), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G16), .A2(G23), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT89), .Z(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(G288), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT33), .B(G1976), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(G22), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT90), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G303), .B2(G16), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G1971), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n720), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n723), .B(KEYINPUT91), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G1971), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n714), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n730), .A2(KEYINPUT34), .B1(KEYINPUT93), .B2(KEYINPUT36), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT34), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n714), .A2(new_n727), .A3(new_n732), .A4(new_n729), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G25), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n473), .A2(G107), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n484), .A2(G119), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n491), .A2(G131), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n734), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT35), .B(G1991), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n743), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n745), .B(new_n735), .C1(new_n741), .C2(new_n734), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n717), .A2(G24), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G290), .B2(G16), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(G1986), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(G1986), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n744), .A2(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AND3_X1   g326(.A1(new_n733), .A2(KEYINPUT92), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(KEYINPUT92), .B1(new_n733), .B2(new_n751), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n731), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(KEYINPUT94), .ZN(new_n755));
  NOR2_X1   g330(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT94), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n757), .B(new_n731), .C1(new_n752), .C2(new_n753), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n734), .A2(G35), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n493), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT29), .ZN(new_n763));
  INV_X1    g338(.A(G2090), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT101), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n717), .A2(G4), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n624), .B2(new_n717), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1348), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n734), .A2(G26), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT28), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n491), .A2(G140), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n484), .A2(G128), .ZN(new_n774));
  OR2_X1    g349(.A1(G104), .A2(G2105), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n775), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n772), .B1(new_n777), .B2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G2067), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n717), .A2(G20), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT23), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  INV_X1    g358(.A(G1956), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OR3_X1    g360(.A1(new_n770), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n763), .A2(new_n764), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n717), .A2(G19), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n560), .B2(new_n717), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT95), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1341), .Z(new_n791));
  NOR3_X1   g366(.A1(new_n786), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT100), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT25), .ZN(new_n795));
  NAND2_X1  g370(.A1(G115), .A2(G2104), .ZN(new_n796));
  INV_X1    g371(.A(G127), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n477), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n795), .B1(G2105), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G139), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n490), .B2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g378(.A(KEYINPUT96), .B(new_n799), .C1(new_n490), .C2(new_n800), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n734), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n734), .B2(G33), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G2072), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n808), .A2(G28), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n734), .B1(new_n808), .B2(G28), .ZN(new_n810));
  AND2_X1   g385(.A1(KEYINPUT31), .A2(G11), .ZN(new_n811));
  NOR2_X1   g386(.A1(KEYINPUT31), .A2(G11), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n717), .A2(G21), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G168), .B2(new_n717), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n813), .B1(new_n815), .B2(G1966), .ZN(new_n816));
  INV_X1    g391(.A(G1961), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n717), .A2(G5), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G301), .B2(G16), .ZN(new_n819));
  OAI221_X1 g394(.A(new_n816), .B1(G1966), .B2(new_n815), .C1(new_n817), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n644), .A2(new_n734), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT99), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OR3_X1    g397(.A1(new_n820), .A2(KEYINPUT99), .A3(new_n821), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n807), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n734), .A2(G32), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n491), .A2(G141), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n484), .A2(G129), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT98), .B(KEYINPUT26), .ZN(new_n828));
  NAND3_X1  g403(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n473), .A2(G105), .A3(G2104), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT97), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n826), .A2(new_n827), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n825), .B1(new_n835), .B2(new_n734), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT27), .B(G1996), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT24), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(G34), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(G34), .ZN(new_n842));
  AOI21_X1  g417(.A(G29), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n481), .B2(G29), .ZN(new_n844));
  INV_X1    g419(.A(G2084), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n819), .A2(new_n817), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n734), .A2(G27), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G164), .B2(new_n734), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G2078), .ZN(new_n849));
  INV_X1    g424(.A(new_n844), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n849), .B1(G2084), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n838), .A2(new_n846), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n793), .B1(new_n824), .B2(new_n852), .ZN(new_n853));
  OR3_X1    g428(.A1(new_n824), .A2(new_n793), .A3(new_n852), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n767), .A2(new_n792), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n756), .B1(new_n755), .B2(new_n758), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n760), .A2(new_n855), .A3(new_n856), .ZN(G311));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n759), .ZN(G150));
  NAND2_X1  g434(.A1(G80), .A2(G543), .ZN(new_n860));
  INV_X1    g435(.A(G67), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n520), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G651), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n524), .A2(G55), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n510), .A2(new_n516), .ZN(new_n865));
  INV_X1    g440(.A(G93), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n863), .B(new_n864), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NOR2_X1   g444(.A1(new_n555), .A2(new_n867), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n559), .B2(new_n867), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT38), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n636), .A2(new_n631), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT102), .ZN(new_n877));
  AOI21_X1  g452(.A(G860), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n877), .A2(KEYINPUT103), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT103), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n869), .B1(new_n879), .B2(new_n880), .ZN(G145));
  XNOR2_X1  g456(.A(new_n493), .B(new_n481), .ZN(new_n882));
  INV_X1    g457(.A(new_n644), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n491), .A2(G142), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT106), .Z(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n888));
  INV_X1    g463(.A(G118), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(G2105), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n484), .B2(G130), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n739), .A2(new_n740), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(new_n649), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n893), .A2(new_n649), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n894), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n887), .A3(new_n891), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n501), .A2(new_n503), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n499), .A2(KEYINPUT104), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(new_n496), .B2(new_n498), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n900), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n803), .A2(KEYINPUT105), .A3(new_n804), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n835), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n834), .A2(KEYINPUT105), .A3(new_n803), .A4(new_n804), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n777), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n777), .B1(new_n906), .B2(new_n907), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n910), .ZN(new_n912));
  INV_X1    g487(.A(new_n904), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n913), .A3(new_n908), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n899), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n911), .A3(new_n899), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT107), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(KEYINPUT107), .B2(new_n916), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n885), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n884), .A2(new_n916), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(new_n915), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT40), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n915), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n916), .A2(KEYINPUT107), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n884), .B1(new_n928), .B2(new_n917), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT40), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n929), .A2(new_n923), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n925), .A2(new_n931), .ZN(G395));
  INV_X1    g507(.A(new_n867), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n556), .B2(new_n558), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n637), .B1(new_n934), .B2(new_n870), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n871), .B1(new_n636), .B2(G559), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n635), .A2(new_n628), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n635), .A2(new_n628), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT41), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n938), .B2(new_n939), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n623), .A2(G299), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n635), .A2(new_n628), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(KEYINPUT41), .A3(new_n945), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n935), .A2(new_n936), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT42), .B1(new_n941), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n935), .B(new_n936), .C1(new_n939), .C2(new_n938), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(G290), .A2(G288), .ZN(new_n953));
  INV_X1    g528(.A(G288), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n594), .A2(new_n595), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT78), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n594), .A2(KEYINPUT78), .A3(new_n595), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n608), .A2(G651), .A3(new_n604), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT77), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n603), .A2(new_n598), .A3(new_n604), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n954), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT108), .B1(new_n953), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(G290), .A2(G288), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n959), .A2(new_n954), .A3(new_n963), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(G303), .B(G305), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n965), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n970), .A2(new_n968), .A3(new_n966), .A4(new_n967), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n948), .A2(new_n952), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n948), .B2(new_n952), .ZN(new_n976));
  OAI21_X1  g551(.A(G868), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n867), .A2(new_n633), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(G295));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n977), .A2(new_n980), .A3(new_n978), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n977), .B2(new_n978), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(G331));
  INV_X1    g558(.A(G90), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n865), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n540), .A2(new_n541), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n533), .B(new_n532), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n536), .A2(G286), .A3(new_n542), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n559), .A2(new_n867), .ZN(new_n990));
  INV_X1    g565(.A(new_n870), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n987), .A2(new_n988), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n934), .A2(new_n993), .A3(new_n870), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n940), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n990), .A2(new_n991), .A3(new_n989), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n993), .B1(new_n934), .B2(new_n870), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n943), .A3(new_n997), .A4(new_n946), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n995), .A2(new_n972), .A3(new_n998), .A4(new_n973), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n999), .A2(new_n921), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(new_n998), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n974), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n995), .A2(new_n998), .A3(KEYINPUT111), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n974), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n1000), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1004), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n1011));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1000), .A2(new_n1012), .A3(new_n1002), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1012), .B1(new_n1008), .B2(new_n1000), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n999), .A2(new_n921), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1001), .A2(new_n1005), .B1(new_n973), .B2(new_n972), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n1007), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1019), .A2(KEYINPUT112), .A3(new_n1012), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT113), .B(new_n1011), .C1(new_n1016), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT112), .B1(new_n1019), .B2(new_n1012), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1009), .A2(new_n1015), .A3(KEYINPUT43), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n1013), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT113), .B1(new_n1025), .B2(new_n1011), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1010), .B1(new_n1022), .B2(new_n1026), .ZN(G397));
  INV_X1    g602(.A(new_n777), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n779), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n777), .A2(G2067), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(KEYINPUT115), .A3(new_n1030), .ZN(new_n1034));
  XOR2_X1   g609(.A(new_n834), .B(G1996), .Z(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT114), .B(G1384), .Z(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT45), .B1(new_n904), .B2(new_n1038), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n474), .A2(G40), .A3(new_n480), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT116), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1036), .A2(new_n1045), .A3(new_n1042), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n741), .A2(new_n743), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n893), .A2(new_n745), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1042), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1044), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(G290), .B(G1986), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1042), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1384), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n501), .A2(new_n503), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n499), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT50), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n904), .A2(new_n1057), .A3(new_n1053), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1040), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(G2084), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n904), .A2(new_n1053), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT45), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(KEYINPUT119), .A3(new_n1040), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G164), .A2(G1384), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(KEYINPUT120), .A3(KEYINPUT45), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT45), .B1(new_n904), .B2(new_n1053), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1040), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1064), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1966), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1060), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g653(.A(KEYINPUT123), .B(new_n1060), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(G286), .A2(G8), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n1084));
  INV_X1    g659(.A(G8), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n1080), .B2(G168), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1060), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1089), .B1(new_n1092), .B2(G8), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1082), .B(new_n1083), .C1(new_n1088), .C2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(KEYINPUT123), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(G168), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1093), .B1(new_n1097), .B2(new_n1086), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT62), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n1102));
  NAND2_X1  g677(.A1(G303), .A2(G8), .ZN(new_n1103));
  MUX2_X1   g678(.A(new_n1101), .B(new_n1102), .S(new_n1103), .Z(new_n1104));
  OAI21_X1  g679(.A(new_n1040), .B1(new_n1055), .B2(KEYINPUT50), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1057), .B1(new_n904), .B2(new_n1053), .ZN(new_n1106));
  OR3_X1    g681(.A1(new_n1105), .A2(G2090), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1055), .A2(new_n1062), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n904), .A2(KEYINPUT45), .A3(new_n1038), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n1040), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n726), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(KEYINPUT118), .B(new_n1104), .C1(new_n1112), .C2(new_n1085), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1040), .A2(new_n1053), .A3(new_n904), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1114), .A2(G8), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n954), .A2(G1976), .ZN(new_n1116));
  INV_X1    g691(.A(G1976), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT52), .B1(G288), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT49), .ZN(new_n1120));
  INV_X1    g695(.A(G1981), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n588), .A2(new_n1121), .A3(new_n592), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n588), .B2(new_n592), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(G305), .A2(G1981), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n588), .A2(new_n1121), .A3(new_n592), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(KEYINPUT49), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1115), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1114), .A2(new_n1116), .A3(G8), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT52), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1119), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1104), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1056), .A2(new_n1058), .A3(new_n764), .A4(new_n1040), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1085), .B1(new_n1111), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1131), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT118), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1085), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(new_n1132), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1113), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1109), .A2(new_n1040), .ZN(new_n1140));
  INV_X1    g715(.A(G2078), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n1141), .A3(new_n1108), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT124), .B(G1961), .Z(new_n1144));
  AOI22_X1  g719(.A1(new_n1142), .A2(new_n1143), .B1(new_n1059), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1143), .A2(G2078), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1064), .A2(new_n1069), .A3(new_n1073), .A4(new_n1146), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1139), .A2(G301), .A3(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1094), .A2(new_n1100), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1151));
  NOR2_X1   g726(.A1(G288), .A2(G1976), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1122), .B1(new_n1128), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1115), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1151), .A2(new_n1131), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1076), .A2(new_n1085), .A3(G286), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1111), .A2(new_n1133), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(G8), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1157), .B1(new_n1159), .B2(new_n1104), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1156), .A2(new_n1135), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT121), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1156), .A2(new_n1135), .A3(new_n1163), .A4(new_n1160), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1156), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1157), .B1(new_n1139), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1155), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n628), .B(KEYINPUT57), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT56), .B(G2072), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1140), .A2(new_n1108), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n784), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1114), .A2(G2067), .ZN(new_n1174));
  INV_X1    g749(.A(G1348), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n1175), .B2(new_n1059), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1176), .A2(new_n636), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1171), .A2(new_n1169), .A3(new_n1172), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1173), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT60), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n636), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(new_n1176), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n624), .A2(KEYINPUT60), .ZN(new_n1183));
  XOR2_X1   g758(.A(KEYINPUT58), .B(G1341), .Z(new_n1184));
  NAND2_X1  g759(.A1(new_n1114), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT122), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT122), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1114), .A2(new_n1187), .A3(new_n1184), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1186), .B(new_n1188), .C1(G1996), .C2(new_n1110), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT59), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1189), .A2(new_n1190), .A3(new_n560), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1190), .B1(new_n1189), .B2(new_n560), .ZN(new_n1192));
  OAI22_X1  g767(.A1(new_n1182), .A2(new_n1183), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1178), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1194), .B1(new_n1195), .B2(new_n1173), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1173), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1197), .A2(KEYINPUT61), .A3(new_n1178), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1179), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(G301), .B(KEYINPUT54), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1039), .A2(new_n1143), .A3(G2078), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(new_n1140), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1201), .B1(new_n1145), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1204), .B1(new_n1148), .B2(new_n1201), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1139), .A2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g781(.A(new_n1200), .B(new_n1206), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1168), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1052), .B1(new_n1150), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1050), .A2(KEYINPUT126), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1044), .A2(new_n1211), .A3(new_n1046), .A4(new_n1049), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1041), .A2(G1986), .A3(G290), .ZN(new_n1213));
  XNOR2_X1  g788(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n1213), .B(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1210), .A2(new_n1212), .A3(new_n1215), .ZN(new_n1216));
  AND3_X1   g791(.A1(new_n1044), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1029), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1042), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1041), .A2(G1996), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1220), .B(KEYINPUT46), .Z(new_n1221));
  NAND3_X1  g796(.A1(new_n1033), .A2(new_n835), .A3(new_n1034), .ZN(new_n1222));
  AND3_X1   g797(.A1(new_n1222), .A2(KEYINPUT125), .A3(new_n1042), .ZN(new_n1223));
  AOI21_X1  g798(.A(KEYINPUT125), .B1(new_n1222), .B2(new_n1042), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1221), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1225), .A2(KEYINPUT47), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT47), .ZN(new_n1227));
  OAI211_X1 g802(.A(new_n1227), .B(new_n1221), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  AND3_X1   g804(.A1(new_n1216), .A2(new_n1219), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1209), .A2(new_n1230), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g806(.A1(new_n920), .A2(new_n924), .ZN(new_n1233));
  NOR4_X1   g807(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1234));
  AND3_X1   g808(.A1(new_n1233), .A2(new_n1025), .A3(new_n1234), .ZN(G308));
  NAND3_X1  g809(.A1(new_n1233), .A2(new_n1025), .A3(new_n1234), .ZN(G225));
endmodule


