//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953;
  INV_X1    g000(.A(G148gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G141gat), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G155gat), .B(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(G155gat), .ZN(new_n208));
  INV_X1    g007(.A(G162gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT2), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AND4_X1   g009(.A1(KEYINPUT73), .A2(new_n206), .A3(new_n207), .A4(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT73), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(new_n203), .B2(new_n205), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n207), .B1(new_n213), .B2(new_n210), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(G127gat), .B(G134gat), .Z(new_n216));
  XNOR2_X1  g015(.A(G113gat), .B(G120gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(KEYINPUT1), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G113gat), .B(G120gat), .Z(new_n219));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n206), .A2(KEYINPUT73), .A3(new_n210), .ZN(new_n224));
  INV_X1    g023(.A(new_n207), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n213), .A2(new_n207), .A3(new_n210), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n215), .A2(new_n223), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G225gat), .A2(G233gat), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n226), .A2(new_n228), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT4), .B1(new_n235), .B2(new_n223), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT74), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(new_n211), .B2(new_n214), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n226), .A2(KEYINPUT74), .A3(new_n228), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n223), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n237), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT78), .B1(new_n234), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n238), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n236), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT78), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n232), .A4(new_n233), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G1gat), .B(G29gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT0), .ZN(new_n251));
  XNOR2_X1  g050(.A(G57gat), .B(G85gat), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n251), .B(new_n252), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n242), .A2(KEYINPUT4), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n238), .B1(new_n235), .B2(new_n223), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n232), .A2(KEYINPUT75), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT75), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n230), .A2(new_n231), .A3(new_n255), .ZN(new_n258));
  AOI211_X1 g057(.A(new_n238), .B(new_n223), .C1(new_n240), .C2(new_n241), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n231), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n211), .A2(new_n214), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n218), .A2(new_n222), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n235), .A2(new_n223), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n233), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT77), .B1(new_n261), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT77), .ZN(new_n272));
  AOI211_X1 g071(.A(new_n272), .B(new_n269), .C1(new_n256), .C2(new_n260), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n249), .B(new_n253), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n253), .B(KEYINPUT81), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n230), .A2(new_n231), .A3(new_n255), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT75), .B1(new_n278), .B2(new_n254), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n258), .A2(new_n259), .A3(new_n257), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n270), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n272), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n261), .A2(KEYINPUT77), .A3(new_n270), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n277), .B1(new_n284), .B2(new_n249), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT84), .B1(new_n276), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n249), .B1(new_n271), .B2(new_n273), .ZN(new_n287));
  INV_X1    g086(.A(new_n277), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT84), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n289), .A2(new_n290), .A3(new_n275), .A4(new_n274), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n253), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n287), .A2(KEYINPUT6), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT79), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n287), .A2(KEYINPUT79), .A3(KEYINPUT6), .A4(new_n293), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G8gat), .B(G36gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT72), .ZN(new_n300));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT23), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308));
  INV_X1    g107(.A(G169gat), .ZN(new_n309));
  INV_X1    g108(.A(G176gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n307), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT64), .ZN(new_n315));
  OAI221_X1 g114(.A(new_n313), .B1(G183gat), .B2(G190gat), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n314), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(KEYINPUT64), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n305), .B(new_n312), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT25), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n311), .A2(new_n308), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n305), .A3(new_n306), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(new_n320), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n317), .B(new_n313), .C1(G183gat), .C2(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n307), .A2(new_n304), .A3(KEYINPUT26), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT26), .ZN(new_n329));
  INV_X1    g128(.A(G183gat), .ZN(new_n330));
  INV_X1    g129(.A(G190gat), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n311), .A2(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(KEYINPUT27), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT27), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G183gat), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(KEYINPUT28), .A3(new_n331), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(new_n336), .A3(new_n331), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(KEYINPUT66), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT66), .B1(new_n339), .B2(new_n340), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n333), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n348));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G211gat), .B(G218gat), .ZN(new_n351));
  INV_X1    g150(.A(G211gat), .ZN(new_n352));
  INV_X1    g151(.A(G218gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT69), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT69), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G218gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT70), .B1(new_n357), .B2(KEYINPUT22), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT70), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT22), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT69), .B(G218gat), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n359), .B(new_n360), .C1(new_n361), .C2(new_n352), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(G197gat), .B(G204gat), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n351), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n351), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n364), .B(new_n367), .C1(new_n358), .C2(new_n362), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n319), .A2(new_n320), .B1(new_n324), .B2(new_n325), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT67), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n344), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(KEYINPUT67), .B(new_n333), .C1(new_n342), .C2(new_n343), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(new_n349), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT29), .B1(new_n327), .B2(new_n344), .ZN(new_n377));
  INV_X1    g176(.A(new_n349), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT71), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n350), .B(new_n370), .C1(new_n376), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n349), .A2(new_n346), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n375), .A2(new_n381), .B1(new_n349), .B2(new_n345), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n369), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n385));
  AOI21_X1  g184(.A(new_n303), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT38), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n376), .A2(new_n379), .ZN(new_n388));
  INV_X1    g187(.A(new_n350), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n369), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n382), .A2(new_n369), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(KEYINPUT37), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(new_n387), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n302), .B1(new_n380), .B2(new_n383), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n380), .A2(new_n383), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT37), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n387), .B1(new_n398), .B2(new_n386), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n292), .A2(new_n298), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G78gat), .B(G106gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(G22gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n229), .A2(new_n346), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n369), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n346), .B1(new_n366), .B2(new_n368), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n408), .A2(new_n227), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n240), .A2(new_n241), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n405), .B(new_n407), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT31), .B(G50gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n407), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n408), .A2(KEYINPUT80), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT80), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n416), .B(new_n346), .C1(new_n366), .C2(new_n368), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n227), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n418), .B2(new_n235), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n411), .B(new_n413), .C1(new_n419), .C2(new_n405), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT3), .B1(new_n408), .B2(KEYINPUT80), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n263), .B1(new_n422), .B2(new_n417), .ZN(new_n423));
  OAI211_X1 g222(.A(G228gat), .B(G233gat), .C1(new_n423), .C2(new_n414), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n413), .B1(new_n424), .B2(new_n411), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n404), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n411), .B1(new_n419), .B2(new_n405), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n412), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n403), .A3(new_n420), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT39), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n246), .A2(new_n230), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT82), .B1(new_n432), .B2(new_n262), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n434));
  AOI211_X1 g233(.A(new_n434), .B(new_n231), .C1(new_n246), .C2(new_n230), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n431), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n230), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n262), .B1(new_n243), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n434), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n432), .A2(KEYINPUT82), .A3(new_n262), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n265), .A2(new_n266), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n431), .B1(new_n441), .B2(new_n231), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n436), .A2(new_n443), .A3(new_n277), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT40), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(KEYINPUT83), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(KEYINPUT83), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n436), .A2(new_n443), .A3(new_n277), .A4(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n446), .A2(new_n289), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n380), .A2(new_n383), .A3(new_n302), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT30), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(new_n394), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n397), .A2(KEYINPUT30), .A3(new_n302), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n430), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n401), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(G227gat), .ZN(new_n457));
  INV_X1    g256(.A(G233gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n375), .A2(new_n264), .ZN(new_n460));
  AOI211_X1 g259(.A(new_n223), .B(new_n371), .C1(new_n373), .C2(new_n374), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G71gat), .B(G99gat), .Z(new_n463));
  XNOR2_X1  g262(.A(G15gat), .B(G43gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(KEYINPUT33), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n462), .A2(KEYINPUT32), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n459), .ZN(new_n470));
  INV_X1    g269(.A(new_n343), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n338), .A3(new_n341), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT67), .B1(new_n472), .B2(new_n333), .ZN(new_n473));
  INV_X1    g272(.A(new_n374), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n327), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n223), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n375), .A2(new_n264), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n470), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT32), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n465), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n478), .A2(KEYINPUT33), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n469), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n476), .A2(new_n477), .A3(new_n470), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT34), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n462), .A2(KEYINPUT32), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT33), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n462), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n488), .A3(new_n465), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT34), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n483), .B(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n491), .A3(new_n469), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n485), .A2(new_n492), .A3(KEYINPUT36), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT36), .B1(new_n485), .B2(new_n492), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n287), .A2(new_n293), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(new_n275), .A3(new_n274), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n296), .A2(new_n497), .A3(new_n297), .ZN(new_n498));
  INV_X1    g297(.A(new_n454), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n495), .B1(new_n500), .B2(new_n430), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n426), .A2(new_n429), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n492), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n498), .A2(new_n502), .A3(new_n499), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n292), .A2(new_n298), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(new_n452), .B2(new_n453), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n430), .A2(new_n509), .A3(new_n503), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n456), .A2(new_n501), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(G29gat), .A2(G36gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G29gat), .A2(G36gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT88), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n515), .A2(KEYINPUT15), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n518), .A2(new_n520), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT15), .B1(new_n515), .B2(new_n517), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT17), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT89), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(KEYINPUT89), .A3(G1gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G8gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n525), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n524), .A2(new_n534), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n536), .A2(KEYINPUT18), .A3(new_n537), .A4(new_n538), .ZN(new_n542));
  OR3_X1    g341(.A1(new_n524), .A2(new_n534), .A3(KEYINPUT90), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT90), .B1(new_n524), .B2(new_n534), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n537), .B(KEYINPUT13), .Z(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n541), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT87), .B(G197gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT11), .B(G169gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT12), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n541), .A2(new_n542), .A3(new_n547), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n298), .A2(KEYINPUT103), .A3(new_n497), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT103), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n498), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n512), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT21), .ZN(new_n565));
  INV_X1    g364(.A(G57gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(G64gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT92), .ZN(new_n568));
  NAND2_X1  g367(.A1(KEYINPUT92), .A2(G57gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(KEYINPUT91), .A3(G64gat), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n566), .A2(G64gat), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n568), .B(new_n570), .C1(KEYINPUT91), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  OR2_X1    g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT9), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT9), .B1(new_n571), .B2(new_n567), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(new_n573), .A3(new_n574), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n535), .B1(new_n565), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT94), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G155gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n582), .B(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(G127gat), .ZN(new_n590));
  XOR2_X1   g389(.A(G183gat), .B(G211gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n585), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT7), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(new_n598), .B2(new_n599), .ZN(new_n602));
  NAND3_X1  g401(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  OR2_X1    g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT96), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n525), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT97), .ZN(new_n612));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT95), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT41), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n608), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n524), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n611), .A2(KEYINPUT97), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n614), .A2(new_n615), .ZN(new_n624));
  XOR2_X1   g423(.A(G134gat), .B(G162gat), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n626), .A3(new_n622), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n596), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n608), .A2(new_n580), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT10), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n606), .A2(new_n577), .A3(new_n579), .A4(new_n607), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT98), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n633), .A2(new_n638), .A3(new_n634), .A4(new_n635), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640));
  OR3_X1    g439(.A1(new_n635), .A2(new_n640), .A3(new_n634), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n640), .B1(new_n635), .B2(new_n634), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n637), .A2(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n633), .A2(new_n635), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n645), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  NOR2_X1   g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n656), .B1(new_n655), .B2(new_n648), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n644), .B1(new_n643), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n637), .A2(new_n639), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n641), .A2(new_n642), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n660), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n657), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g464(.A(KEYINPUT102), .B(new_n657), .C1(new_n659), .C2(new_n662), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n654), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n632), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n564), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g470(.A1(new_n512), .A2(new_n668), .A3(new_n559), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n454), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT104), .Z(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(G8gat), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT16), .B(G8gat), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n677));
  INV_X1    g476(.A(new_n676), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  OAI221_X1 g478(.A(new_n675), .B1(new_n673), .B2(new_n677), .C1(new_n679), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g479(.A(new_n672), .ZN(new_n681));
  INV_X1    g480(.A(new_n495), .ZN(new_n682));
  OAI21_X1  g481(.A(G15gat), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n503), .A2(G15gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n681), .B2(new_n684), .ZN(G1326gat));
  NAND2_X1  g484(.A1(new_n672), .A2(new_n430), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  INV_X1    g487(.A(G29gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n660), .A2(new_n661), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT100), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n643), .A2(new_n658), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n692), .A3(new_n644), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT102), .B1(new_n693), .B2(new_n657), .ZN(new_n694));
  INV_X1    g493(.A(new_n666), .ZN(new_n695));
  OAI22_X1  g494(.A1(new_n694), .A2(new_n695), .B1(new_n653), .B2(new_n650), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n595), .A2(new_n630), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n564), .A2(new_n689), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n512), .B2(new_n630), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n456), .A2(new_n501), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n506), .A2(new_n511), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(KEYINPUT44), .A3(new_n631), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n559), .A2(new_n595), .A3(new_n696), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n701), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n563), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n699), .A2(new_n708), .ZN(G1328gat));
  AND3_X1   g508(.A1(new_n704), .A2(new_n558), .A3(new_n697), .ZN(new_n710));
  AOI21_X1  g509(.A(G36gat), .B1(KEYINPUT105), .B2(KEYINPUT46), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n454), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G36gat), .B1(new_n707), .B2(new_n499), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1329gat));
  OAI21_X1  g515(.A(G43gat), .B1(new_n707), .B2(new_n682), .ZN(new_n717));
  INV_X1    g516(.A(G43gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n710), .A2(new_n718), .A3(new_n504), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g520(.A(G50gat), .B1(new_n707), .B2(new_n502), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n502), .A2(G50gat), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT106), .Z(new_n724));
  NAND2_X1  g523(.A1(new_n710), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT48), .Z(G1331gat));
  NAND4_X1  g526(.A1(new_n704), .A2(new_n632), .A3(new_n696), .A4(new_n559), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n563), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT107), .B(G57gat), .Z(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1332gat));
  NOR2_X1   g530(.A1(new_n728), .A2(new_n499), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT49), .B(G64gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT108), .ZN(G1333gat));
  OR3_X1    g536(.A1(new_n728), .A2(G71gat), .A3(new_n503), .ZN(new_n738));
  OAI21_X1  g537(.A(G71gat), .B1(new_n728), .B2(new_n682), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g540(.A1(new_n728), .A2(new_n502), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT109), .B(G78gat), .Z(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1335gat));
  NOR2_X1   g543(.A1(new_n595), .A2(new_n558), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n704), .A2(KEYINPUT51), .A3(new_n631), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT111), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n745), .ZN(new_n749));
  AOI211_X1 g548(.A(new_n630), .B(new_n749), .C1(new_n702), .C2(new_n703), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(KEYINPUT51), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n563), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(new_n598), .A3(new_n696), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n749), .A2(new_n667), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n701), .A2(new_n705), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT110), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n701), .A2(new_n705), .A3(new_n758), .A4(new_n755), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n757), .A2(new_n753), .A3(new_n759), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n752), .A2(new_n754), .B1(new_n760), .B2(new_n598), .ZN(G1336gat));
  NOR3_X1   g560(.A1(new_n499), .A2(new_n667), .A3(G92gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n751), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764));
  OAI21_X1  g563(.A(G92gat), .B1(new_n756), .B2(new_n499), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n757), .A2(new_n454), .A3(new_n759), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G92gat), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT112), .B1(new_n750), .B2(KEYINPUT51), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n704), .A2(new_n631), .A3(new_n745), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n762), .B1(new_n747), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n768), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT113), .B1(new_n776), .B2(KEYINPUT52), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n778), .B(new_n764), .C1(new_n768), .C2(new_n775), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n766), .B1(new_n777), .B2(new_n779), .ZN(G1337gat));
  INV_X1    g579(.A(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n504), .A2(new_n696), .A3(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n757), .A2(new_n495), .A3(new_n759), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n752), .A2(new_n782), .B1(new_n783), .B2(new_n781), .ZN(G1338gat));
  OAI21_X1  g583(.A(G106gat), .B1(new_n756), .B2(new_n502), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  OR3_X1    g585(.A1(new_n502), .A2(G106gat), .A3(new_n667), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n785), .B(new_n786), .C1(new_n752), .C2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n757), .A2(new_n430), .A3(new_n759), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n789), .A2(new_n790), .A3(G106gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n789), .B2(G106gat), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n769), .A2(new_n773), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n787), .B1(new_n748), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n788), .B1(new_n795), .B2(new_n786), .ZN(G1339gat));
  AOI21_X1  g595(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n545), .A2(new_n546), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n553), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n557), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(new_n696), .A3(KEYINPUT117), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n557), .A2(new_n799), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(new_n667), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n643), .A2(new_n645), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT54), .B(new_n806), .C1(new_n659), .C2(new_n662), .ZN(new_n807));
  XOR2_X1   g606(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n808));
  AOI21_X1  g607(.A(new_n653), .B1(new_n646), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(KEYINPUT55), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n694), .B2(new_n695), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n810), .B(new_n813), .C1(new_n694), .C2(new_n695), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n807), .A2(new_n809), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n812), .A2(new_n558), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n631), .B1(new_n805), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n630), .A2(new_n803), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n820), .A2(new_n814), .A3(new_n812), .A4(new_n817), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n596), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n668), .A2(new_n558), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n430), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  AND4_X1   g625(.A1(new_n499), .A2(new_n826), .A3(new_n504), .A4(new_n753), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n558), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n696), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n595), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g632(.A1(new_n827), .A2(new_n631), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n834), .A2(G134gat), .B1(new_n835), .B2(KEYINPUT56), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(KEYINPUT119), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n835), .B(KEYINPUT56), .C1(new_n834), .C2(G134gat), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n834), .A2(G134gat), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(KEYINPUT118), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(KEYINPUT118), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n838), .B(new_n839), .C1(new_n841), .C2(new_n842), .ZN(G1343gat));
  AOI21_X1  g642(.A(new_n502), .B1(new_n823), .B2(new_n825), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n563), .A2(new_n495), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR4_X1   g645(.A1(new_n846), .A2(G141gat), .A3(new_n454), .A4(new_n559), .ZN(new_n847));
  XOR2_X1   g646(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n800), .A2(new_n696), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n558), .A2(new_n817), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n811), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n630), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n595), .B1(new_n854), .B2(new_n821), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n430), .B1(new_n855), .B2(new_n824), .ZN(new_n856));
  OAI22_X1  g655(.A1(new_n844), .A2(new_n849), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n845), .A2(new_n499), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT121), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n857), .A2(new_n862), .A3(new_n859), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n558), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n847), .B1(new_n864), .B2(G141gat), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n846), .A2(KEYINPUT122), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n846), .A2(KEYINPUT122), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n867), .A2(new_n868), .A3(new_n454), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n869), .A2(new_n204), .A3(new_n558), .ZN(new_n870));
  OAI21_X1  g669(.A(G141gat), .B1(new_n860), .B2(new_n559), .ZN(new_n871));
  XOR2_X1   g670(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI22_X1  g672(.A1(new_n865), .A2(new_n866), .B1(new_n870), .B2(new_n873), .ZN(G1344gat));
  INV_X1    g673(.A(new_n863), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n862), .B1(new_n857), .B2(new_n859), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n878), .A3(new_n696), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n818), .A2(new_n804), .A3(new_n801), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n630), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n595), .B1(new_n881), .B2(new_n821), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n430), .B(new_n849), .C1(new_n882), .C2(new_n824), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n856), .A2(new_n850), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n696), .A3(new_n859), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n202), .B1(new_n886), .B2(KEYINPUT59), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n696), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n878), .A2(G148gat), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n879), .A2(new_n887), .B1(new_n888), .B2(new_n889), .ZN(G1345gat));
  NAND3_X1  g689(.A1(new_n869), .A2(new_n208), .A3(new_n595), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n875), .A2(new_n596), .A3(new_n876), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n208), .ZN(G1346gat));
  AOI21_X1  g692(.A(G162gat), .B1(new_n869), .B2(new_n631), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n630), .A2(new_n209), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n877), .B2(new_n895), .ZN(G1347gat));
  NOR3_X1   g695(.A1(new_n753), .A2(new_n499), .A3(new_n503), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n826), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n826), .A2(KEYINPUT124), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(new_n309), .A3(new_n559), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n753), .B1(new_n823), .B2(new_n825), .ZN(new_n904));
  AND4_X1   g703(.A1(new_n502), .A2(new_n904), .A3(new_n454), .A4(new_n504), .ZN(new_n905));
  AOI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n558), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n903), .A2(new_n906), .ZN(G1348gat));
  OAI21_X1  g706(.A(G176gat), .B1(new_n902), .B2(new_n667), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n310), .A3(new_n696), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1349gat));
  OAI21_X1  g709(.A(G183gat), .B1(new_n902), .B2(new_n596), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n905), .A2(new_n595), .A3(new_n337), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT60), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n631), .A3(new_n901), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(G190gat), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n331), .A3(new_n631), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT125), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(G1351gat));
  NOR3_X1   g723(.A1(new_n753), .A2(new_n499), .A3(new_n495), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n926), .B1(new_n883), .B2(new_n884), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(G197gat), .A3(new_n558), .ZN(new_n928));
  AND4_X1   g727(.A1(new_n430), .A2(new_n904), .A3(new_n454), .A4(new_n682), .ZN(new_n929));
  AOI21_X1  g728(.A(G197gat), .B1(new_n929), .B2(new_n558), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n928), .A2(new_n930), .ZN(G1352gat));
  INV_X1    g730(.A(G204gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n929), .A2(new_n932), .A3(new_n696), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT62), .Z(new_n934));
  INV_X1    g733(.A(new_n927), .ZN(new_n935));
  OAI21_X1  g734(.A(G204gat), .B1(new_n935), .B2(new_n667), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1353gat));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n885), .A2(new_n939), .A3(new_n595), .A4(new_n925), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n927), .B2(new_n595), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n885), .A2(new_n595), .A3(new_n925), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n945), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n940), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n943), .A2(KEYINPUT127), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n948), .B(new_n938), .C1(new_n941), .C2(new_n942), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n929), .A2(new_n352), .A3(new_n595), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(G1354gat));
  AOI21_X1  g750(.A(G218gat), .B1(new_n929), .B2(new_n631), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n630), .A2(new_n361), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n927), .B2(new_n953), .ZN(G1355gat));
endmodule


