//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n558, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT67), .A4(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(new_n470), .B2(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NOR3_X1   g048(.A1(new_n473), .A2(new_n463), .A3(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(KEYINPUT69), .B1(new_n475), .B2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n465), .B1(new_n463), .B2(KEYINPUT68), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n477), .A2(G101), .B1(new_n481), .B2(G137), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n472), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  AOI21_X1  g059(.A(new_n475), .B1(new_n478), .B2(new_n480), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(new_n486), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  MUX2_X1   g065(.A(G100), .B(G112), .S(G2105), .Z(new_n491));
  AOI22_X1  g066(.A1(new_n481), .A2(G136), .B1(new_n491), .B2(G2104), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n490), .A2(new_n492), .ZN(G162));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n495), .A2(new_n464), .A3(new_n466), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT72), .B(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI211_X1 g073(.A(new_n494), .B(G2105), .C1(new_n478), .C2(new_n480), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT71), .A2(G114), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT71), .A2(G114), .ZN(new_n503));
  OAI21_X1  g078(.A(G2105), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n475), .A2(G102), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G2104), .B1(new_n485), .B2(G126), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT73), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XOR2_X1   g090(.A(new_n515), .B(KEYINPUT74), .Z(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n514), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n519), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n511), .B2(new_n513), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  OAI211_X1 g100(.A(G88), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  OAI211_X1 g101(.A(G50), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n521), .A2(new_n526), .A3(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NOR2_X1   g104(.A1(new_n524), .A2(new_n525), .ZN(new_n530));
  INV_X1    g105(.A(new_n522), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(G543), .B1(new_n524), .B2(new_n525), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n522), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n533), .A2(new_n536), .A3(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n532), .A2(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n535), .A2(G52), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n514), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(new_n532), .A2(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n535), .A2(G43), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n547), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  OAI211_X1 g137(.A(G53), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  OAI211_X1 g139(.A(G91), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n531), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n566), .A2(KEYINPUT75), .B1(G651), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n564), .A2(new_n570), .A3(new_n572), .ZN(G299));
  OAI21_X1  g148(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g151(.A(KEYINPUT76), .B(G651), .C1(new_n522), .C2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g153(.A(G87), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(new_n579));
  OAI211_X1 g154(.A(G49), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  OAI211_X1 g156(.A(G48), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n582));
  OAI211_X1 g157(.A(G86), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n518), .B2(new_n519), .ZN(new_n585));
  AND2_X1   g160(.A1(G73), .A2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n514), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n582), .A2(new_n583), .A3(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT77), .A4(new_n587), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n531), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n595), .A2(new_n596), .A3(new_n514), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT78), .B1(new_n598), .B2(new_n547), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g175(.A(G47), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n601));
  OAI211_X1 g176(.A(G85), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n600), .A2(new_n603), .ZN(G290));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(G301), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT79), .B(G66), .Z(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(new_n522), .B1(G79), .B2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G54), .ZN(new_n609));
  OAI22_X1  g184(.A1(new_n510), .A2(new_n608), .B1(new_n534), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g185(.A(G92), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n606), .B1(new_n605), .B2(new_n615), .ZN(G284));
  AOI21_X1  g191(.A(new_n606), .B1(new_n605), .B2(new_n615), .ZN(G321));
  NOR2_X1   g192(.A1(G286), .A2(new_n605), .ZN(new_n618));
  AND3_X1   g193(.A1(new_n564), .A2(new_n572), .A3(new_n570), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n605), .ZN(G297));
  AOI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(new_n605), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  NOR2_X1   g198(.A1(new_n555), .A2(G868), .ZN(new_n624));
  INV_X1    g199(.A(new_n615), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n625), .A2(G559), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n624), .B1(new_n626), .B2(G868), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n477), .A2(new_n470), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OAI22_X1  g207(.A1(new_n630), .A2(new_n631), .B1(KEYINPUT80), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(new_n631), .B2(new_n630), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G2100), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n634), .A2(KEYINPUT80), .A3(new_n632), .ZN(new_n638));
  MUX2_X1   g213(.A(G99), .B(G111), .S(G2105), .Z(new_n639));
  AOI22_X1  g214(.A1(new_n481), .A2(G135), .B1(new_n639), .B2(G2104), .ZN(new_n640));
  INV_X1    g215(.A(new_n489), .ZN(new_n641));
  INV_X1    g216(.A(G123), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n637), .A2(new_n638), .A3(new_n644), .ZN(G156));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT15), .B(G2435), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2427), .ZN(new_n649));
  INV_X1    g224(.A(G2430), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n649), .ZN(new_n652));
  XOR2_X1   g227(.A(G2443), .B(G2446), .Z(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT82), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n652), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2084), .B(G2090), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT83), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT84), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n666), .B(KEYINPUT17), .Z(new_n670));
  INV_X1    g245(.A(new_n667), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(KEYINPUT84), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n667), .A2(new_n664), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n671), .A2(new_n664), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n666), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT18), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G2096), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n682), .A2(G2100), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(G2100), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n687), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n687), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n699), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  NOR2_X1   g279(.A1(G4), .A2(G16), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT88), .Z(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n625), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1348), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(G32), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n481), .A2(G141), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n712), .B(new_n715), .C1(G105), .C2(new_n477), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n489), .A2(G129), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT92), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n711), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT27), .B(G1996), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n710), .A2(G35), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT96), .Z(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G162), .B2(new_n710), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT29), .Z(new_n728));
  INV_X1    g303(.A(G2090), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n709), .B(new_n724), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n722), .B2(new_n723), .ZN(new_n732));
  AND2_X1   g307(.A1(KEYINPUT24), .A2(G34), .ZN(new_n733));
  NOR2_X1   g308(.A1(KEYINPUT24), .A2(G34), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n710), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n483), .B2(new_n710), .ZN(new_n736));
  INV_X1    g311(.A(G2084), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(G164), .A2(G29), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G27), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT95), .B(G2078), .ZN(new_n741));
  NOR2_X1   g316(.A1(G168), .A2(new_n707), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n707), .B2(G21), .ZN(new_n743));
  INV_X1    g318(.A(G1966), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n738), .B1(new_n740), .B2(new_n741), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n743), .A2(new_n744), .B1(new_n737), .B2(new_n736), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n707), .A2(G5), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G171), .B2(new_n707), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n749), .A2(new_n750), .B1(new_n740), .B2(new_n741), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n730), .A2(new_n732), .A3(new_n745), .A4(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT25), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G139), .B2(new_n481), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT90), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(new_n475), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(new_n710), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n710), .B2(G33), .ZN(new_n763));
  INV_X1    g338(.A(G2072), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT91), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n707), .A2(G19), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT89), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n556), .B2(new_n707), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G1341), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n710), .A2(G26), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT28), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n489), .A2(G128), .ZN(new_n774));
  MUX2_X1   g349(.A(G104), .B(G116), .S(G2105), .Z(new_n775));
  AOI22_X1  g350(.A1(new_n481), .A2(G140), .B1(new_n775), .B2(G2104), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n773), .B1(new_n777), .B2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2067), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT31), .B(G11), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT94), .B(G28), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(KEYINPUT30), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(KEYINPUT30), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(new_n710), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n780), .B1(new_n782), .B2(new_n784), .C1(new_n643), .C2(new_n710), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G1961), .B2(new_n748), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n767), .A2(new_n771), .A3(new_n779), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n766), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n707), .A2(G20), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT23), .Z(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G299), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1956), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n753), .A2(new_n788), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n489), .A2(G119), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n481), .A2(G131), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT85), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G95), .B(G107), .S(G2105), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G2104), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n794), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT86), .Z(new_n801));
  MUX2_X1   g376(.A(G25), .B(new_n801), .S(G29), .Z(new_n802));
  XOR2_X1   g377(.A(KEYINPUT35), .B(G1991), .Z(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n802), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n707), .A2(G24), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT87), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G290), .B2(G16), .ZN(new_n808));
  INV_X1    g383(.A(G1986), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G6), .A2(G16), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n590), .A2(new_n591), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(G16), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT32), .B(G1981), .Z(new_n815));
  XOR2_X1   g390(.A(new_n814), .B(new_n815), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n707), .A2(G23), .ZN(new_n817));
  INV_X1    g392(.A(G288), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n707), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT33), .B(G1976), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(G16), .A2(G22), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G166), .B2(G16), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1971), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n816), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT34), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n811), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT36), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n811), .A2(new_n828), .A3(new_n831), .A4(new_n827), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n793), .B1(new_n830), .B2(new_n832), .ZN(G311));
  NAND2_X1  g408(.A1(new_n830), .A2(new_n832), .ZN(new_n834));
  INV_X1    g409(.A(new_n793), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(G150));
  NAND2_X1  g411(.A1(new_n532), .A2(G93), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n535), .A2(G55), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(new_n547), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  OR2_X1    g418(.A1(new_n555), .A2(new_n841), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n555), .A2(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n625), .A2(new_n622), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  INV_X1    g425(.A(G860), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n843), .B1(new_n850), .B2(new_n852), .ZN(G145));
  MUX2_X1   g428(.A(G106), .B(G118), .S(G2105), .Z(new_n854));
  AOI22_X1  g429(.A1(new_n481), .A2(G142), .B1(new_n854), .B2(G2104), .ZN(new_n855));
  INV_X1    g430(.A(G130), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n641), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n630), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n800), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n761), .B(new_n716), .C1(new_n720), .C2(new_n719), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n721), .A2(new_n760), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n777), .B(G164), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n860), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT98), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n860), .A2(new_n870), .A3(new_n866), .A4(new_n867), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n866), .A2(new_n867), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n859), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(G162), .B(new_n483), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n643), .B(KEYINPUT97), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(KEYINPUT99), .B(G37), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n868), .A2(new_n877), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(new_n873), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n879), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(G395));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n891));
  AND3_X1   g466(.A1(G299), .A2(new_n891), .A3(new_n615), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(G299), .B2(new_n615), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n619), .A2(new_n625), .A3(KEYINPUT102), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(G299), .B2(new_n615), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n890), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n846), .A2(new_n626), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n844), .B(new_n845), .C1(G559), .C2(new_n625), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  OAI221_X1 g479(.A(new_n904), .B1(G299), .B2(new_n615), .C1(new_n892), .C2(new_n893), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(G290), .A2(G288), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n535), .A2(G49), .B1(new_n576), .B2(new_n577), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n908), .A2(new_n600), .A3(new_n579), .A4(new_n603), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(G305), .A2(G166), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n813), .A2(G303), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n813), .A2(G303), .ZN(new_n914));
  AOI21_X1  g489(.A(G166), .B1(new_n590), .B2(new_n591), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n907), .B(new_n909), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n913), .A2(new_n916), .A3(KEYINPUT104), .A4(KEYINPUT42), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n913), .A2(new_n916), .ZN(new_n918));
  XNOR2_X1  g493(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(G299), .A2(new_n615), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n894), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n900), .A3(new_n901), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n906), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n920), .B1(new_n906), .B2(new_n923), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(KEYINPUT105), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n927));
  AOI211_X1 g502(.A(new_n927), .B(new_n920), .C1(new_n923), .C2(new_n906), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n841), .A2(new_n605), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n932));
  NAND2_X1  g507(.A1(G331), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(G295));
  NAND2_X1  g510(.A1(G168), .A2(G171), .ZN(new_n936));
  NAND2_X1  g511(.A1(G301), .A2(G286), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n844), .A2(new_n936), .A3(new_n845), .A4(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n844), .A2(new_n845), .B1(new_n936), .B2(new_n937), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT41), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n894), .A2(new_n898), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n936), .A2(new_n937), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n846), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n903), .B1(new_n944), .B2(new_n938), .ZN(new_n945));
  OAI22_X1  g520(.A1(new_n941), .A2(new_n942), .B1(new_n945), .B2(new_n922), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n881), .B1(new_n946), .B2(new_n918), .ZN(new_n947));
  INV_X1    g522(.A(new_n918), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n939), .A2(new_n940), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n894), .B2(new_n921), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n899), .A2(new_n905), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n948), .B(new_n950), .C1(new_n951), .C2(new_n949), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n950), .B1(new_n951), .B2(new_n949), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n918), .ZN(new_n957));
  INV_X1    g532(.A(G37), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n957), .A2(new_n952), .A3(KEYINPUT43), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT44), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n958), .A3(new_n952), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(KEYINPUT43), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n960), .B1(KEYINPUT44), .B2(new_n963), .ZN(G397));
  NOR2_X1   g539(.A1(G290), .A2(G1986), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n809), .B1(new_n600), .B2(new_n603), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n965), .A2(KEYINPUT107), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(G1384), .B1(new_n501), .B2(new_n507), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(KEYINPUT45), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n472), .A2(G40), .A3(new_n482), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n966), .A2(KEYINPUT107), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n967), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n971), .B(KEYINPUT108), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n777), .A2(G2067), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  INV_X1    g551(.A(G2067), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n774), .B2(new_n776), .ZN(new_n978));
  OR3_X1    g553(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n976), .B1(new_n975), .B2(new_n978), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n974), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n974), .A2(G1996), .A3(new_n721), .ZN(new_n982));
  INV_X1    g557(.A(G1996), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n969), .A2(new_n983), .A3(new_n970), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n721), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n800), .B(new_n804), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n973), .B(new_n986), .C1(new_n974), .C2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n472), .A2(G40), .A3(new_n482), .ZN(new_n989));
  INV_X1    g564(.A(G1384), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n479), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT3), .B1(new_n479), .B2(G2104), .ZN(new_n992));
  OAI211_X1 g567(.A(G138), .B(new_n475), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n993), .A2(KEYINPUT4), .B1(new_n496), .B2(new_n497), .ZN(new_n994));
  OAI211_X1 g569(.A(G126), .B(G2105), .C1(new_n991), .C2(new_n992), .ZN(new_n995));
  INV_X1    g570(.A(new_n505), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT71), .B(G114), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n996), .B1(new_n997), .B2(G2105), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n995), .B1(new_n998), .B2(new_n463), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n990), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n989), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n508), .A2(new_n1003), .A3(KEYINPUT45), .A4(new_n990), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT45), .B(new_n990), .C1(new_n994), .C2(new_n999), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT110), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1971), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT111), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n968), .A2(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1000), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n989), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n729), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1007), .A2(new_n1016), .A3(new_n1008), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1010), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G303), .A2(G8), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT55), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(G8), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n970), .A2(new_n968), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n588), .A2(G1981), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT113), .B(G1981), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n582), .A2(new_n583), .A3(new_n587), .A4(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(KEYINPUT49), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(new_n1027), .A3(G8), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT49), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT114), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1000), .A2(new_n989), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1029), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1027), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n578), .A2(G1976), .A3(new_n579), .A4(new_n580), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(G8), .C1(new_n1000), .C2(new_n989), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G288), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1039), .A2(KEYINPUT52), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1040), .A2(new_n1046), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1037), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1020), .B1(new_n1051), .B2(new_n1032), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1022), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n970), .B1(new_n968), .B2(KEYINPUT45), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1005), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n744), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT50), .B1(new_n508), .B2(new_n990), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n1012), .B(G1384), .C1(new_n501), .C2(new_n507), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n737), .B(new_n970), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1059), .A3(G168), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(KEYINPUT120), .A3(G8), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT51), .ZN(new_n1062));
  AOI21_X1  g637(.A(G168), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(KEYINPUT51), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1063), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1062), .B1(new_n1066), .B2(new_n1032), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n1068));
  INV_X1    g643(.A(G2078), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1002), .A2(new_n1006), .A3(new_n1069), .A4(new_n1004), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n970), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n750), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1072), .B(new_n1074), .C1(new_n1075), .C2(new_n1070), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1068), .B1(new_n1076), .B2(G171), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT125), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1002), .A2(new_n1069), .A3(new_n1005), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1002), .A2(KEYINPUT121), .A3(new_n1069), .A4(new_n1005), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(KEYINPUT53), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1070), .A2(new_n1071), .B1(new_n1073), .B2(new_n750), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(G301), .A3(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1077), .A2(new_n1078), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1078), .B1(new_n1077), .B2(new_n1085), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1053), .B(new_n1067), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT56), .B(G2072), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1002), .A2(new_n1006), .A3(new_n1004), .A4(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1014), .B2(G1956), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G299), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT115), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(G299), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1348), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1073), .A2(new_n1098), .B1(new_n977), .B2(new_n1031), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n615), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1097), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n983), .A2(new_n1002), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT116), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1000), .B2(new_n989), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(KEYINPUT117), .B(new_n1106), .C1(new_n1000), .C2(new_n989), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n556), .B1(new_n1104), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(KEYINPUT59), .B(new_n556), .C1(new_n1104), .C2(new_n1111), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1099), .A2(KEYINPUT60), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1031), .A2(new_n977), .ZN(new_n1118));
  OAI211_X1 g693(.A(KEYINPUT60), .B(new_n1118), .C1(new_n1014), .C2(G1348), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT119), .B1(new_n1119), .B2(new_n615), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1099), .A2(new_n1121), .A3(KEYINPUT60), .A4(new_n625), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n615), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1116), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1002), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1126));
  INV_X1    g701(.A(G1956), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1126), .A2(new_n1089), .B1(new_n1127), .B2(new_n1073), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1096), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT61), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1091), .A2(KEYINPUT118), .A3(new_n1096), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT118), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1097), .A2(KEYINPUT61), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1103), .B1(new_n1125), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1137), .B1(new_n1138), .B2(G171), .ZN(new_n1139));
  AOI211_X1 g714(.A(KEYINPUT123), .B(G301), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(G171), .B1(new_n1073), .B2(new_n750), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1142), .B(new_n1072), .C1(new_n1075), .C2(new_n1070), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT124), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT54), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1088), .A2(new_n1136), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1061), .A2(KEYINPUT51), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(G286), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1032), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1147), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1062), .B(KEYINPUT62), .C1(new_n1066), .C2(new_n1032), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1141), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(new_n1156), .A3(new_n1053), .ZN(new_n1157));
  AOI211_X1 g732(.A(new_n1032), .B(G286), .C1(new_n1056), .C2(new_n1059), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1022), .A2(new_n1050), .A3(new_n1052), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1018), .A2(G8), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1020), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1158), .A2(KEYINPUT63), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n1022), .A4(new_n1050), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1022), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1037), .A2(new_n1042), .A3(new_n818), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1026), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1167), .A2(new_n1050), .B1(new_n1169), .B2(new_n1033), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1157), .A2(new_n1166), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n988), .B1(new_n1146), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n986), .B1(new_n974), .B2(new_n987), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n965), .A2(new_n970), .A3(new_n969), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT48), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n801), .A2(new_n804), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n986), .A2(new_n1176), .B1(G2067), .B2(new_n777), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1173), .A2(new_n1175), .B1(new_n1177), .B2(new_n974), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n984), .B(KEYINPUT46), .Z(new_n1179));
  NAND2_X1  g754(.A1(new_n974), .A2(new_n721), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n981), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n981), .A2(KEYINPUT126), .A3(new_n1180), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1179), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT47), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1178), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1172), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g766(.A1(new_n955), .A2(new_n959), .ZN(new_n1193));
  NOR2_X1   g767(.A1(G401), .A2(new_n461), .ZN(new_n1194));
  NAND4_X1  g768(.A1(new_n683), .A2(new_n684), .A3(new_n703), .A4(new_n1194), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n1195), .B1(new_n879), .B2(new_n883), .ZN(new_n1196));
  AND2_X1   g770(.A1(new_n1193), .A2(new_n1196), .ZN(G308));
  NAND2_X1  g771(.A1(new_n1193), .A2(new_n1196), .ZN(G225));
endmodule


