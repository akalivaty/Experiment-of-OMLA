//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AND2_X1   g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G116), .ZN(new_n222));
  INV_X1    g0022(.A(G270), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n202), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n215), .B1(new_n217), .B2(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND2_X1  g0046(.A1(G1), .A2(G13), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n247), .B1(G33), .B2(G41), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G226), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n253), .B1(new_n216), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n250), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G222), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n259), .B1(new_n260), .B2(new_n258), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n257), .B1(new_n264), .B2(new_n248), .ZN(new_n265));
  INV_X1    g0065(.A(G200), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(G190), .B2(new_n265), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n247), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n273), .A2(new_n274), .B1(new_n202), .B2(new_n270), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n210), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n276), .A2(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(G20), .B2(new_n203), .ZN(new_n282));
  INV_X1    g0082(.A(new_n272), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n275), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT67), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT9), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n287), .B(new_n275), .C1(new_n282), .C2(new_n283), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n286), .B1(new_n285), .B2(new_n288), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n268), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT10), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT10), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n268), .B(new_n293), .C1(new_n289), .C2(new_n290), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G97), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n296), .B(new_n297), .C1(new_n262), .C2(new_n221), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n248), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT13), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n251), .A2(G238), .B1(new_n250), .B2(new_n255), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n303));
  OAI21_X1  g0103(.A(G200), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n269), .A2(G68), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT12), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT68), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n306), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n308), .B2(new_n309), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n209), .A2(G20), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n273), .A2(G68), .A3(new_n312), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n280), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n277), .A2(new_n260), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n272), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n316), .A2(KEYINPUT11), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(KEYINPUT11), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n311), .B(new_n313), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n299), .A2(new_n301), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(G190), .A3(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n304), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(G169), .B1(new_n302), .B2(new_n303), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT14), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n322), .A2(G179), .A3(new_n323), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n329), .B(G169), .C1(new_n302), .C2(new_n303), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n325), .B1(new_n331), .B2(new_n319), .ZN(new_n332));
  INV_X1    g0132(.A(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT3), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G33), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n334), .A2(new_n336), .A3(G232), .A4(new_n261), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n334), .A2(new_n336), .A3(G238), .A4(G1698), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n338), .C1(new_n206), .C2(new_n258), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n248), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n251), .A2(G244), .B1(new_n250), .B2(new_n255), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n340), .A2(KEYINPUT66), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT66), .B1(new_n340), .B2(new_n341), .ZN(new_n343));
  OAI21_X1  g0143(.A(G190), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n341), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT66), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT66), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(G200), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n276), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n279), .B1(G20), .B2(G77), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT15), .B(G87), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n277), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n272), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n312), .A2(G77), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n273), .A2(new_n356), .B1(new_n260), .B2(new_n270), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n344), .A2(new_n349), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(KEYINPUT65), .A2(G179), .ZN(new_n359));
  NOR2_X1   g0159(.A1(KEYINPUT65), .A2(G179), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n342), .B2(new_n343), .ZN(new_n362));
  INV_X1    g0162(.A(G169), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n347), .A2(new_n363), .A3(new_n348), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n354), .A2(new_n357), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n265), .A2(new_n361), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(new_n284), .C1(G169), .C2(new_n265), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n295), .A2(new_n332), .A3(new_n367), .A4(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n276), .B1(new_n209), .B2(G20), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(new_n273), .B1(new_n270), .B2(new_n276), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n334), .A2(new_n336), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT7), .B1(new_n374), .B2(new_n210), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  AOI211_X1 g0176(.A(new_n376), .B(G20), .C1(new_n334), .C2(new_n336), .ZN(new_n377));
  OAI21_X1  g0177(.A(G68), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G58), .ZN(new_n379));
  INV_X1    g0179(.A(G68), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(G20), .B1(new_n381), .B2(new_n201), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n279), .A2(G159), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n283), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n378), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n373), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n334), .A2(new_n336), .A3(G226), .A4(G1698), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n334), .A2(new_n336), .A3(G223), .A4(new_n261), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n248), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n216), .A2(new_n254), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(G232), .A3(new_n249), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n256), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n395), .A2(new_n398), .A3(new_n361), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n256), .A2(new_n397), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n248), .B2(new_n394), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n399), .B1(new_n401), .B2(G169), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT18), .B1(new_n390), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n376), .B1(new_n258), .B2(G20), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n374), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n380), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n387), .B1(new_n406), .B2(new_n384), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n389), .A2(new_n407), .A3(new_n272), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n402), .B1(new_n408), .B2(new_n372), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G190), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n395), .A2(new_n398), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n401), .B2(G200), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n414), .A3(new_n372), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n408), .A2(new_n414), .A3(KEYINPUT17), .A4(new_n372), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n403), .A2(new_n411), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  XOR2_X1   g0219(.A(new_n419), .B(KEYINPUT69), .Z(new_n420));
  NAND4_X1  g0220(.A1(new_n334), .A2(new_n336), .A3(G257), .A4(new_n261), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT75), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n258), .A2(KEYINPUT75), .A3(G257), .A4(new_n261), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n374), .A2(G303), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n258), .A2(G264), .A3(G1698), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n423), .A2(new_n424), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n248), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n209), .A2(G45), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT5), .B(G41), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n248), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n430), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n432), .A2(G270), .B1(new_n434), .B2(new_n255), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n209), .A2(G33), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n269), .A2(new_n437), .A3(new_n247), .A4(new_n271), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G116), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(G116), .B2(new_n270), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G283), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT71), .B(G97), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n210), .B(new_n441), .C1(new_n442), .C2(G33), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n271), .A2(new_n247), .B1(G20), .B2(new_n222), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT20), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n205), .A2(KEYINPUT71), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT71), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G97), .ZN(new_n448));
  AOI21_X1  g0248(.A(G33), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n441), .A2(new_n210), .ZN(new_n450));
  OAI211_X1 g0250(.A(KEYINPUT20), .B(new_n444), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n440), .B1(new_n445), .B2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n436), .A2(KEYINPUT21), .A3(new_n453), .A4(G169), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n255), .A2(new_n430), .A3(new_n431), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n433), .A2(new_n396), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n223), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(new_n248), .B2(new_n427), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(G179), .A3(new_n453), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT21), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n436), .A2(G169), .A3(new_n453), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n460), .A2(KEYINPUT76), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT76), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n454), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n453), .B1(new_n436), .B2(G200), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n412), .B2(new_n436), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n352), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(new_n269), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT19), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n442), .B2(new_n277), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G87), .A2(G107), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n446), .A2(new_n448), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n210), .B1(new_n297), .B2(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n258), .A2(new_n210), .A3(G68), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n472), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n470), .B1(new_n478), .B2(new_n272), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n352), .B(KEYINPUT74), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(new_n273), .A3(new_n437), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n258), .A2(G244), .A3(G1698), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G116), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n334), .A2(new_n336), .A3(G238), .A4(new_n261), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n248), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n429), .A2(G250), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n396), .A2(new_n488), .B1(new_n255), .B2(new_n430), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n361), .A3(new_n489), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n487), .A2(new_n489), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n482), .B(new_n490), .C1(new_n491), .C2(G169), .ZN(new_n492));
  INV_X1    g0292(.A(G87), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n438), .A2(new_n493), .ZN(new_n494));
  AOI211_X1 g0294(.A(new_n470), .B(new_n494), .C1(new_n478), .C2(new_n272), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n487), .A2(G190), .A3(new_n489), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n496), .C1(new_n491), .C2(new_n266), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n433), .A2(G264), .A3(new_n396), .ZN(new_n498));
  MUX2_X1   g0298(.A(G250), .B(G257), .S(G1698), .Z(new_n499));
  AOI22_X1  g0299(.A1(new_n499), .A2(new_n258), .B1(G33), .B2(G294), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n498), .B(new_n455), .C1(new_n500), .C2(new_n396), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n501), .A2(new_n412), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(G200), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OR3_X1    g0304(.A1(new_n269), .A2(KEYINPUT25), .A3(G107), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT25), .B1(new_n269), .B2(G107), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n505), .B(new_n506), .C1(new_n206), .C2(new_n438), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT77), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n438), .A2(new_n206), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n510), .A2(KEYINPUT77), .A3(new_n505), .A4(new_n506), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT23), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n210), .B2(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G20), .B2(new_n484), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n334), .A2(new_n336), .A3(new_n210), .A4(G87), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT22), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT22), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n258), .A2(new_n520), .A3(new_n210), .A4(G87), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n517), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n272), .B1(new_n522), .B2(KEYINPUT24), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(new_n521), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n484), .A2(G20), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n514), .B2(new_n515), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT24), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n512), .B1(new_n523), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n492), .B(new_n497), .C1(new_n504), .C2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n501), .A2(new_n363), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n501), .A2(G179), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n530), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n334), .A2(new_n336), .A3(G244), .A4(new_n261), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n258), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n441), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n248), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n433), .A2(G257), .A3(new_n396), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n455), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n361), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n248), .B2(new_n542), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n363), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n446), .B2(new_n448), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT6), .B1(new_n207), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(G20), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n279), .A2(G77), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n556), .B(KEYINPUT70), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n206), .B1(new_n404), .B2(new_n405), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n272), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n438), .A2(G97), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n269), .A2(new_n205), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT72), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n561), .A2(KEYINPUT72), .A3(new_n562), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT73), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n560), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n568), .B1(new_n560), .B2(new_n567), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n550), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n560), .A2(new_n567), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n549), .A2(G190), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n266), .C2(new_n549), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n532), .A2(new_n536), .A3(new_n571), .A4(new_n574), .ZN(new_n575));
  NOR4_X1   g0375(.A1(new_n370), .A2(new_n420), .A3(new_n468), .A4(new_n575), .ZN(G372));
  NOR2_X1   g0376(.A1(new_n420), .A2(new_n370), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT78), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n532), .A2(new_n578), .A3(new_n571), .A4(new_n574), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n571), .A2(new_n574), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT78), .B1(new_n580), .B2(new_n531), .ZN(new_n581));
  INV_X1    g0381(.A(new_n460), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n462), .A2(new_n461), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n536), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT79), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n582), .A2(KEYINPUT79), .A3(new_n583), .A4(new_n536), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n579), .A2(new_n581), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n560), .A2(new_n567), .ZN(new_n589));
  INV_X1    g0389(.A(new_n548), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n363), .B1(new_n543), .B2(new_n546), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT80), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n492), .A2(new_n497), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT26), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n550), .A2(KEYINPUT80), .A3(new_n589), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n492), .A2(new_n497), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT26), .B1(new_n571), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n598), .A2(new_n492), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n588), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n577), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g0403(.A(new_n603), .B(KEYINPUT81), .Z(new_n604));
  XNOR2_X1  g0404(.A(new_n409), .B(KEYINPUT18), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n330), .A2(new_n328), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n322), .A2(new_n323), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n329), .B1(new_n608), .B2(G169), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n319), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n325), .B2(new_n366), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n417), .A2(new_n418), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n295), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n369), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT82), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(KEYINPUT82), .B(new_n369), .C1(new_n613), .C2(new_n614), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n604), .A2(new_n619), .ZN(G369));
  NAND2_X1  g0420(.A1(new_n582), .A2(new_n583), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(G213), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(G343), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n453), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n468), .B2(new_n628), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(G330), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n283), .B1(new_n527), .B2(new_n528), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n528), .B2(new_n527), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(new_n512), .A3(new_n502), .A4(new_n503), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n530), .A2(new_n627), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n536), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n627), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n637), .B1(new_n536), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n536), .A2(new_n627), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n627), .B1(new_n463), .B2(new_n465), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n635), .A2(new_n536), .A3(new_n636), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n640), .A2(new_n644), .ZN(G399));
  INV_X1    g0445(.A(new_n213), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(G41), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n474), .A2(G116), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n647), .A2(new_n209), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n219), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n650), .A2(KEYINPUT83), .B1(new_n651), .B2(new_n647), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(KEYINPUT83), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT28), .ZN(new_n654));
  INV_X1    g0454(.A(G330), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n463), .A2(new_n465), .A3(new_n467), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n580), .A2(new_n531), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n656), .A2(new_n536), .A3(new_n657), .A4(new_n638), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n487), .A2(new_n489), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n549), .B1(KEYINPUT84), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n501), .A2(new_n361), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n458), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n659), .A2(KEYINPUT84), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT30), .ZN(new_n665));
  INV_X1    g0465(.A(new_n500), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n666), .A2(new_n248), .B1(G264), .B2(new_n432), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n491), .A2(new_n549), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n458), .A2(G179), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n665), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n667), .A2(new_n487), .A3(new_n489), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n428), .A2(G179), .A3(new_n435), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(KEYINPUT30), .A3(new_n672), .A4(new_n549), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n664), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n627), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT31), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT31), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n677), .A3(new_n627), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n655), .B1(new_n658), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n602), .A2(new_n638), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT26), .ZN(new_n685));
  INV_X1    g0485(.A(new_n570), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n560), .A2(new_n567), .A3(new_n568), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n595), .A2(new_n550), .A3(new_n688), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n685), .B(new_n492), .C1(KEYINPUT26), .C2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n463), .A2(new_n465), .A3(new_n536), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n657), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI211_X1 g0493(.A(KEYINPUT29), .B(new_n638), .C1(new_n690), .C2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n680), .B1(new_n683), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n654), .B1(new_n695), .B2(G1), .ZN(G364));
  AND2_X1   g0496(.A1(new_n210), .A2(G13), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n209), .B1(new_n697), .B2(G45), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n647), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n632), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(G330), .B2(new_n630), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n646), .A2(new_n374), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G355), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(G116), .B2(new_n213), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n646), .A2(new_n258), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G45), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n651), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n242), .A2(new_n708), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n705), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G13), .A2(G33), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n247), .B1(G20), .B2(new_n363), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n700), .B1(new_n711), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n210), .A2(new_n266), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n547), .A2(G190), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n210), .A2(new_n412), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n547), .A2(new_n266), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI22_X1  g0524(.A1(G50), .A2(new_n721), .B1(new_n724), .B2(G58), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n210), .A2(G190), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n547), .A2(new_n266), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n260), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT85), .Z(new_n729));
  NOR2_X1   g0529(.A1(new_n266), .A2(G179), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n722), .A2(new_n730), .ZN(new_n732));
  OAI221_X1 g0532(.A(new_n258), .B1(new_n731), .B2(new_n206), .C1(new_n493), .C2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G179), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n726), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G159), .ZN(new_n736));
  OR3_X1    g0536(.A1(new_n735), .A2(KEYINPUT32), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT32), .B1(new_n735), .B2(new_n736), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n210), .B1(new_n734), .B2(G190), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G97), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n737), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n547), .A2(new_n412), .A3(new_n719), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n733), .B(new_n742), .C1(G68), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n729), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n732), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n747), .A2(KEYINPUT87), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(KEYINPUT87), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G303), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT33), .B(G317), .ZN(new_n752));
  INV_X1    g0552(.A(new_n727), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n744), .A2(new_n752), .B1(new_n753), .B2(G311), .ZN(new_n754));
  INV_X1    g0554(.A(G294), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n739), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G283), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n374), .B1(new_n731), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n735), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n756), .B(new_n758), .C1(G329), .C2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(KEYINPUT86), .B(G326), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G322), .A2(new_n724), .B1(new_n721), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n751), .A2(new_n754), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT88), .B1(new_n746), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n715), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n746), .A2(KEYINPUT88), .A3(new_n763), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n718), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n714), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n630), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n702), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(G396));
  OAI21_X1  g0572(.A(new_n258), .B1(new_n731), .B2(new_n380), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(G132), .B2(new_n759), .ZN(new_n774));
  INV_X1    g0574(.A(new_n750), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n774), .B1(new_n379), .B2(new_n739), .C1(new_n775), .C2(new_n202), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G137), .A2(new_n721), .B1(new_n744), .B2(G150), .ZN(new_n778));
  XNOR2_X1  g0578(.A(KEYINPUT92), .B(G143), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n778), .B1(new_n736), .B2(new_n727), .C1(new_n723), .C2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT34), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n741), .B1(new_n723), .B2(new_n755), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT90), .Z(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n374), .B1(new_n735), .B2(new_n784), .C1(new_n493), .C2(new_n731), .ZN(new_n785));
  XOR2_X1   g0585(.A(KEYINPUT89), .B(G283), .Z(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n785), .B1(new_n744), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n750), .A2(G107), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G303), .A2(new_n721), .B1(new_n753), .B2(G116), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n783), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT91), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n777), .A2(new_n781), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n715), .ZN(new_n795));
  INV_X1    g0595(.A(new_n700), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n715), .A2(new_n712), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n796), .B1(new_n260), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n365), .A2(new_n627), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT94), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n364), .A2(new_n365), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT95), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n801), .A2(new_n802), .A3(new_n362), .A4(new_n627), .ZN(new_n803));
  OAI21_X1  g0603(.A(KEYINPUT95), .B1(new_n366), .B2(new_n638), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n367), .A2(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n795), .B(new_n798), .C1(new_n713), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n681), .A2(new_n805), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n627), .B1(new_n588), .B2(new_n601), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n806), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n680), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT96), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(KEYINPUT96), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n808), .A2(new_n680), .A3(new_n810), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n814), .A2(new_n796), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n807), .B1(new_n813), .B2(new_n816), .ZN(G384));
  NOR2_X1   g0617(.A1(new_n217), .A2(new_n222), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n552), .A2(new_n554), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT97), .Z(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT35), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(new_n822), .B2(new_n821), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT36), .ZN(new_n825));
  OR3_X1    g0625(.A1(new_n219), .A2(new_n260), .A3(new_n381), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n202), .A2(G68), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n209), .B(G13), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n325), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n319), .A2(new_n627), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n610), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n319), .B(new_n627), .C1(new_n331), .C2(new_n325), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n803), .A2(new_n804), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n367), .A2(new_n800), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n832), .A2(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n575), .A2(new_n468), .A3(new_n627), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n674), .A2(new_n677), .A3(new_n627), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n677), .B1(new_n674), .B2(new_n627), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n836), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n408), .A2(new_n372), .ZN(new_n843));
  INV_X1    g0643(.A(new_n402), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n625), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n845), .A2(new_n847), .A3(new_n415), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT37), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n408), .A2(new_n372), .A3(new_n414), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n409), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n852), .A3(new_n847), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n847), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n419), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n854), .A2(new_n856), .A3(KEYINPUT38), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT38), .B1(new_n854), .B2(new_n856), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT98), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT98), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n852), .B1(new_n851), .B2(new_n847), .ZN(new_n862));
  AND4_X1   g0662(.A1(new_n852), .A2(new_n845), .A3(new_n847), .A4(new_n415), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n847), .B1(new_n605), .B2(new_n612), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n854), .A2(new_n856), .A3(KEYINPUT38), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n860), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n842), .B1(new_n859), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT99), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT40), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT98), .B1(new_n857), .B2(new_n858), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n866), .A2(new_n860), .A3(new_n867), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n841), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT99), .B1(new_n875), .B2(KEYINPUT40), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n871), .B1(new_n866), .B2(new_n867), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n842), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT100), .Z(new_n881));
  OAI21_X1  g0681(.A(new_n577), .B1(new_n837), .B2(new_n840), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n655), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n881), .B2(new_n883), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n866), .A2(new_n867), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT39), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n866), .A2(KEYINPUT39), .A3(new_n867), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n331), .A2(new_n319), .A3(new_n638), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n890), .A2(new_n891), .B1(new_n605), .B2(new_n846), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n832), .A2(new_n833), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n366), .A2(new_n627), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n895), .B1(new_n810), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n873), .A2(new_n874), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n683), .A2(new_n577), .A3(new_n694), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n619), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n901), .B(new_n903), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n885), .A2(new_n904), .B1(new_n209), .B2(new_n697), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT101), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n885), .A2(new_n904), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n905), .A2(KEYINPUT101), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n829), .B1(new_n908), .B2(new_n909), .ZN(G367));
  NAND2_X1  g0710(.A1(new_n706), .A2(new_n238), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(new_n716), .C1(new_n213), .C2(new_n352), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n750), .A2(KEYINPUT46), .A3(G116), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT108), .Z(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT46), .B1(new_n747), .B2(G116), .ZN(new_n915));
  INV_X1    g0715(.A(G317), .ZN(new_n916));
  OAI221_X1 g0716(.A(new_n374), .B1(new_n735), .B2(new_n916), .C1(new_n442), .C2(new_n731), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n915), .B(new_n917), .C1(G107), .C2(new_n740), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n743), .A2(new_n755), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n720), .A2(new_n784), .ZN(new_n920));
  INV_X1    g0720(.A(G303), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n723), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n727), .A2(new_n786), .ZN(new_n923));
  NOR4_X1   g0723(.A1(new_n919), .A2(new_n920), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n914), .A2(new_n918), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT109), .ZN(new_n926));
  AOI22_X1  g0726(.A1(G150), .A2(new_n724), .B1(new_n753), .B2(G50), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n927), .B1(new_n736), .B2(new_n743), .C1(new_n720), .C2(new_n779), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n739), .A2(new_n380), .ZN(new_n929));
  INV_X1    g0729(.A(G137), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n258), .B1(new_n735), .B2(new_n930), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n732), .A2(new_n379), .B1(new_n731), .B2(new_n260), .ZN(new_n932));
  NOR4_X1   g0732(.A1(new_n928), .A2(new_n929), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n926), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT47), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n700), .B(new_n912), .C1(new_n935), .C2(new_n765), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n937), .A2(KEYINPUT110), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n495), .A2(new_n638), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT102), .Z(new_n940));
  NOR2_X1   g0740(.A1(new_n940), .A2(new_n595), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n492), .B2(new_n940), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n714), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n937), .A2(KEYINPUT110), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n938), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT107), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n571), .B(new_n574), .C1(new_n572), .C2(new_n638), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n550), .A2(new_n589), .A3(new_n627), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT105), .B1(new_n644), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n460), .A2(KEYINPUT76), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(new_n465), .A3(new_n583), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n643), .A3(new_n638), .ZN(new_n954));
  INV_X1    g0754(.A(new_n641), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT105), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n948), .A2(new_n949), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n951), .A2(KEYINPUT44), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT44), .ZN(new_n961));
  AOI211_X1 g0761(.A(KEYINPUT105), .B(new_n950), .C1(new_n954), .C2(new_n955), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT104), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n644), .A2(new_n965), .A3(new_n950), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n954), .A2(new_n955), .A3(new_n950), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT104), .ZN(new_n968));
  XNOR2_X1  g0768(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n969), .B1(new_n966), .B2(new_n968), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n960), .B(new_n964), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n640), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n966), .A2(new_n968), .ZN(new_n975));
  INV_X1    g0775(.A(new_n969), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n979), .A2(new_n640), .A3(new_n960), .A4(new_n964), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n642), .A2(new_n639), .ZN(new_n981));
  INV_X1    g0781(.A(new_n954), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(new_n631), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n631), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n680), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n694), .B1(KEYINPUT29), .B2(new_n809), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n974), .A2(new_n980), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n695), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n647), .B(KEYINPUT41), .Z(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(KEYINPUT106), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n990), .B2(new_n695), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT106), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n995), .A2(new_n698), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n982), .A2(new_n950), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n571), .B1(new_n958), .B2(new_n536), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(KEYINPUT42), .A2(new_n1000), .B1(new_n1001), .B2(new_n638), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT42), .B2(new_n1000), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT43), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n943), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n640), .A2(new_n958), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1009));
  AND3_X1   g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1008), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n947), .B1(new_n999), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n698), .B1(new_n996), .B2(new_n997), .ZN(new_n1014));
  AOI211_X1 g0814(.A(KEYINPUT106), .B(new_n992), .C1(new_n990), .C2(new_n695), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n947), .B(new_n1012), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n946), .B1(new_n1013), .B2(new_n1017), .ZN(G387));
  AOI21_X1  g0818(.A(new_n707), .B1(new_n235), .B2(G45), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n649), .B2(new_n703), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT50), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n350), .B2(new_n202), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n276), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n708), .B1(new_n380), .B2(new_n260), .ZN(new_n1024));
  NOR4_X1   g0824(.A1(new_n649), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1020), .A2(new_n1025), .B1(G107), .B2(new_n213), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n796), .B1(new_n1026), .B2(new_n716), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n639), .B2(new_n769), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n380), .A2(new_n727), .B1(new_n743), .B2(new_n276), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT111), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n258), .B1(new_n731), .B2(new_n205), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n732), .A2(new_n260), .B1(new_n735), .B2(new_n278), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n721), .C2(G159), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n724), .A2(G50), .B1(new_n480), .B2(new_n740), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1030), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n786), .A2(new_n739), .B1(new_n732), .B2(new_n755), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G311), .A2(new_n744), .B1(new_n721), .B2(G322), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n921), .B2(new_n727), .C1(new_n916), .C2(new_n723), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT48), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n1039), .B2(new_n1038), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT49), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(KEYINPUT112), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n374), .B1(new_n731), .B2(new_n222), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n759), .B2(new_n761), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1042), .A2(KEYINPUT112), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1035), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT113), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n765), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1028), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n699), .B2(new_n986), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n695), .A2(new_n986), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n989), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n647), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1053), .B1(new_n1054), .B2(new_n1056), .ZN(G393));
  INV_X1    g0857(.A(new_n974), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n980), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1060), .A2(new_n647), .A3(new_n990), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n974), .A2(new_n980), .A3(new_n699), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n716), .B1(new_n213), .B2(new_n442), .C1(new_n707), .C2(new_n245), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n700), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n784), .A2(new_n723), .B1(new_n720), .B2(new_n916), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT52), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n374), .B1(new_n731), .B2(new_n206), .ZN(new_n1067));
  INV_X1    g0867(.A(G322), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n786), .A2(new_n732), .B1(new_n735), .B2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(G116), .C2(new_n740), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G303), .A2(new_n744), .B1(new_n753), .B2(G294), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1066), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n278), .A2(new_n720), .B1(new_n723), .B2(new_n736), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT51), .Z(new_n1074));
  OAI21_X1  g0874(.A(new_n258), .B1(new_n731), .B2(new_n493), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n732), .A2(new_n380), .B1(new_n735), .B2(new_n779), .ZN(new_n1076));
  OR3_X1    g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n753), .A2(new_n350), .B1(G77), .B2(new_n740), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n202), .B2(new_n743), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT114), .Z(new_n1080));
  OAI21_X1  g0880(.A(new_n1072), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1064), .B1(new_n1081), .B2(new_n715), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n769), .B2(new_n950), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1061), .A2(new_n1062), .A3(new_n1083), .ZN(G390));
  NAND3_X1  g0884(.A1(new_n680), .A2(new_n806), .A3(new_n894), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n627), .B(new_n805), .C1(new_n588), .C2(new_n601), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n894), .B1(new_n1087), .B2(new_n896), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1088), .A2(new_n891), .B1(new_n888), .B2(new_n889), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n886), .A2(new_n891), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n684), .A2(KEYINPUT26), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n492), .B1(new_n689), .B2(KEYINPUT26), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n627), .B1(new_n1093), .B2(new_n692), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n806), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n897), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1090), .B1(new_n1096), .B2(new_n894), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1086), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n891), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n890), .B1(new_n898), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n896), .B1(new_n1094), .B2(new_n806), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n886), .B(new_n891), .C1(new_n1101), .C2(new_n895), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1085), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1098), .A2(new_n699), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT116), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1104), .B(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(G330), .B(new_n806), .C1(new_n837), .C2(new_n840), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n895), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT115), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1101), .A2(new_n1108), .A3(new_n1085), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1101), .A2(new_n1108), .A3(new_n1085), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1112), .A2(KEYINPUT115), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1108), .A2(new_n1085), .B1(new_n810), .B2(new_n897), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1111), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n577), .A2(new_n680), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n902), .A2(new_n619), .A3(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1116), .A2(new_n1098), .A3(new_n1103), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1112), .A2(KEYINPUT115), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1118), .B(new_n1110), .C1(new_n1114), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1119), .A2(new_n1123), .A3(new_n647), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n797), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n700), .B1(new_n350), .B2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT117), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1128), .A2(new_n753), .B1(new_n724), .B2(G132), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n930), .B2(new_n743), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n732), .A2(new_n278), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n720), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n731), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n374), .B1(new_n1135), .B2(G50), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n759), .A2(G125), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(new_n1137), .C1(new_n736), .C2(new_n739), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1130), .A2(new_n1134), .A3(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT118), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n775), .A2(new_n493), .B1(new_n222), .B2(new_n723), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G283), .B2(new_n721), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n374), .B1(new_n735), .B2(new_n755), .C1(new_n380), .C2(new_n731), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G77), .B2(new_n740), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n206), .A2(new_n743), .B1(new_n727), .B2(new_n442), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT119), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1142), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT120), .B1(new_n1140), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1148), .A2(new_n765), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1140), .A2(KEYINPUT120), .A3(new_n1147), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1126), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n890), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1151), .B1(new_n1152), .B2(new_n713), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1106), .A2(new_n1124), .A3(new_n1153), .ZN(G378));
  NAND2_X1  g0954(.A1(new_n295), .A2(new_n369), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n625), .B1(new_n285), .B2(new_n288), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n879), .A2(G330), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1165), .B1(new_n877), .B2(new_n1167), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1166), .B(new_n1164), .C1(new_n872), .C2(new_n876), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n901), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n902), .A2(new_n619), .A3(new_n1117), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT123), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n870), .B1(new_n869), .B2(new_n871), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n875), .A2(KEYINPUT99), .A3(KEYINPUT40), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1167), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1164), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n901), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n877), .A2(new_n1167), .A3(new_n1165), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1170), .A2(new_n1174), .A3(new_n1181), .A4(KEYINPUT57), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n901), .A2(KEYINPUT122), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT122), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n893), .B2(new_n900), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1178), .A2(new_n1180), .A3(new_n1186), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1184), .A2(new_n1187), .B1(new_n1119), .B2(new_n1173), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n647), .B(new_n1182), .C1(new_n1188), .C2(KEYINPUT57), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1165), .A2(new_n712), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n700), .B1(G50), .B2(new_n1125), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n258), .A2(G41), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n480), .A2(new_n753), .B1(new_n721), .B2(G116), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G97), .A2(new_n744), .B1(new_n724), .B2(G107), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1193), .B1(new_n379), .B2(new_n731), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n732), .A2(new_n260), .B1(new_n735), .B2(new_n757), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1198), .A2(new_n1199), .A3(new_n929), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1196), .A2(new_n1197), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT58), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1195), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT121), .B(G124), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G33), .B(G41), .C1(new_n759), .C2(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G132), .A2(new_n744), .B1(new_n753), .B2(G137), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G125), .A2(new_n721), .B1(new_n724), .B2(G128), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1128), .A2(new_n747), .B1(G150), .B2(new_n740), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT59), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1205), .B1(new_n736), .B2(new_n731), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1209), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1203), .B1(new_n1202), .B2(new_n1201), .C1(new_n1211), .C2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1192), .B1(new_n1214), .B2(new_n715), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1190), .A2(new_n699), .B1(new_n1191), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1189), .A2(new_n1216), .ZN(G375));
  OAI21_X1  g1017(.A(new_n1110), .B1(new_n1121), .B2(new_n1114), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1171), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(new_n993), .A3(new_n1122), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n895), .A2(new_n712), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n700), .B1(G68), .B2(new_n1125), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n757), .A2(new_n723), .B1(new_n720), .B2(new_n755), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n750), .B2(G97), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n374), .B1(new_n735), .B2(new_n921), .C1(new_n260), .C2(new_n731), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n480), .B2(new_n740), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G116), .A2(new_n744), .B1(new_n753), .B2(G107), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n750), .A2(G159), .B1(G128), .B2(new_n759), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT124), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G132), .A2(new_n721), .B1(new_n753), .B2(G150), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n724), .A2(G137), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n258), .B1(new_n731), .B2(new_n379), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G50), .B2(new_n740), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n744), .A2(new_n1128), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1231), .A2(new_n1232), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1228), .B1(new_n1230), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1222), .B1(new_n1237), .B2(new_n715), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1116), .A2(new_n699), .B1(new_n1221), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1220), .A2(new_n1239), .ZN(G381));
  OR2_X1    g1040(.A1(G393), .A2(G396), .ZN(new_n1241));
  OR4_X1    g1041(.A1(G384), .A2(new_n1241), .A3(G390), .A4(G381), .ZN(new_n1242));
  OR4_X1    g1042(.A1(G387), .A2(new_n1242), .A3(G378), .A4(G375), .ZN(G407));
  AND3_X1   g1043(.A1(new_n1106), .A2(new_n1124), .A3(new_n1153), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n626), .ZN(new_n1245));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(G375), .C2(new_n1245), .ZN(G409));
  NAND3_X1  g1046(.A1(new_n1189), .A2(G378), .A3(new_n1216), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1190), .A2(new_n993), .A3(new_n1174), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1170), .A2(new_n1181), .A3(new_n699), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1191), .A2(new_n1215), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1244), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1247), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1122), .A2(KEYINPUT60), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1256), .A2(new_n1219), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n647), .B1(new_n1256), .B2(new_n1219), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1239), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G384), .B(new_n1239), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1247), .A2(new_n1252), .A3(KEYINPUT125), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n626), .A2(G213), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1255), .A2(new_n1264), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1261), .A2(KEYINPUT63), .A3(new_n1262), .ZN(new_n1270));
  AND4_X1   g1070(.A1(KEYINPUT126), .A2(new_n1253), .A3(new_n1266), .A4(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1266), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1247), .B2(new_n1252), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT126), .B1(new_n1273), .B2(new_n1270), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1255), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1272), .A2(G2897), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1261), .A2(new_n1262), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1276), .A2(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(G393), .B(new_n771), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT107), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1016), .ZN(new_n1287));
  AOI21_X1  g1087(.A(G390), .B1(new_n1287), .B2(new_n946), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n946), .ZN(new_n1289));
  INV_X1    g1089(.A(G390), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1289), .B(new_n1290), .C1(new_n1286), .C2(new_n1016), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1284), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G387), .A2(new_n1290), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1287), .A2(new_n946), .A3(G390), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1283), .A3(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1292), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1269), .A2(new_n1275), .A3(new_n1282), .A4(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1280), .B2(new_n1273), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1267), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1273), .A2(KEYINPUT62), .A3(new_n1264), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1299), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1292), .A2(new_n1295), .A3(KEYINPUT127), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1298), .B1(new_n1303), .B2(new_n1308), .ZN(G405));
  INV_X1    g1109(.A(new_n1307), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT127), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1247), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G378), .B1(new_n1189), .B2(new_n1216), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1264), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1313), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(new_n1263), .A3(new_n1247), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1310), .A2(new_n1311), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1317), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1319), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1318), .A2(new_n1320), .ZN(G402));
endmodule


