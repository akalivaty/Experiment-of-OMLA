//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g035(.A(G261), .ZN(G325));
  NAND2_X1  g036(.A1(new_n456), .A2(G2106), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n458), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  AND2_X1   g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OR2_X1    g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n472), .A2(G136), .ZN(new_n478));
  INV_X1    g053(.A(G124), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n473), .B1(new_n470), .B2(new_n471), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n478), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g059(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G112), .B2(new_n473), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND3_X1  g064(.A1(new_n466), .A2(G126), .A3(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(G114), .B2(new_n473), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n471), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n473), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n472), .A2(new_n499), .A3(G138), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(G543), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(KEYINPUT72), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT70), .B1(new_n509), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  AND3_X1   g089(.A1(new_n507), .A2(new_n508), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n502), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n507), .A2(new_n508), .A3(new_n514), .A4(new_n519), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n518), .A2(new_n524), .ZN(G166));
  INV_X1    g100(.A(new_n522), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n520), .A2(G51), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n507), .A2(new_n508), .A3(new_n514), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n527), .A2(new_n534), .ZN(G168));
  NAND4_X1  g110(.A1(new_n507), .A2(G64), .A3(new_n508), .A4(new_n514), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n502), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT73), .B(G52), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n520), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n522), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT74), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n544), .B(new_n540), .C1(new_n522), .C2(new_n541), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n538), .B1(new_n543), .B2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n526), .A2(G81), .B1(G43), .B2(new_n520), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n532), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G651), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n520), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n526), .A2(G91), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n507), .A2(G65), .A3(new_n508), .A4(new_n514), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n563), .B1(new_n566), .B2(G651), .ZN(new_n567));
  AOI211_X1 g142(.A(KEYINPUT76), .B(new_n502), .C1(new_n564), .C2(new_n565), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n561), .B(new_n562), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n569), .A2(KEYINPUT77), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(KEYINPUT77), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n543), .A2(new_n545), .ZN(new_n574));
  INV_X1    g149(.A(new_n538), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI211_X1 g151(.A(KEYINPUT78), .B(new_n538), .C1(new_n543), .C2(new_n545), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  OR2_X1    g154(.A1(new_n518), .A2(new_n524), .ZN(G303));
  AOI22_X1  g155(.A1(new_n526), .A2(G87), .B1(G49), .B2(new_n520), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  INV_X1    g157(.A(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n532), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n582), .B1(new_n584), .B2(G651), .ZN(new_n585));
  AOI211_X1 g160(.A(KEYINPUT79), .B(new_n502), .C1(new_n532), .C2(new_n583), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n581), .B1(new_n585), .B2(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n532), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n526), .A2(G86), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n520), .A2(G48), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT80), .ZN(G305));
  XNOR2_X1  g170(.A(KEYINPUT81), .B(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n520), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n522), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n532), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n599), .B1(G651), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n522), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n532), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G301), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G284));
  AOI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(G299), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G280));
  AND2_X1   g195(.A1(new_n607), .A2(new_n611), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT82), .B(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(G860), .B2(new_n622), .ZN(G148));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n466), .A2(new_n474), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT13), .Z(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n472), .A2(G135), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT83), .Z(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n480), .B2(G123), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n631), .A2(G2100), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n632), .A2(new_n641), .A3(new_n642), .A4(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT85), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT84), .B(G2438), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OR3_X1    g226(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n651), .B1(new_n648), .B2(new_n649), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n662), .A3(new_n660), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(new_n665), .A3(G14), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT86), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n668));
  NAND4_X1  g243(.A1(new_n664), .A2(new_n665), .A3(new_n668), .A4(G14), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT18), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n677), .A2(new_n672), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n674), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n673), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n680), .A2(new_n681), .A3(new_n672), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G2096), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT88), .B(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n689), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n689), .B2(new_n695), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT89), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n703), .B(new_n704), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(G229));
  NOR2_X1   g281(.A1(G6), .A2(G16), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT80), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n594), .B(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n707), .B1(new_n709), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT32), .B(G1981), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G23), .ZN(new_n715));
  INV_X1    g290(.A(G288), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n714), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT33), .B(G1976), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(G303), .A2(G16), .ZN(new_n720));
  INV_X1    g295(.A(G22), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(G16), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G1971), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n717), .A2(new_n718), .ZN(new_n724));
  INV_X1    g299(.A(G1971), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n720), .B(new_n725), .C1(G16), .C2(new_n721), .ZN(new_n726));
  AND4_X1   g301(.A1(new_n719), .A2(new_n723), .A3(new_n724), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n713), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(KEYINPUT34), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n713), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT91), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n472), .A2(G131), .ZN(new_n735));
  INV_X1    g310(.A(G119), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(new_n481), .ZN(new_n737));
  NOR2_X1   g312(.A1(G95), .A2(G2105), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT90), .Z(new_n739));
  OAI21_X1  g314(.A(G2104), .B1(new_n473), .B2(G107), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n734), .B1(new_n742), .B2(new_n733), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT35), .B(G1991), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n714), .A2(G24), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n603), .B2(new_n714), .ZN(new_n747));
  INV_X1    g322(.A(G1986), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n745), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AND3_X1   g326(.A1(new_n731), .A2(new_n732), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n732), .B1(new_n731), .B2(new_n751), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n729), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(KEYINPUT36), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n756), .B(new_n729), .C1(new_n752), .C2(new_n753), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n472), .A2(G141), .B1(G105), .B2(new_n474), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n480), .A2(G129), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT26), .Z(new_n762));
  AND3_X1   g337(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(new_n733), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n733), .B2(G32), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G29), .A2(G33), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT25), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n466), .A2(G127), .ZN(new_n771));
  NAND2_X1  g346(.A1(G115), .A2(G2104), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n473), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n770), .B(new_n773), .C1(G139), .C2(new_n472), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n768), .B1(new_n774), .B2(G29), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G2072), .ZN(new_n776));
  INV_X1    g351(.A(G2084), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT24), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n733), .B1(new_n778), .B2(G34), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(KEYINPUT94), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(G34), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n779), .B2(KEYINPUT94), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n476), .A2(new_n733), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n767), .B(new_n776), .C1(new_n777), .C2(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n775), .A2(G2072), .ZN(new_n785));
  NAND2_X1  g360(.A1(G164), .A2(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G27), .B2(G29), .ZN(new_n787));
  INV_X1    g362(.A(G2078), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(G28), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n733), .B1(new_n791), .B2(G28), .ZN(new_n793));
  AND2_X1   g368(.A1(KEYINPUT31), .A2(G11), .ZN(new_n794));
  NOR2_X1   g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n792), .A2(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n639), .B2(G29), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n785), .A2(new_n789), .A3(new_n790), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n733), .A2(G35), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G162), .B2(new_n733), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT29), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n784), .B(new_n798), .C1(G2090), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n714), .A2(G21), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G168), .B2(new_n714), .ZN(new_n804));
  INV_X1    g379(.A(G1966), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n714), .A2(G19), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n553), .B2(new_n714), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G1341), .Z(new_n809));
  NAND3_X1  g384(.A1(new_n802), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n733), .A2(G26), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT93), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT28), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n472), .A2(G140), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n480), .A2(G128), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n473), .A2(G116), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n814), .B(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT92), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n813), .B1(new_n822), .B2(G29), .ZN(new_n823));
  INV_X1    g398(.A(G2067), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n801), .A2(G2090), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(KEYINPUT97), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n621), .A2(G16), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G4), .B2(G16), .ZN(new_n829));
  INV_X1    g404(.A(G1348), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n827), .B(new_n831), .C1(KEYINPUT97), .C2(new_n826), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n714), .A2(G5), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G171), .B2(new_n714), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT95), .Z(new_n835));
  INV_X1    g410(.A(G1961), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n829), .A2(new_n830), .ZN(new_n838));
  NOR4_X1   g413(.A1(new_n810), .A2(new_n832), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n714), .A2(G20), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT23), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n618), .B2(new_n714), .ZN(new_n842));
  INV_X1    g417(.A(G1956), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n783), .A2(new_n777), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n765), .B2(new_n766), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n835), .B2(new_n836), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT96), .Z(new_n848));
  NAND3_X1  g423(.A1(new_n839), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT98), .B1(new_n758), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n852));
  AOI211_X1 g427(.A(new_n852), .B(new_n849), .C1(new_n755), .C2(new_n757), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n851), .A2(new_n853), .ZN(G311));
  NAND2_X1  g429(.A1(new_n758), .A2(new_n850), .ZN(G150));
  NAND2_X1  g430(.A1(new_n621), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n526), .A2(G93), .B1(G55), .B2(new_n520), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n507), .A2(G67), .A3(new_n508), .A4(new_n514), .ZN(new_n859));
  NAND2_X1  g434(.A1(G80), .A2(G543), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G651), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n552), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n547), .A2(new_n858), .A3(new_n551), .A4(new_n862), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n857), .B(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n868), .A2(new_n869), .A3(G860), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n863), .A2(G860), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT99), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT37), .Z(new_n873));
  OR2_X1    g448(.A1(new_n870), .A2(new_n873), .ZN(G145));
  OR2_X1    g449(.A1(new_n737), .A2(new_n741), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n742), .A2(KEYINPUT101), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n629), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n774), .B(new_n763), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  INV_X1    g459(.A(new_n822), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(G164), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n500), .A2(new_n498), .ZN(new_n887));
  INV_X1    g462(.A(G114), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n491), .B1(new_n888), .B2(G2105), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n480), .B2(G126), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n822), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  INV_X1    g468(.A(G118), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n893), .A2(KEYINPUT100), .B1(new_n894), .B2(G2105), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(KEYINPUT100), .B2(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n472), .A2(G142), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n480), .A2(G130), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n886), .A2(new_n892), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n899), .B1(new_n886), .B2(new_n892), .ZN(new_n901));
  OAI22_X1  g476(.A1(new_n883), .A2(new_n884), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n881), .A2(new_n882), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n900), .A2(new_n901), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n881), .A2(new_n882), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n488), .B(G160), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n639), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n907), .B2(new_n909), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g488(.A1(new_n864), .A2(new_n865), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n624), .B(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n566), .A2(G651), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT76), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n566), .A2(new_n563), .A3(G651), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT77), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n920), .A2(new_n921), .A3(new_n561), .A4(new_n562), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n569), .A2(KEYINPUT77), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n922), .A2(new_n621), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n621), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n916), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n612), .B1(new_n570), .B2(new_n571), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n621), .A3(new_n923), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(KEYINPUT41), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n915), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n624), .B(new_n866), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n924), .A2(new_n925), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n930), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(G303), .A2(new_n603), .ZN(new_n936));
  NAND2_X1  g511(.A1(G166), .A2(G290), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(G305), .A2(G288), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n709), .A2(new_n716), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n941), .B2(new_n942), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n935), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n931), .B1(new_n930), .B2(new_n934), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n926), .A2(new_n929), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n932), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n927), .A2(new_n928), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n915), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(KEYINPUT102), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n948), .A2(new_n949), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n947), .A2(new_n955), .A3(G868), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G868), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n863), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n947), .A2(new_n955), .A3(KEYINPUT103), .A4(G868), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(G331));
  XNOR2_X1  g537(.A(G331), .B(KEYINPUT104), .ZN(G295));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n965));
  OAI21_X1  g540(.A(G168), .B1(new_n576), .B2(new_n577), .ZN(new_n966));
  NOR2_X1   g541(.A1(G171), .A2(G168), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n965), .B1(new_n969), .B2(new_n914), .ZN(new_n970));
  AOI211_X1 g545(.A(KEYINPUT105), .B(new_n866), .C1(new_n966), .C2(new_n968), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n966), .A2(new_n866), .A3(new_n968), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n952), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n545), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT71), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n509), .ZN(new_n977));
  NAND2_X1  g552(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n512), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n979), .A2(KEYINPUT72), .B1(new_n510), .B2(new_n513), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n980), .A2(G90), .A3(new_n507), .A4(new_n519), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n544), .B1(new_n981), .B2(new_n540), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n575), .B1(new_n975), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT78), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n574), .A2(new_n573), .A3(new_n575), .ZN(new_n985));
  AOI21_X1  g560(.A(G286), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n914), .B1(new_n986), .B2(new_n967), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n973), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n972), .A2(new_n974), .B1(new_n950), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(KEYINPUT106), .B(new_n964), .C1(new_n989), .C2(new_n943), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n924), .A2(new_n925), .A3(new_n916), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT41), .B1(new_n927), .B2(new_n928), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n988), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n987), .A2(KEYINPUT105), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n965), .B(new_n914), .C1(new_n986), .C2(new_n967), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(new_n952), .A3(new_n973), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n943), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n991), .B1(new_n998), .B2(G37), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n989), .A2(new_n943), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n990), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n1003));
  AOI21_X1  g578(.A(G37), .B1(new_n989), .B2(new_n943), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n993), .A2(KEYINPUT107), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n993), .A2(KEYINPUT107), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n929), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n972), .A2(new_n973), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1007), .A2(new_n1008), .B1(new_n987), .B2(new_n974), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1003), .B(new_n1004), .C1(new_n1009), .C2(new_n943), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1002), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n990), .A2(new_n999), .A3(new_n1003), .A4(new_n1000), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(KEYINPUT108), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1004), .B1(new_n1009), .B2(new_n943), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1012), .B1(new_n1016), .B2(KEYINPUT43), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(KEYINPUT108), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1013), .B1(new_n1015), .B2(new_n1019), .ZN(G397));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n891), .A2(new_n1021), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1022), .A2(KEYINPUT109), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n1022), .B2(KEYINPUT109), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n469), .A2(G40), .A3(new_n475), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n822), .B(new_n824), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n763), .B2(new_n1031), .ZN(new_n1032));
  OR3_X1    g607(.A1(new_n1030), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT46), .B1(new_n1030), .B2(G1996), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT47), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1037));
  XOR2_X1   g612(.A(new_n1037), .B(KEYINPUT111), .Z(new_n1038));
  INV_X1    g613(.A(new_n1030), .ZN(new_n1039));
  XOR2_X1   g614(.A(new_n763), .B(G1996), .Z(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n875), .A2(new_n744), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n885), .A2(new_n824), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1030), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n875), .A2(new_n744), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1039), .B1(new_n1046), .B2(new_n1042), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1030), .A2(G1986), .A3(G290), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  AOI211_X1 g626(.A(new_n1036), .B(new_n1045), .C1(new_n1048), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n561), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(KEYINPUT117), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n920), .A2(new_n1056), .A3(new_n562), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n569), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(KEYINPUT118), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1059), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1065), .B1(new_n1067), .B2(new_n1062), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n469), .A2(G40), .A3(new_n475), .ZN(new_n1069));
  AOI21_X1  g644(.A(G1384), .B1(new_n887), .B2(new_n890), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(KEYINPUT45), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT50), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1069), .B1(new_n1070), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1077), .B2(new_n1070), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n843), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1064), .A2(new_n1068), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1070), .B2(new_n1077), .ZN(new_n1084));
  OAI211_X1 g659(.A(KEYINPUT112), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n1078), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1086), .B2(new_n1078), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1088), .A2(new_n1089), .A3(G1348), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1022), .A2(new_n1069), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(G2067), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n621), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(KEYINPUT120), .B(new_n621), .C1(new_n1090), .C2(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1081), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1082), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1064), .A2(new_n1068), .A3(new_n1081), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(new_n1099), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1089), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1086), .A2(new_n1087), .A3(new_n1078), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n830), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1093), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n612), .A2(KEYINPUT60), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT58), .B(G1341), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1073), .A2(G1996), .B1(new_n1091), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n553), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1111), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1108), .A2(new_n612), .A3(new_n1109), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1094), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1119), .B2(KEYINPUT60), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1081), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT118), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1067), .A2(new_n1065), .A3(new_n1062), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(KEYINPUT61), .A3(new_n1082), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1105), .A2(new_n1120), .A3(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(KEYINPUT121), .B(new_n1082), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1102), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n1074), .B2(new_n788), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(new_n836), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1029), .B1(new_n1070), .B2(KEYINPUT45), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1070), .A2(KEYINPUT114), .A3(new_n1025), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1132), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(KEYINPUT53), .A3(new_n788), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1131), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT54), .B1(new_n1138), .B2(new_n614), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1029), .A2(KEYINPUT53), .A3(new_n788), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT45), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1027), .B(new_n1140), .C1(new_n1141), .C2(new_n1022), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n983), .B1(new_n1131), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1138), .A2(new_n614), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1131), .A2(G301), .A3(new_n1142), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT54), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1086), .A2(new_n777), .A3(new_n1078), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1136), .B2(G1966), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G8), .ZN(new_n1150));
  NAND2_X1  g725(.A1(G286), .A2(G8), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(G8), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1069), .B1(new_n1022), .B2(new_n1141), .ZN(new_n1156));
  NOR4_X1   g731(.A1(G164), .A2(new_n1133), .A3(G1384), .A4(new_n1024), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT114), .B1(new_n1070), .B2(new_n1025), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n805), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1155), .B1(new_n1160), .B2(new_n1148), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(G286), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1163), .A2(KEYINPUT51), .ZN(new_n1164));
  OAI211_X1 g739(.A(G8), .B(new_n1164), .C1(new_n1149), .C2(G286), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1154), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT113), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(KEYINPUT49), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n594), .A2(G1981), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n594), .A2(G1981), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1168), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1171), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1168), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1173), .A2(new_n1169), .A3(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1091), .A2(new_n1155), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1172), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1086), .A2(new_n1078), .ZN(new_n1178));
  OAI22_X1  g753(.A1(new_n1178), .A2(G2090), .B1(new_n1074), .B2(G1971), .ZN(new_n1179));
  NAND3_X1  g754(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT55), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(G166), .B2(new_n1155), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1179), .A2(new_n1183), .A3(G8), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT52), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n581), .B(G1976), .C1(new_n585), .C2(new_n586), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1185), .B1(new_n1176), .B2(new_n1186), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1176), .A2(new_n1186), .ZN(new_n1188));
  INV_X1    g763(.A(G1976), .ZN(new_n1189));
  AOI21_X1  g764(.A(KEYINPUT52), .B1(G288), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1187), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1177), .A2(new_n1184), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1183), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1079), .A2(G2090), .ZN(new_n1194));
  AOI21_X1  g769(.A(G1971), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1195));
  OAI21_X1  g770(.A(G8), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1166), .A2(new_n1192), .A3(new_n1197), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1144), .A2(new_n1147), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1128), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1166), .A2(KEYINPUT62), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(KEYINPUT123), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1166), .A2(new_n1203), .A3(KEYINPUT62), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1197), .A2(new_n1177), .A3(new_n1184), .A4(new_n1191), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1145), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1154), .A2(new_n1207), .A3(new_n1162), .A4(new_n1165), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1202), .A2(new_n1204), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n716), .A2(new_n1189), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1171), .B1(new_n1177), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1176), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1177), .A2(new_n1191), .ZN(new_n1214));
  OAI22_X1  g789(.A1(new_n1212), .A2(new_n1213), .B1(new_n1214), .B2(new_n1184), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT63), .ZN(new_n1216));
  AND4_X1   g791(.A1(KEYINPUT115), .A2(new_n1149), .A3(G8), .A4(G168), .ZN(new_n1217));
  AOI21_X1  g792(.A(KEYINPUT115), .B1(new_n1161), .B2(G168), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1216), .B1(new_n1219), .B2(new_n1205), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1179), .A2(G8), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1216), .B1(new_n1221), .B2(new_n1193), .ZN(new_n1222));
  OAI211_X1 g797(.A(new_n1192), .B(new_n1222), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1215), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1209), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g800(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1200), .A2(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n603), .B(new_n748), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1039), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1048), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g805(.A(new_n1230), .ZN(new_n1231));
  AOI21_X1  g806(.A(KEYINPUT124), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1225), .B1(new_n1128), .B2(new_n1199), .ZN(new_n1233));
  INV_X1    g808(.A(KEYINPUT124), .ZN(new_n1234));
  NOR3_X1   g809(.A1(new_n1233), .A2(new_n1234), .A3(new_n1230), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1052), .B1(new_n1232), .B2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g811(.A(KEYINPUT127), .ZN(new_n1238));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n1239));
  NOR2_X1   g813(.A1(G227), .A2(new_n464), .ZN(new_n1240));
  AND3_X1   g814(.A1(new_n670), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g815(.A(new_n1239), .B1(new_n670), .B2(new_n1240), .ZN(new_n1242));
  OAI211_X1 g816(.A(new_n705), .B(new_n912), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1243));
  INV_X1    g817(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g818(.A(new_n1238), .B1(new_n1011), .B2(new_n1244), .ZN(new_n1245));
  AOI211_X1 g819(.A(KEYINPUT127), .B(new_n1243), .C1(new_n1002), .C2(new_n1010), .ZN(new_n1246));
  NOR2_X1   g820(.A1(new_n1245), .A2(new_n1246), .ZN(G308));
  NAND2_X1  g821(.A1(new_n1011), .A2(new_n1244), .ZN(G225));
endmodule


