

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n545), .A2(n544), .ZN(G160) );
  BUF_X1 U553 ( .A(n582), .Z(n538) );
  BUF_X1 U554 ( .A(n705), .Z(n706) );
  NOR2_X1 U555 ( .A1(G168), .A2(n597), .ZN(n599) );
  XNOR2_X1 U556 ( .A(n537), .B(n536), .ZN(n582) );
  XNOR2_X1 U557 ( .A(n535), .B(KEYINPUT70), .ZN(n536) );
  NOR2_X1 U558 ( .A1(n660), .A2(n664), .ZN(n595) );
  INV_X1 U559 ( .A(KEYINPUT94), .ZN(n598) );
  INV_X1 U560 ( .A(KEYINPUT96), .ZN(n659) );
  XNOR2_X1 U561 ( .A(n667), .B(n659), .ZN(n661) );
  INV_X1 U562 ( .A(KEYINPUT97), .ZN(n662) );
  NOR2_X1 U563 ( .A1(G1384), .A2(G164), .ZN(n590) );
  INV_X1 U564 ( .A(KEYINPUT17), .ZN(n535) );
  XOR2_X1 U565 ( .A(KEYINPUT66), .B(G2104), .Z(n541) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n790) );
  XNOR2_X1 U567 ( .A(n542), .B(KEYINPUT67), .ZN(n705) );
  NOR2_X1 U568 ( .A1(G651), .A2(n571), .ZN(n787) );
  XOR2_X1 U569 ( .A(KEYINPUT0), .B(G543), .Z(n571) );
  INV_X1 U570 ( .A(G651), .ZN(n522) );
  NOR2_X1 U571 ( .A1(n571), .A2(n522), .ZN(n791) );
  NAND2_X1 U572 ( .A1(n791), .A2(G76), .ZN(n517) );
  XNOR2_X1 U573 ( .A(KEYINPUT74), .B(n517), .ZN(n520) );
  NAND2_X1 U574 ( .A1(n790), .A2(G89), .ZN(n518) );
  XNOR2_X1 U575 ( .A(KEYINPUT4), .B(n518), .ZN(n519) );
  NAND2_X1 U576 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U577 ( .A(n521), .B(KEYINPUT5), .ZN(n528) );
  NOR2_X1 U578 ( .A1(G543), .A2(n522), .ZN(n523) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n523), .Z(n786) );
  NAND2_X1 U580 ( .A1(G63), .A2(n786), .ZN(n525) );
  NAND2_X1 U581 ( .A1(G51), .A2(n787), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U583 ( .A(KEYINPUT6), .B(n526), .Z(n527) );
  NAND2_X1 U584 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U585 ( .A(n529), .B(KEYINPUT7), .ZN(G168) );
  AND2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n852) );
  NAND2_X1 U587 ( .A1(G113), .A2(n852), .ZN(n530) );
  XNOR2_X1 U588 ( .A(n530), .B(KEYINPUT69), .ZN(n534) );
  INV_X1 U589 ( .A(n541), .ZN(n581) );
  INV_X1 U590 ( .A(G2105), .ZN(n580) );
  AND2_X1 U591 ( .A1(G101), .A2(n580), .ZN(n531) );
  NAND2_X1 U592 ( .A1(n581), .A2(n531), .ZN(n532) );
  XNOR2_X1 U593 ( .A(KEYINPUT23), .B(n532), .ZN(n533) );
  NOR2_X1 U594 ( .A1(n534), .A2(n533), .ZN(n540) );
  NOR2_X1 U595 ( .A1(G2104), .A2(G2105), .ZN(n537) );
  NAND2_X1 U596 ( .A1(G137), .A2(n538), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G2105), .A2(n541), .ZN(n542) );
  NAND2_X1 U599 ( .A1(G125), .A2(n705), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT68), .B(n543), .Z(n544) );
  NAND2_X1 U601 ( .A1(G61), .A2(n786), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G86), .A2(n790), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n791), .A2(G73), .ZN(n548) );
  XOR2_X1 U605 ( .A(KEYINPUT2), .B(n548), .Z(n549) );
  NOR2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n787), .A2(G48), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(G305) );
  NAND2_X1 U609 ( .A1(n790), .A2(G90), .ZN(n553) );
  XNOR2_X1 U610 ( .A(n553), .B(KEYINPUT72), .ZN(n555) );
  NAND2_X1 U611 ( .A1(G77), .A2(n791), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U613 ( .A(n556), .B(KEYINPUT9), .ZN(n558) );
  NAND2_X1 U614 ( .A1(G64), .A2(n786), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G52), .A2(n787), .ZN(n559) );
  XNOR2_X1 U617 ( .A(KEYINPUT71), .B(n559), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n561), .A2(n560), .ZN(G171) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U620 ( .A1(G88), .A2(n790), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G75), .A2(n791), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U623 ( .A1(G62), .A2(n786), .ZN(n565) );
  NAND2_X1 U624 ( .A1(G50), .A2(n787), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U626 ( .A1(n567), .A2(n566), .ZN(G166) );
  INV_X1 U627 ( .A(G166), .ZN(G303) );
  NAND2_X1 U628 ( .A1(G49), .A2(n787), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G74), .A2(G651), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U631 ( .A1(n786), .A2(n570), .ZN(n573) );
  NAND2_X1 U632 ( .A1(n571), .A2(G87), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n573), .A2(n572), .ZN(G288) );
  NAND2_X1 U634 ( .A1(G85), .A2(n790), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G72), .A2(n791), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U637 ( .A1(G60), .A2(n786), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G47), .A2(n787), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n578) );
  OR2_X1 U640 ( .A1(n579), .A2(n578), .ZN(G290) );
  INV_X1 U641 ( .A(G8), .ZN(n592) );
  AND2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n858) );
  NAND2_X1 U643 ( .A1(n858), .A2(G102), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n582), .A2(G138), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT83), .B(n583), .Z(n584) );
  NAND2_X1 U646 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U647 ( .A1(G114), .A2(n852), .ZN(n587) );
  NAND2_X1 U648 ( .A1(G126), .A2(n705), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U650 ( .A1(n589), .A2(n588), .ZN(G164) );
  XNOR2_X1 U651 ( .A(n590), .B(KEYINPUT64), .ZN(n591) );
  INV_X1 U652 ( .A(n591), .ZN(n725) );
  NAND2_X1 U653 ( .A1(G160), .A2(G40), .ZN(n726) );
  NOR2_X4 U654 ( .A1(n725), .A2(n726), .ZN(n642) );
  OR2_X2 U655 ( .A1(n592), .A2(n642), .ZN(n698) );
  NOR2_X1 U656 ( .A1(G1981), .A2(G305), .ZN(n593) );
  XOR2_X1 U657 ( .A(n593), .B(KEYINPUT24), .Z(n594) );
  NOR2_X1 U658 ( .A1(n698), .A2(n594), .ZN(n704) );
  NOR2_X1 U659 ( .A1(G1966), .A2(n698), .ZN(n660) );
  INV_X1 U660 ( .A(n642), .ZN(n668) );
  NOR2_X1 U661 ( .A1(G2084), .A2(n668), .ZN(n664) );
  NAND2_X1 U662 ( .A1(n595), .A2(G8), .ZN(n596) );
  XNOR2_X1 U663 ( .A(n596), .B(KEYINPUT30), .ZN(n597) );
  XNOR2_X1 U664 ( .A(n599), .B(n598), .ZN(n605) );
  XOR2_X1 U665 ( .A(G2078), .B(KEYINPUT25), .Z(n1005) );
  NOR2_X1 U666 ( .A1(n668), .A2(n1005), .ZN(n601) );
  NOR2_X1 U667 ( .A1(n642), .A2(G1961), .ZN(n600) );
  NOR2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U669 ( .A(KEYINPUT91), .B(n602), .ZN(n607) );
  NOR2_X1 U670 ( .A1(G171), .A2(n607), .ZN(n603) );
  XNOR2_X1 U671 ( .A(KEYINPUT95), .B(n603), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U673 ( .A(n606), .B(KEYINPUT31), .ZN(n658) );
  NAND2_X1 U674 ( .A1(n607), .A2(G171), .ZN(n656) );
  NAND2_X1 U675 ( .A1(G65), .A2(n786), .ZN(n609) );
  NAND2_X1 U676 ( .A1(G53), .A2(n787), .ZN(n608) );
  NAND2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U678 ( .A1(G91), .A2(n790), .ZN(n611) );
  NAND2_X1 U679 ( .A1(G78), .A2(n791), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U681 ( .A1(n613), .A2(n612), .ZN(n917) );
  NAND2_X1 U682 ( .A1(n642), .A2(G2072), .ZN(n614) );
  XNOR2_X1 U683 ( .A(n614), .B(KEYINPUT27), .ZN(n616) );
  INV_X1 U684 ( .A(G1956), .ZN(n975) );
  NOR2_X1 U685 ( .A1(n975), .A2(n642), .ZN(n615) );
  NOR2_X1 U686 ( .A1(n616), .A2(n615), .ZN(n619) );
  NOR2_X1 U687 ( .A1(n917), .A2(n619), .ZN(n618) );
  XOR2_X1 U688 ( .A(KEYINPUT92), .B(KEYINPUT28), .Z(n617) );
  XNOR2_X1 U689 ( .A(n618), .B(n617), .ZN(n653) );
  NAND2_X1 U690 ( .A1(n917), .A2(n619), .ZN(n651) );
  NAND2_X1 U691 ( .A1(G56), .A2(n786), .ZN(n620) );
  XOR2_X1 U692 ( .A(KEYINPUT14), .B(n620), .Z(n626) );
  NAND2_X1 U693 ( .A1(n790), .A2(G81), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n621), .B(KEYINPUT12), .ZN(n623) );
  NAND2_X1 U695 ( .A1(G68), .A2(n791), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U697 ( .A(KEYINPUT13), .B(n624), .Z(n625) );
  NOR2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U699 ( .A1(n787), .A2(G43), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n949) );
  NAND2_X1 U701 ( .A1(n642), .A2(G1996), .ZN(n630) );
  XOR2_X1 U702 ( .A(KEYINPUT26), .B(KEYINPUT93), .Z(n629) );
  XNOR2_X1 U703 ( .A(n630), .B(n629), .ZN(n632) );
  NAND2_X1 U704 ( .A1(n668), .A2(G1341), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U706 ( .A1(n949), .A2(n633), .ZN(n634) );
  XNOR2_X1 U707 ( .A(KEYINPUT65), .B(n634), .ZN(n646) );
  NAND2_X1 U708 ( .A1(G66), .A2(n786), .ZN(n636) );
  NAND2_X1 U709 ( .A1(G92), .A2(n790), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U711 ( .A1(G79), .A2(n791), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G54), .A2(n787), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U715 ( .A(KEYINPUT15), .B(n641), .Z(n952) );
  INV_X1 U716 ( .A(n952), .ZN(n761) );
  NAND2_X1 U717 ( .A1(G2067), .A2(n642), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G1348), .A2(n668), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n647) );
  OR2_X1 U720 ( .A1(n761), .A2(n647), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n761), .A2(n647), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U726 ( .A(KEYINPUT29), .B(n654), .Z(n655) );
  NAND2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n667) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U730 ( .A(n663), .B(n662), .ZN(n666) );
  NAND2_X1 U731 ( .A1(G8), .A2(n664), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n677) );
  NAND2_X1 U733 ( .A1(G286), .A2(n667), .ZN(n673) );
  NOR2_X1 U734 ( .A1(G1971), .A2(n698), .ZN(n670) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n668), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U737 ( .A1(n671), .A2(G303), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U739 ( .A1(G8), .A2(n674), .ZN(n675) );
  XNOR2_X1 U740 ( .A(KEYINPUT32), .B(n675), .ZN(n676) );
  NAND2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n697) );
  NOR2_X1 U742 ( .A1(G1971), .A2(G303), .ZN(n678) );
  NOR2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n964) );
  NOR2_X1 U744 ( .A1(n678), .A2(n964), .ZN(n680) );
  INV_X1 U745 ( .A(KEYINPUT33), .ZN(n679) );
  AND2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U747 ( .A1(n697), .A2(n681), .ZN(n694) );
  INV_X1 U748 ( .A(n698), .ZN(n682) );
  NAND2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n967) );
  AND2_X1 U750 ( .A1(n682), .A2(n967), .ZN(n683) );
  AND2_X1 U751 ( .A1(n683), .A2(KEYINPUT98), .ZN(n684) );
  NOR2_X1 U752 ( .A1(KEYINPUT33), .A2(n684), .ZN(n691) );
  INV_X1 U753 ( .A(KEYINPUT98), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n685), .A2(n964), .ZN(n688) );
  NAND2_X1 U755 ( .A1(n964), .A2(KEYINPUT33), .ZN(n686) );
  NAND2_X1 U756 ( .A1(n686), .A2(KEYINPUT98), .ZN(n687) );
  NAND2_X1 U757 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U758 ( .A1(n698), .A2(n689), .ZN(n690) );
  NOR2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n957) );
  AND2_X1 U761 ( .A1(n692), .A2(n957), .ZN(n693) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n701) );
  NOR2_X1 U763 ( .A1(G2090), .A2(G303), .ZN(n695) );
  NAND2_X1 U764 ( .A1(G8), .A2(n695), .ZN(n696) );
  NAND2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U768 ( .A(KEYINPUT99), .B(n702), .Z(n703) );
  NOR2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n740) );
  XNOR2_X1 U770 ( .A(KEYINPUT88), .B(G1991), .ZN(n1004) );
  NAND2_X1 U771 ( .A1(G107), .A2(n852), .ZN(n708) );
  NAND2_X1 U772 ( .A1(G119), .A2(n706), .ZN(n707) );
  NAND2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U774 ( .A(KEYINPUT86), .B(n709), .ZN(n712) );
  NAND2_X1 U775 ( .A1(G95), .A2(n858), .ZN(n710) );
  XNOR2_X1 U776 ( .A(KEYINPUT87), .B(n710), .ZN(n711) );
  NOR2_X1 U777 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U778 ( .A1(G131), .A2(n538), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n714), .A2(n713), .ZN(n866) );
  AND2_X1 U780 ( .A1(n1004), .A2(n866), .ZN(n724) );
  NAND2_X1 U781 ( .A1(G105), .A2(n858), .ZN(n715) );
  XNOR2_X1 U782 ( .A(n715), .B(KEYINPUT38), .ZN(n722) );
  NAND2_X1 U783 ( .A1(n706), .A2(G129), .ZN(n717) );
  NAND2_X1 U784 ( .A1(G141), .A2(n538), .ZN(n716) );
  NAND2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U786 ( .A1(G117), .A2(n852), .ZN(n718) );
  XNOR2_X1 U787 ( .A(KEYINPUT89), .B(n718), .ZN(n719) );
  NOR2_X1 U788 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U789 ( .A1(n722), .A2(n721), .ZN(n851) );
  AND2_X1 U790 ( .A1(n851), .A2(G1996), .ZN(n723) );
  OR2_X1 U791 ( .A1(n724), .A2(n723), .ZN(n922) );
  NOR2_X1 U792 ( .A1(n726), .A2(n591), .ZN(n752) );
  AND2_X1 U793 ( .A1(n922), .A2(n752), .ZN(n745) );
  XOR2_X1 U794 ( .A(KEYINPUT90), .B(n745), .Z(n738) );
  XNOR2_X1 U795 ( .A(KEYINPUT37), .B(G2067), .ZN(n750) );
  XNOR2_X1 U796 ( .A(KEYINPUT35), .B(KEYINPUT85), .ZN(n730) );
  NAND2_X1 U797 ( .A1(G116), .A2(n852), .ZN(n728) );
  NAND2_X1 U798 ( .A1(G128), .A2(n706), .ZN(n727) );
  NAND2_X1 U799 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U800 ( .A(n730), .B(n729), .ZN(n736) );
  NAND2_X1 U801 ( .A1(n858), .A2(G104), .ZN(n731) );
  XNOR2_X1 U802 ( .A(n731), .B(KEYINPUT84), .ZN(n733) );
  NAND2_X1 U803 ( .A1(G140), .A2(n538), .ZN(n732) );
  NAND2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U805 ( .A(KEYINPUT34), .B(n734), .ZN(n735) );
  NOR2_X1 U806 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U807 ( .A(KEYINPUT36), .B(n737), .ZN(n871) );
  NOR2_X1 U808 ( .A1(n750), .A2(n871), .ZN(n923) );
  NAND2_X1 U809 ( .A1(n752), .A2(n923), .ZN(n748) );
  NAND2_X1 U810 ( .A1(n738), .A2(n748), .ZN(n739) );
  NOR2_X1 U811 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X1 U812 ( .A(G1986), .B(G290), .ZN(n954) );
  NAND2_X1 U813 ( .A1(n954), .A2(n752), .ZN(n741) );
  NAND2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n755) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n851), .ZN(n919) );
  NOR2_X1 U816 ( .A1(n1004), .A2(n866), .ZN(n928) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n743) );
  NOR2_X1 U818 ( .A1(n928), .A2(n743), .ZN(n744) );
  NOR2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n919), .A2(n746), .ZN(n747) );
  XNOR2_X1 U821 ( .A(n747), .B(KEYINPUT39), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n749), .A2(n748), .ZN(n751) );
  NAND2_X1 U823 ( .A1(n750), .A2(n871), .ZN(n933) );
  NAND2_X1 U824 ( .A1(n751), .A2(n933), .ZN(n753) );
  NAND2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U827 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U828 ( .A(G57), .ZN(G237) );
  INV_X1 U829 ( .A(G132), .ZN(G219) );
  INV_X1 U830 ( .A(G82), .ZN(G220) );
  NAND2_X1 U831 ( .A1(G94), .A2(G452), .ZN(n758) );
  XNOR2_X1 U832 ( .A(n758), .B(KEYINPUT73), .ZN(G173) );
  NAND2_X1 U833 ( .A1(G7), .A2(G661), .ZN(n759) );
  XNOR2_X1 U834 ( .A(n759), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U835 ( .A(G223), .ZN(n825) );
  NAND2_X1 U836 ( .A1(n825), .A2(G567), .ZN(n760) );
  XOR2_X1 U837 ( .A(KEYINPUT11), .B(n760), .Z(G234) );
  INV_X1 U838 ( .A(G860), .ZN(n767) );
  OR2_X1 U839 ( .A1(n949), .A2(n767), .ZN(G153) );
  INV_X1 U840 ( .A(G171), .ZN(G301) );
  NAND2_X1 U841 ( .A1(G868), .A2(G301), .ZN(n763) );
  INV_X1 U842 ( .A(G868), .ZN(n806) );
  NAND2_X1 U843 ( .A1(n761), .A2(n806), .ZN(n762) );
  NAND2_X1 U844 ( .A1(n763), .A2(n762), .ZN(G284) );
  NAND2_X1 U845 ( .A1(n917), .A2(n806), .ZN(n764) );
  XNOR2_X1 U846 ( .A(n764), .B(KEYINPUT75), .ZN(n766) );
  NOR2_X1 U847 ( .A1(n806), .A2(G286), .ZN(n765) );
  NOR2_X1 U848 ( .A1(n766), .A2(n765), .ZN(G297) );
  NAND2_X1 U849 ( .A1(n767), .A2(G559), .ZN(n768) );
  NAND2_X1 U850 ( .A1(n768), .A2(n952), .ZN(n769) );
  XNOR2_X1 U851 ( .A(n769), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U852 ( .A1(G868), .A2(n949), .ZN(n772) );
  NAND2_X1 U853 ( .A1(G868), .A2(n952), .ZN(n770) );
  NOR2_X1 U854 ( .A1(G559), .A2(n770), .ZN(n771) );
  NOR2_X1 U855 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U856 ( .A(KEYINPUT76), .B(n773), .ZN(G282) );
  NAND2_X1 U857 ( .A1(n858), .A2(G99), .ZN(n775) );
  NAND2_X1 U858 ( .A1(G135), .A2(n538), .ZN(n774) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n782) );
  NAND2_X1 U860 ( .A1(G111), .A2(n852), .ZN(n776) );
  XNOR2_X1 U861 ( .A(n776), .B(KEYINPUT78), .ZN(n780) );
  XOR2_X1 U862 ( .A(KEYINPUT18), .B(KEYINPUT77), .Z(n778) );
  NAND2_X1 U863 ( .A1(G123), .A2(n706), .ZN(n777) );
  XNOR2_X1 U864 ( .A(n778), .B(n777), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U866 ( .A1(n782), .A2(n781), .ZN(n927) );
  XNOR2_X1 U867 ( .A(G2096), .B(n927), .ZN(n784) );
  INV_X1 U868 ( .A(G2100), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(G156) );
  NAND2_X1 U870 ( .A1(n952), .A2(G559), .ZN(n804) );
  XNOR2_X1 U871 ( .A(n949), .B(n804), .ZN(n785) );
  NOR2_X1 U872 ( .A1(n785), .A2(G860), .ZN(n796) );
  NAND2_X1 U873 ( .A1(G67), .A2(n786), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G55), .A2(n787), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n795) );
  NAND2_X1 U876 ( .A1(G93), .A2(n790), .ZN(n793) );
  NAND2_X1 U877 ( .A1(G80), .A2(n791), .ZN(n792) );
  NAND2_X1 U878 ( .A1(n793), .A2(n792), .ZN(n794) );
  OR2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n807) );
  XOR2_X1 U880 ( .A(n796), .B(n807), .Z(G145) );
  XNOR2_X1 U881 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n798) );
  XNOR2_X1 U882 ( .A(G305), .B(G166), .ZN(n797) );
  XNOR2_X1 U883 ( .A(n798), .B(n797), .ZN(n801) );
  XNOR2_X1 U884 ( .A(n917), .B(n949), .ZN(n799) );
  XNOR2_X1 U885 ( .A(n799), .B(G288), .ZN(n800) );
  XNOR2_X1 U886 ( .A(n801), .B(n800), .ZN(n803) );
  XOR2_X1 U887 ( .A(G290), .B(n807), .Z(n802) );
  XNOR2_X1 U888 ( .A(n803), .B(n802), .ZN(n877) );
  XOR2_X1 U889 ( .A(n877), .B(n804), .Z(n805) );
  NAND2_X1 U890 ( .A1(G868), .A2(n805), .ZN(n809) );
  NAND2_X1 U891 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U892 ( .A1(n809), .A2(n808), .ZN(G295) );
  NAND2_X1 U893 ( .A1(G2084), .A2(G2078), .ZN(n811) );
  XOR2_X1 U894 ( .A(KEYINPUT80), .B(KEYINPUT20), .Z(n810) );
  XNOR2_X1 U895 ( .A(n811), .B(n810), .ZN(n812) );
  NAND2_X1 U896 ( .A1(n812), .A2(G2090), .ZN(n813) );
  XOR2_X1 U897 ( .A(KEYINPUT81), .B(n813), .Z(n814) );
  XNOR2_X1 U898 ( .A(KEYINPUT21), .B(n814), .ZN(n815) );
  NAND2_X1 U899 ( .A1(n815), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U900 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U901 ( .A1(G220), .A2(G219), .ZN(n816) );
  XOR2_X1 U902 ( .A(KEYINPUT22), .B(n816), .Z(n817) );
  NOR2_X1 U903 ( .A1(G218), .A2(n817), .ZN(n818) );
  XNOR2_X1 U904 ( .A(KEYINPUT82), .B(n818), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n819), .A2(G96), .ZN(n831) );
  NAND2_X1 U906 ( .A1(n831), .A2(G2106), .ZN(n823) );
  NAND2_X1 U907 ( .A1(G120), .A2(G69), .ZN(n820) );
  NOR2_X1 U908 ( .A1(G237), .A2(n820), .ZN(n821) );
  NAND2_X1 U909 ( .A1(G108), .A2(n821), .ZN(n832) );
  NAND2_X1 U910 ( .A1(n832), .A2(G567), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n823), .A2(n822), .ZN(n889) );
  NAND2_X1 U912 ( .A1(G661), .A2(G483), .ZN(n824) );
  NOR2_X1 U913 ( .A1(n889), .A2(n824), .ZN(n829) );
  NAND2_X1 U914 ( .A1(n829), .A2(G36), .ZN(G176) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n825), .ZN(G217) );
  NAND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n826) );
  XNOR2_X1 U917 ( .A(KEYINPUT101), .B(n826), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n827), .A2(G661), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n828) );
  XNOR2_X1 U920 ( .A(KEYINPUT102), .B(n828), .ZN(n830) );
  NAND2_X1 U921 ( .A1(n830), .A2(n829), .ZN(G188) );
  XNOR2_X1 U922 ( .A(G69), .B(KEYINPUT103), .ZN(G235) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  NOR2_X1 U926 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  NAND2_X1 U928 ( .A1(n706), .A2(G124), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n833), .B(KEYINPUT44), .ZN(n835) );
  NAND2_X1 U930 ( .A1(G136), .A2(n538), .ZN(n834) );
  NAND2_X1 U931 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U932 ( .A(KEYINPUT106), .B(n836), .ZN(n840) );
  NAND2_X1 U933 ( .A1(G112), .A2(n852), .ZN(n838) );
  NAND2_X1 U934 ( .A1(G100), .A2(n858), .ZN(n837) );
  NAND2_X1 U935 ( .A1(n838), .A2(n837), .ZN(n839) );
  NOR2_X1 U936 ( .A1(n840), .A2(n839), .ZN(G162) );
  NAND2_X1 U937 ( .A1(n858), .A2(G106), .ZN(n842) );
  NAND2_X1 U938 ( .A1(G142), .A2(n538), .ZN(n841) );
  NAND2_X1 U939 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n843), .B(KEYINPUT45), .ZN(n848) );
  NAND2_X1 U941 ( .A1(G118), .A2(n852), .ZN(n845) );
  NAND2_X1 U942 ( .A1(G130), .A2(n706), .ZN(n844) );
  NAND2_X1 U943 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U944 ( .A(KEYINPUT107), .B(n846), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n849), .B(n927), .ZN(n850) );
  XOR2_X1 U947 ( .A(n851), .B(n850), .Z(n870) );
  XOR2_X1 U948 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n864) );
  XNOR2_X1 U949 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n857) );
  NAND2_X1 U950 ( .A1(G115), .A2(n852), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G127), .A2(n706), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n855), .B(KEYINPUT47), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n862) );
  NAND2_X1 U955 ( .A1(n858), .A2(G103), .ZN(n860) );
  NAND2_X1 U956 ( .A1(G139), .A2(n538), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U958 ( .A1(n862), .A2(n861), .ZN(n938) );
  XNOR2_X1 U959 ( .A(G164), .B(n938), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U961 ( .A(n865), .B(G162), .Z(n868) );
  XOR2_X1 U962 ( .A(G160), .B(n866), .Z(n867) );
  XNOR2_X1 U963 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U964 ( .A(n870), .B(n869), .ZN(n872) );
  XOR2_X1 U965 ( .A(n872), .B(n871), .Z(n873) );
  NOR2_X1 U966 ( .A1(G37), .A2(n873), .ZN(G395) );
  XOR2_X1 U967 ( .A(KEYINPUT110), .B(G286), .Z(n875) );
  XNOR2_X1 U968 ( .A(G171), .B(n952), .ZN(n874) );
  XNOR2_X1 U969 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U970 ( .A(n877), .B(n876), .Z(n878) );
  NOR2_X1 U971 ( .A1(G37), .A2(n878), .ZN(G397) );
  XNOR2_X1 U972 ( .A(G1341), .B(G2454), .ZN(n879) );
  XNOR2_X1 U973 ( .A(n879), .B(G2430), .ZN(n880) );
  XNOR2_X1 U974 ( .A(n880), .B(G1348), .ZN(n886) );
  XOR2_X1 U975 ( .A(G2443), .B(G2427), .Z(n882) );
  XNOR2_X1 U976 ( .A(G2438), .B(G2446), .ZN(n881) );
  XNOR2_X1 U977 ( .A(n882), .B(n881), .ZN(n884) );
  XOR2_X1 U978 ( .A(G2451), .B(G2435), .Z(n883) );
  XNOR2_X1 U979 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U980 ( .A(n886), .B(n885), .ZN(n887) );
  NAND2_X1 U981 ( .A1(n887), .A2(G14), .ZN(n888) );
  XOR2_X1 U982 ( .A(KEYINPUT100), .B(n888), .Z(G401) );
  INV_X1 U983 ( .A(n889), .ZN(G319) );
  XOR2_X1 U984 ( .A(G2096), .B(KEYINPUT104), .Z(n891) );
  XNOR2_X1 U985 ( .A(G2090), .B(KEYINPUT43), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U987 ( .A(n892), .B(KEYINPUT42), .Z(n894) );
  XNOR2_X1 U988 ( .A(G2067), .B(G2072), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n898) );
  XOR2_X1 U990 ( .A(G2678), .B(G2100), .Z(n896) );
  XNOR2_X1 U991 ( .A(G2084), .B(G2078), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(G227) );
  XOR2_X1 U994 ( .A(G1976), .B(G1966), .Z(n900) );
  XNOR2_X1 U995 ( .A(G1986), .B(G1981), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U997 ( .A(G1971), .B(G1956), .Z(n902) );
  XNOR2_X1 U998 ( .A(G1996), .B(G1991), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1001 ( .A(KEYINPUT105), .B(G2474), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1003 ( .A(G1961), .B(KEYINPUT41), .Z(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(G229) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n909) );
  XOR2_X1 U1006 ( .A(KEYINPUT113), .B(n909), .Z(n916) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(KEYINPUT111), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n912), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT112), .B(n914), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(n917), .ZN(G299) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1017 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(KEYINPUT117), .B(n920), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n921), .B(KEYINPUT51), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n936) );
  XOR2_X1 U1023 ( .A(G160), .B(G2084), .Z(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT114), .B(n926), .ZN(n931) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n929), .B(KEYINPUT115), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(n932), .B(KEYINPUT116), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1031 ( .A(KEYINPUT118), .B(n937), .Z(n944) );
  XNOR2_X1 U1032 ( .A(G2072), .B(n938), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(n939), .B(KEYINPUT119), .ZN(n941) );
  XOR2_X1 U1034 ( .A(G2078), .B(G164), .Z(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1036 ( .A(KEYINPUT50), .B(n942), .Z(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(n945), .B(KEYINPUT121), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(n946), .B(KEYINPUT52), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n947), .B(KEYINPUT120), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n948), .A2(G29), .ZN(n1003) );
  INV_X1 U1042 ( .A(G16), .ZN(n972) );
  XNOR2_X1 U1043 ( .A(G301), .B(G1961), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(n949), .B(G1341), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n963) );
  XNOR2_X1 U1046 ( .A(n952), .B(G1348), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(G1956), .B(G299), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n961) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G168), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1052 ( .A(KEYINPUT57), .B(n959), .Z(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1054 ( .A1(n963), .A2(n962), .ZN(n971) );
  XOR2_X1 U1055 ( .A(n964), .B(KEYINPUT125), .Z(n966) );
  XOR2_X1 U1056 ( .A(G166), .B(G1971), .Z(n965) );
  NOR2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n968) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(KEYINPUT126), .B(n969), .ZN(n970) );
  NOR2_X1 U1060 ( .A1(n971), .A2(n970), .ZN(n996) );
  NOR2_X1 U1061 ( .A1(n972), .A2(n996), .ZN(n973) );
  NAND2_X1 U1062 ( .A1(KEYINPUT56), .A2(n973), .ZN(n974) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n974), .ZN(n1001) );
  XNOR2_X1 U1064 ( .A(G20), .B(n975), .ZN(n979) );
  XNOR2_X1 U1065 ( .A(G1981), .B(G6), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(G19), .B(G1341), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1069 ( .A(KEYINPUT59), .B(G1348), .Z(n980) );
  XNOR2_X1 U1070 ( .A(G4), .B(n980), .ZN(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(KEYINPUT60), .B(n983), .ZN(n987) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G21), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(G5), .B(G1961), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n994) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(G23), .B(G1976), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n991) );
  XOR2_X1 U1080 ( .A(G1986), .B(G24), .Z(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(KEYINPUT58), .B(n992), .ZN(n993) );
  NOR2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n995), .B(KEYINPUT61), .ZN(n998) );
  NOR2_X1 U1085 ( .A1(KEYINPUT56), .A2(n996), .ZN(n997) );
  NOR2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(G16), .A2(n999), .ZN(n1000) );
  NOR2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1027) );
  XNOR2_X1 U1090 ( .A(n1004), .B(G25), .ZN(n1015) );
  XOR2_X1 U1091 ( .A(G2072), .B(G33), .Z(n1010) );
  XNOR2_X1 U1092 ( .A(G1996), .B(G32), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(n1005), .B(G27), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(KEYINPUT122), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G26), .B(G2067), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(KEYINPUT123), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1101 ( .A1(G28), .A2(n1016), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(n1017), .B(KEYINPUT53), .ZN(n1020) );
  XOR2_X1 U1103 ( .A(G2084), .B(G34), .Z(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT54), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(G35), .B(G2090), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(n1023), .B(KEYINPUT124), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(G29), .A2(n1024), .ZN(n1025) );
  XOR2_X1 U1110 ( .A(KEYINPUT55), .B(n1025), .Z(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

