//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(G355));
  NAND2_X1  g0009(.A1(new_n206), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G77), .A2(G244), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G97), .A2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G87), .A2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G50), .A2(G226), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G116), .A2(G270), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G68), .A2(G238), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G58), .A2(G232), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G1), .ZN(new_n225));
  OAI22_X1  g0025(.A1(new_n219), .A2(new_n224), .B1(new_n225), .B2(new_n213), .ZN(new_n226));
  AOI22_X1  g0026(.A1(new_n211), .A2(new_n214), .B1(KEYINPUT1), .B2(new_n226), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n225), .A2(new_n213), .A3(G13), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(G250), .B1(G257), .B2(G264), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n232), .A2(KEYINPUT0), .ZN(new_n233));
  OR2_X1    g0033(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(KEYINPUT0), .ZN(new_n235));
  AND4_X1   g0035(.A1(new_n227), .A2(new_n233), .A3(new_n234), .A4(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G97), .B(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n203), .A2(G50), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n247), .B(new_n253), .ZN(G351));
  XNOR2_X1  g0054(.A(KEYINPUT68), .B(G45), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT67), .A2(G41), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT67), .A2(G41), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(G1), .B(G13), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n225), .B1(G41), .B2(G45), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G222), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G77), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G223), .ZN(new_n273));
  OAI221_X1 g0073(.A(new_n270), .B1(new_n271), .B2(new_n268), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n275));
  AOI211_X1 g0075(.A(new_n261), .B(new_n267), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G179), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n212), .ZN(new_n280));
  INV_X1    g0080(.A(new_n206), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n213), .B1(new_n281), .B2(new_n248), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n213), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G150), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n283), .A2(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n280), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n225), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n280), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(G1), .B2(new_n213), .ZN(new_n292));
  MUX2_X1   g0092(.A(new_n290), .B(new_n292), .S(G50), .Z(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n278), .B(new_n294), .C1(G169), .C2(new_n276), .ZN(new_n295));
  INV_X1    g0095(.A(new_n294), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n296), .A2(KEYINPUT9), .B1(new_n276), .B2(G190), .ZN(new_n297));
  INV_X1    g0097(.A(G200), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n297), .B1(KEYINPUT9), .B2(new_n296), .C1(new_n298), .C2(new_n276), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G97), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n268), .A2(new_n269), .ZN(new_n304));
  INV_X1    g0104(.A(G226), .ZN(new_n305));
  INV_X1    g0105(.A(G232), .ZN(new_n306));
  OAI221_X1 g0106(.A(new_n303), .B1(new_n304), .B2(new_n305), .C1(new_n306), .C2(new_n272), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n275), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n261), .B1(G238), .B2(new_n266), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT13), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n310), .B1(new_n308), .B2(new_n309), .ZN(new_n313));
  OAI21_X1  g0113(.A(G200), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n308), .A2(new_n309), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(G190), .A3(new_n311), .ZN(new_n317));
  INV_X1    g0117(.A(new_n290), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n203), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT70), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n320), .A2(KEYINPUT12), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(KEYINPUT12), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n323), .A2(KEYINPUT71), .B1(KEYINPUT12), .B2(new_n319), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(KEYINPUT71), .B2(new_n323), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n287), .A2(new_n248), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n284), .A2(new_n271), .B1(new_n213), .B2(G68), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n280), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n329), .A2(new_n330), .B1(new_n203), .B2(new_n292), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n314), .A2(new_n317), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT72), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n314), .A2(new_n317), .A3(KEYINPUT72), .A4(new_n332), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n332), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n316), .A2(G179), .A3(new_n311), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n316), .B2(new_n311), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n342), .B(G169), .C1(new_n312), .C2(new_n313), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n338), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n337), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n283), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(new_n318), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n292), .B2(new_n348), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT3), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G33), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT7), .B1(new_n355), .B2(new_n213), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT7), .ZN(new_n357));
  AOI211_X1 g0157(.A(new_n357), .B(G20), .C1(new_n352), .C2(new_n354), .ZN(new_n358));
  OAI21_X1  g0158(.A(G68), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G58), .A2(G68), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n204), .A2(new_n205), .A3(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(G20), .B1(G159), .B2(new_n286), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT16), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n291), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(KEYINPUT16), .A3(new_n362), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT73), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n357), .B1(new_n268), .B2(G20), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n355), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n203), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n361), .A2(G20), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n286), .A2(G159), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n364), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n366), .A2(new_n374), .A3(KEYINPUT73), .A4(new_n280), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n351), .B1(new_n367), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n266), .A2(G232), .B1(new_n258), .B2(new_n260), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n352), .A2(new_n354), .A3(G226), .A4(G1698), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n352), .A2(new_n354), .A3(G223), .A4(new_n269), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n275), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n340), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT75), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n382), .A2(KEYINPUT74), .A3(new_n275), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT74), .B1(new_n382), .B2(new_n275), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n258), .A2(new_n260), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n264), .A2(G232), .A3(new_n265), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n277), .A3(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n385), .B(new_n386), .C1(new_n389), .C2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT74), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n383), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n382), .A2(KEYINPUT74), .A3(new_n275), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(G169), .B1(new_n378), .B2(new_n383), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT75), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT18), .B1(new_n377), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n366), .A2(new_n374), .A3(new_n280), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT73), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n350), .B1(new_n404), .B2(new_n375), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n393), .A2(new_n399), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT18), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n404), .A2(new_n375), .ZN(new_n410));
  INV_X1    g0210(.A(G190), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(new_n378), .C1(new_n387), .C2(new_n388), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n384), .A2(new_n298), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND4_X1   g0214(.A1(new_n409), .A2(new_n410), .A3(new_n351), .A4(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n409), .B1(new_n405), .B2(new_n414), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n401), .A2(new_n408), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n318), .A2(new_n271), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n292), .B2(new_n271), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n283), .A2(new_n287), .B1(new_n213), .B2(new_n271), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT15), .B(G87), .Z(new_n421));
  INV_X1    g0221(.A(new_n284), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n420), .B1(KEYINPUT69), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(KEYINPUT69), .B2(new_n423), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n419), .B1(new_n425), .B2(new_n280), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n261), .B1(G244), .B2(new_n266), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n268), .A2(G238), .A3(G1698), .ZN(new_n428));
  INV_X1    g0228(.A(G107), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n428), .B1(new_n429), .B2(new_n268), .C1(new_n304), .C2(new_n306), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n275), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n426), .B1(new_n340), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n432), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n277), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n432), .A2(new_n411), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n426), .B1(new_n434), .B2(new_n298), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR4_X1   g0239(.A1(new_n302), .A2(new_n347), .A3(new_n417), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n225), .A2(G33), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n290), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT79), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(new_n291), .A4(G116), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n290), .A2(new_n441), .A3(new_n212), .A4(new_n279), .ZN(new_n445));
  INV_X1    g0245(.A(G116), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT79), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n444), .A2(new_n447), .B1(new_n446), .B2(new_n318), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G283), .ZN(new_n449));
  INV_X1    g0249(.A(G97), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n449), .B(new_n213), .C1(G33), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n446), .A2(G20), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n280), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT80), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT20), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n455), .B2(new_n453), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n453), .B2(new_n455), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n448), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT5), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n225), .B(G45), .C1(new_n460), .C2(G41), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT67), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n263), .ZN(new_n464));
  NAND2_X1  g0264(.A1(KEYINPUT67), .A2(G41), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n460), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n275), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n257), .A2(new_n256), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n461), .B1(new_n468), .B2(new_n460), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n467), .A2(G270), .B1(new_n469), .B2(G274), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n352), .A2(new_n354), .A3(G264), .A4(G1698), .ZN(new_n471));
  INV_X1    g0271(.A(G303), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(new_n268), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n268), .A2(G257), .A3(new_n269), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n275), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n340), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n459), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT21), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n470), .A2(new_n475), .A3(G179), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n477), .A2(new_n478), .B1(new_n459), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT81), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n477), .B2(new_n478), .ZN(new_n483));
  INV_X1    g0283(.A(new_n459), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n470), .A2(new_n475), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G200), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n484), .B(new_n486), .C1(new_n411), .C2(new_n485), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n459), .A2(new_n476), .A3(KEYINPUT81), .A4(KEYINPUT21), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n481), .A2(new_n483), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT19), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n213), .B1(new_n303), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G87), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n450), .A3(new_n429), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n352), .A2(new_n354), .A3(new_n213), .A4(G68), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n490), .B1(new_n284), .B2(new_n450), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n280), .ZN(new_n498));
  INV_X1    g0298(.A(new_n421), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n318), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT78), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT78), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n498), .A2(new_n503), .A3(new_n500), .ZN(new_n504));
  INV_X1    g0304(.A(new_n445), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n502), .A2(new_n504), .B1(G87), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n225), .A2(G45), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n259), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n507), .B(KEYINPUT77), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n264), .A2(G250), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n352), .A2(new_n354), .A3(G244), .A4(G1698), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n352), .A2(new_n354), .A3(G238), .A4(new_n269), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n275), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n298), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n511), .A2(new_n516), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(G190), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n506), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n352), .A2(new_n354), .A3(G244), .A4(new_n269), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n269), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n449), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n275), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n467), .A2(G257), .B1(new_n469), .B2(G274), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G200), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n531), .A2(new_n450), .A3(G107), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n531), .B2(new_n246), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n533), .A2(new_n213), .B1(new_n271), .B2(new_n287), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n429), .B1(new_n368), .B2(new_n369), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n280), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n505), .A2(G97), .ZN(new_n537));
  OR3_X1    g0337(.A1(new_n290), .A2(KEYINPUT76), .A3(G97), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT76), .B1(new_n290), .B2(G97), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n527), .A2(G190), .A3(new_n528), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n530), .A2(new_n536), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(G169), .B1(new_n511), .B2(new_n516), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n277), .B2(new_n518), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n505), .A2(new_n421), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n498), .A2(new_n503), .A3(new_n500), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n503), .B1(new_n498), .B2(new_n500), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n529), .A2(new_n340), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n536), .A2(new_n541), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n527), .A2(new_n277), .A3(new_n528), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n520), .A2(new_n543), .A3(new_n550), .A4(new_n554), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n489), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n352), .A2(new_n354), .A3(G250), .A4(new_n269), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n352), .A2(new_n354), .A3(G257), .A4(G1698), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G294), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n275), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n469), .A2(G274), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n462), .A2(new_n466), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(G264), .A3(new_n264), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n277), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n275), .A2(new_n560), .B1(new_n467), .B2(G264), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT84), .B1(new_n567), .B2(new_n562), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n561), .A2(KEYINPUT84), .A3(new_n564), .A4(new_n562), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(G169), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n566), .B1(new_n571), .B2(KEYINPUT85), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT84), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n565), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n340), .B1(new_n574), .B2(new_n569), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT85), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n352), .A2(new_n354), .A3(new_n213), .A4(G87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT22), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT22), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n268), .A2(new_n580), .A3(new_n213), .A4(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n514), .A2(G20), .ZN(new_n583));
  OR2_X1    g0383(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n584));
  NAND2_X1  g0384(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(new_n585), .C1(new_n213), .C2(G107), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n429), .A2(KEYINPUT82), .A3(KEYINPUT23), .A4(G20), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT24), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n582), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n582), .B2(new_n588), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n280), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT83), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT83), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n594), .B(new_n280), .C1(new_n590), .C2(new_n591), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n318), .A2(KEYINPUT25), .A3(new_n429), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT25), .B1(new_n318), .B2(new_n429), .ZN(new_n599));
  OAI22_X1  g0399(.A1(new_n598), .A2(new_n599), .B1(new_n429), .B2(new_n445), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n572), .A2(new_n577), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n574), .A2(new_n411), .A3(new_n569), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n565), .A2(new_n298), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n596), .A2(new_n605), .A3(new_n601), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT86), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n582), .A2(new_n588), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT24), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n582), .A2(new_n588), .A3(new_n589), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n594), .B1(new_n611), .B2(new_n280), .ZN(new_n612));
  INV_X1    g0412(.A(new_n595), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n601), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n577), .ZN(new_n615));
  INV_X1    g0415(.A(new_n566), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n575), .B2(new_n576), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n614), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT86), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n596), .A2(new_n605), .A3(new_n601), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n556), .B1(new_n607), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n440), .A2(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n555), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n481), .A2(new_n483), .A3(new_n488), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n620), .B(new_n624), .C1(new_n602), .C2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n550), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n520), .A2(new_n550), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(new_n554), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n506), .A2(new_n519), .B1(new_n545), .B2(new_n549), .ZN(new_n631));
  INV_X1    g0431(.A(new_n554), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(KEYINPUT26), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n627), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n440), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n295), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n351), .B(new_n414), .C1(new_n367), .C2(new_n376), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT17), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n405), .A2(new_n409), .A3(new_n414), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n436), .B1(new_n335), .B2(new_n336), .ZN(new_n642));
  INV_X1    g0442(.A(new_n346), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n377), .A2(new_n400), .A3(KEYINPUT18), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n407), .B1(new_n405), .B2(new_n406), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n300), .A2(new_n301), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n637), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n636), .A2(new_n650), .ZN(G369));
  AND2_X1   g0451(.A1(new_n213), .A2(G13), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n225), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n484), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n625), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT87), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n660), .B1(new_n489), .B2(KEYINPUT88), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(KEYINPUT88), .B2(new_n489), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g0465(.A(new_n665), .B(KEYINPUT89), .Z(new_n666));
  NAND2_X1  g0466(.A1(new_n614), .A2(new_n658), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n602), .A2(new_n606), .A3(KEYINPUT86), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n619), .B1(new_n618), .B2(new_n620), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n602), .A2(new_n658), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n666), .A2(G330), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n625), .A2(new_n659), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n607), .B2(new_n621), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n618), .A2(new_n658), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n677), .ZN(G399));
  NOR2_X1   g0478(.A1(new_n229), .A2(new_n468), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n493), .A2(G116), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n210), .B2(new_n680), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n635), .A2(KEYINPUT92), .A3(new_n659), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n658), .B1(new_n626), .B2(new_n634), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(KEYINPUT92), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n685), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT93), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g0491(.A(KEYINPUT93), .B(new_n685), .C1(new_n686), .C2(new_n688), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n550), .B(KEYINPUT94), .Z(new_n693));
  AND2_X1   g0493(.A1(new_n481), .A2(new_n483), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n618), .A2(new_n488), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n606), .A2(new_n555), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT26), .B1(new_n631), .B2(new_n632), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n633), .B1(new_n698), .B2(KEYINPUT95), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT95), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n631), .A2(new_n700), .A3(KEYINPUT26), .A4(new_n632), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n658), .B1(new_n697), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n691), .A2(new_n692), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n518), .A2(new_n567), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n706), .A2(new_n529), .A3(new_n479), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(KEYINPUT30), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT91), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n518), .A2(G179), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n565), .A3(new_n529), .A4(new_n485), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n707), .A2(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n709), .ZN(new_n715));
  INV_X1    g0515(.A(new_n708), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n659), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n489), .A2(new_n555), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n719), .B(new_n659), .C1(new_n668), .C2(new_n669), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n718), .B1(new_n720), .B2(KEYINPUT31), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n716), .A2(new_n714), .A3(new_n712), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT90), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(G330), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n705), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n684), .B1(new_n728), .B2(G1), .ZN(G364));
  AOI21_X1  g0529(.A(new_n225), .B1(new_n652), .B2(G45), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n680), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n662), .A2(new_n664), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n212), .B1(G20), .B2(new_n340), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G179), .A2(G200), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n213), .B1(new_n738), .B2(G190), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n450), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n738), .A2(G20), .A3(new_n411), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G159), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT32), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n213), .A2(new_n277), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G190), .ZN(new_n747));
  AOI211_X1 g0547(.A(new_n740), .B(new_n744), .C1(G68), .C2(new_n747), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n745), .A2(KEYINPUT98), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n745), .A2(KEYINPUT98), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G190), .A2(G200), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G77), .ZN(new_n754));
  NOR4_X1   g0554(.A1(new_n213), .A2(new_n411), .A3(new_n298), .A4(G179), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n492), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n746), .A2(new_n411), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n355), .B(new_n757), .C1(G50), .C2(new_n758), .ZN(new_n759));
  NOR4_X1   g0559(.A1(new_n213), .A2(new_n298), .A3(G179), .A4(G190), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT99), .Z(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n411), .A2(G200), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n749), .A2(new_n750), .A3(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n762), .A2(G107), .B1(G58), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n748), .A2(new_n754), .A3(new_n759), .A4(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n762), .A2(G283), .B1(G322), .B2(new_n765), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n747), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n739), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n758), .A2(G326), .B1(G294), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n742), .A2(G329), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n355), .B(new_n773), .C1(new_n756), .C2(new_n472), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(G311), .B2(new_n753), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n768), .A2(new_n770), .A3(new_n772), .A4(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n737), .B1(new_n767), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n734), .A2(new_n736), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT97), .Z(new_n779));
  NOR2_X1   g0579(.A1(new_n229), .A2(new_n355), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G355), .A2(new_n780), .B1(new_n446), .B2(new_n229), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n355), .A2(new_n228), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT96), .Z(new_n783));
  INV_X1    g0583(.A(new_n255), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n210), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G45), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n253), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n781), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n777), .B1(new_n779), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n731), .B1(new_n735), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n666), .B(G330), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(new_n791), .B2(new_n731), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT100), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G396));
  INV_X1    g0594(.A(new_n731), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n433), .A2(new_n435), .A3(new_n658), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(KEYINPUT104), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n796), .A2(KEYINPUT104), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n426), .A2(new_n659), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n798), .A2(new_n799), .B1(new_n439), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n686), .B2(new_n688), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n687), .A2(new_n801), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n795), .B1(new_n805), .B2(new_n726), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n726), .B2(new_n805), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n736), .A2(new_n732), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n795), .B1(G77), .B2(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n762), .A2(G87), .B1(G116), .B2(new_n753), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT101), .B(G283), .Z(new_n812));
  NAND2_X1  g0612(.A1(new_n747), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n740), .B1(new_n758), .B2(G303), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n355), .B1(new_n741), .B2(new_n815), .C1(new_n756), .C2(new_n429), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G294), .B2(new_n765), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n811), .A2(new_n813), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G132), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n268), .B1(new_n741), .B2(new_n819), .C1(new_n756), .C2(new_n248), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n761), .A2(new_n203), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(G58), .C2(new_n771), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT103), .Z(new_n823));
  AOI22_X1  g0623(.A1(new_n747), .A2(G150), .B1(new_n758), .B2(G137), .ZN(new_n824));
  INV_X1    g0624(.A(G143), .ZN(new_n825));
  INV_X1    g0625(.A(G159), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n824), .B1(new_n825), .B2(new_n764), .C1(new_n826), .C2(new_n752), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT102), .B(KEYINPUT34), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n818), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n810), .B1(new_n830), .B2(new_n736), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n801), .B2(new_n733), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n807), .A2(new_n832), .ZN(G384));
  INV_X1    g0633(.A(new_n533), .ZN(new_n834));
  OAI211_X1 g0634(.A(G116), .B(new_n214), .C1(new_n834), .C2(KEYINPUT35), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(KEYINPUT35), .B2(new_n834), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT36), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n211), .A2(G77), .A3(new_n360), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n225), .B(G13), .C1(new_n838), .C2(new_n249), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n718), .A2(KEYINPUT31), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT31), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n622), .B2(new_n659), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n841), .B1(new_n843), .B2(new_n718), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n440), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT108), .Z(new_n846));
  NAND2_X1  g0646(.A1(new_n338), .A2(new_n658), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n337), .B2(new_n346), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n337), .A2(new_n346), .A3(new_n847), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n802), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n718), .A2(KEYINPUT31), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n721), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n405), .A2(new_n406), .ZN(new_n855));
  AOI221_X4 g0655(.A(new_n350), .B1(new_n413), .B2(new_n412), .C1(new_n404), .C2(new_n375), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n858));
  INV_X1    g0658(.A(new_n656), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n377), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n857), .A2(KEYINPUT107), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n377), .A2(new_n400), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(new_n860), .A3(new_n638), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n405), .A2(new_n656), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n858), .B1(new_n864), .B2(KEYINPUT107), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n860), .B1(new_n647), .B2(new_n641), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n854), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n374), .A2(new_n280), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT105), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT105), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n374), .A2(new_n872), .A3(new_n280), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n366), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n656), .B1(new_n874), .B2(new_n351), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n417), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n858), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n862), .A2(new_n860), .A3(new_n638), .A4(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n406), .A2(new_n656), .B1(new_n874), .B2(new_n351), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n879), .B2(new_n856), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n869), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT40), .B1(new_n853), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n878), .A2(new_n880), .ZN(new_n885));
  INV_X1    g0685(.A(new_n875), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n647), .B2(new_n641), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n854), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT40), .B1(new_n888), .B2(new_n882), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n844), .A2(new_n889), .A3(new_n851), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(G330), .B1(new_n846), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n891), .B2(new_n846), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n691), .A2(new_n440), .A3(new_n692), .A4(new_n704), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n650), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n893), .B(new_n895), .Z(new_n896));
  NOR3_X1   g0696(.A1(new_n885), .A2(new_n887), .A3(new_n854), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n876), .B2(new_n881), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT39), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n869), .A2(new_n900), .A3(new_n882), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n643), .A2(new_n659), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n436), .A2(new_n658), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n687), .B2(new_n801), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n849), .A2(new_n850), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n907), .B(new_n908), .C1(new_n897), .C2(new_n898), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n647), .B2(new_n859), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n896), .A2(new_n911), .B1(new_n225), .B2(new_n652), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n896), .A2(new_n911), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n840), .B1(new_n912), .B2(new_n913), .ZN(G367));
  XNOR2_X1  g0714(.A(new_n730), .B(KEYINPUT112), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n632), .A2(new_n658), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n552), .A2(new_n658), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n543), .A2(new_n554), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n677), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT44), .ZN(new_n921));
  INV_X1    g0721(.A(new_n919), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n675), .A2(new_n676), .A3(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT45), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n673), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n673), .A2(new_n921), .A3(new_n924), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n666), .A2(G330), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n675), .A2(KEYINPUT110), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n672), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n675), .B1(new_n934), .B2(new_n674), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT110), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n931), .B(new_n933), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(G330), .A3(new_n666), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n930), .A2(KEYINPUT111), .A3(new_n728), .A4(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT111), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n728), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n942), .B1(new_n943), .B2(new_n929), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n727), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n679), .B(KEYINPUT41), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n915), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n506), .A2(new_n659), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT109), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n629), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n627), .B2(new_n950), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT43), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n675), .A2(new_n919), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n554), .B1(new_n618), .B2(new_n918), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n955), .A2(KEYINPUT42), .B1(new_n659), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n954), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n952), .A2(new_n953), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n673), .A2(new_n922), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n948), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n952), .A2(new_n734), .ZN(new_n965));
  INV_X1    g0765(.A(new_n760), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n355), .B1(new_n966), .B2(new_n450), .ZN(new_n967));
  INV_X1    g0767(.A(new_n758), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n968), .A2(new_n815), .B1(new_n739), .B2(new_n429), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n967), .B(new_n969), .C1(G317), .C2(new_n742), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT46), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n756), .B2(new_n446), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n755), .A2(KEYINPUT46), .A3(G116), .ZN(new_n973));
  INV_X1    g0773(.A(G294), .ZN(new_n974));
  INV_X1    g0774(.A(new_n747), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n972), .B(new_n973), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT113), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  INV_X1    g0779(.A(new_n812), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n472), .A2(new_n764), .B1(new_n752), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n970), .A2(new_n978), .A3(new_n979), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n771), .A2(G68), .ZN(new_n984));
  INV_X1    g0784(.A(G137), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n984), .B1(new_n985), .B2(new_n741), .C1(new_n756), .C2(new_n202), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n355), .B1(new_n760), .B2(G77), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT114), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n248), .A2(new_n752), .B1(new_n764), .B2(new_n285), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n975), .A2(new_n826), .B1(new_n968), .B2(new_n825), .ZN(new_n990));
  OR4_X1    g0790(.A1(new_n986), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n983), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT47), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(KEYINPUT47), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(new_n736), .A3(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n783), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n778), .B1(new_n228), .B2(new_n499), .C1(new_n996), .C2(new_n243), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n995), .A2(new_n795), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n965), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n964), .A2(new_n1000), .ZN(G387));
  NOR2_X1   g0801(.A1(new_n283), .A2(G50), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(KEYINPUT115), .B2(new_n681), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n786), .B1(new_n203), .B2(new_n271), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1005), .B(new_n1007), .C1(KEYINPUT115), .C2(new_n681), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1008), .B(new_n783), .C1(new_n240), .C2(new_n255), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n780), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1009), .B1(G107), .B2(new_n228), .C1(new_n681), .C2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n731), .B1(new_n1011), .B2(new_n779), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n771), .A2(new_n421), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n975), .B2(new_n283), .C1(new_n826), .C2(new_n968), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n761), .A2(new_n450), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n755), .A2(G77), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1016), .B(new_n268), .C1(new_n285), .C2(new_n741), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n248), .A2(new_n764), .B1(new_n752), .B2(new_n203), .ZN(new_n1018));
  NOR4_X1   g0818(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n747), .A2(G311), .B1(new_n758), .B2(G322), .ZN(new_n1020));
  INV_X1    g0820(.A(G317), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n472), .B2(new_n752), .C1(new_n1021), .C2(new_n764), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n974), .B2(new_n756), .C1(new_n739), .C2(new_n980), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT49), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n966), .A2(new_n446), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n268), .B(new_n1026), .C1(G326), .C2(new_n742), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1019), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1012), .B1(new_n1028), .B2(new_n737), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT117), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n934), .B2(new_n734), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n915), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1031), .B1(new_n940), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n943), .A2(new_n679), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n940), .A2(new_n728), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(G393));
  NAND2_X1  g0836(.A1(new_n930), .A2(new_n1032), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n922), .A2(new_n734), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n765), .A2(G311), .B1(G317), .B2(new_n758), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT52), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n268), .B1(new_n742), .B2(G322), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n756), .B2(new_n980), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n975), .A2(new_n472), .B1(new_n739), .B2(new_n446), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n761), .A2(new_n429), .B1(new_n974), .B2(new_n752), .ZN(new_n1044));
  NOR4_X1   g0844(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n739), .A2(new_n271), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n268), .B1(new_n741), .B2(new_n825), .C1(new_n756), .C2(new_n203), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(G50), .C2(new_n747), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n826), .A2(new_n764), .B1(new_n968), .B2(new_n285), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT51), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n762), .A2(G87), .B1(new_n348), .B2(new_n753), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1048), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n736), .B1(new_n1045), .B2(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n778), .B1(new_n450), .B2(new_n228), .C1(new_n996), .C2(new_n247), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1038), .A2(new_n795), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1037), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n941), .A2(new_n944), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n680), .B1(new_n943), .B2(new_n929), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(G390));
  INV_X1    g0863(.A(KEYINPUT118), .ZN(new_n1064));
  INV_X1    g0864(.A(G330), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n802), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n908), .B(new_n1066), .C1(new_n721), .C2(new_n725), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n905), .B1(new_n703), .B2(new_n801), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n908), .B1(new_n844), .B2(new_n1066), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1064), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n337), .A2(new_n346), .A3(new_n847), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1072), .A2(new_n848), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n720), .A2(KEYINPUT31), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n718), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n852), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1066), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1078), .A2(KEYINPUT118), .A3(new_n1068), .A4(new_n1067), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1071), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1066), .B1(new_n721), .B2(new_n725), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n1073), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n844), .A2(G330), .A3(new_n851), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n906), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n903), .B1(new_n906), .B2(new_n1073), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(new_n899), .A3(new_n901), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n869), .A2(new_n882), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1089), .B(new_n903), .C1(new_n1068), .C2(new_n1073), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1083), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1088), .A2(new_n1090), .A3(new_n1067), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n844), .A2(G330), .A3(new_n440), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n894), .A2(new_n650), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1086), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1084), .B1(new_n1071), .B2(new_n1079), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n1097), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1099), .A2(new_n679), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n902), .A2(new_n732), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n795), .B1(new_n348), .B2(new_n809), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n975), .A2(new_n429), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1046), .B(new_n1106), .C1(G283), .C2(new_n758), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n268), .B(new_n757), .C1(G294), .C2(new_n742), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n821), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G97), .A2(new_n753), .B1(new_n765), .B2(G116), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n739), .A2(new_n826), .ZN(new_n1112));
  INV_X1    g0912(.A(G125), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n268), .B1(new_n1113), .B2(new_n741), .C1(new_n966), .C2(new_n248), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1112), .B(new_n1114), .C1(G128), .C2(new_n758), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT54), .B(G143), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT119), .Z(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1115), .B1(new_n819), .B2(new_n764), .C1(new_n752), .C2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1120));
  OR3_X1    g0920(.A1(new_n756), .A2(new_n285), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n756), .B2(new_n285), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(new_n985), .C2(new_n975), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1111), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1105), .B1(new_n1124), .B2(new_n736), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1095), .A2(new_n1032), .B1(new_n1104), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1103), .A2(new_n1126), .ZN(G378));
  OAI21_X1  g0927(.A(new_n1098), .B1(new_n1101), .B2(new_n1100), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n296), .A2(new_n656), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT124), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n302), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n302), .A2(new_n1132), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1131), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n302), .A2(new_n1132), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n1133), .A3(new_n1130), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n844), .A2(new_n1089), .A3(new_n851), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n801), .B1(new_n1072), .B2(new_n848), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n841), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1140), .A2(KEYINPUT40), .B1(new_n1143), .B2(new_n889), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1139), .B1(new_n1144), .B2(new_n1065), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1139), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n891), .A2(G330), .A3(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n904), .A2(new_n910), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1128), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n680), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1128), .A2(KEYINPUT57), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1146), .B1(new_n891), .B2(G330), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1065), .B(new_n1139), .C1(new_n884), .C2(new_n890), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n911), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT125), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1158), .A2(KEYINPUT125), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1154), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1153), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1032), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n731), .B1(new_n248), .B2(new_n808), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n984), .B1(new_n975), .B2(new_n450), .C1(new_n446), .C2(new_n968), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n966), .A2(new_n202), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n468), .A2(new_n268), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1016), .A2(new_n1167), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(G283), .C2(new_n742), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n429), .B2(new_n764), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1165), .B(new_n1170), .C1(new_n421), .C2(new_n753), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT122), .Z(new_n1172));
  OR2_X1    g0972(.A1(new_n1172), .A2(KEYINPUT58), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(KEYINPUT58), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G50), .B(new_n1167), .C1(new_n262), .C2(new_n263), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT121), .Z(new_n1176));
  AOI22_X1  g0976(.A1(new_n753), .A2(G137), .B1(G132), .B2(new_n747), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n765), .A2(G128), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n756), .C2(new_n1118), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n758), .A2(G125), .B1(G150), .B2(new_n771), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT123), .Z(new_n1181));
  NOR2_X1   g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n262), .B(new_n263), .C1(new_n966), .C2(new_n826), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G124), .B2(new_n742), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  AND4_X1   g0988(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .A4(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1164), .B1(new_n1146), .B2(new_n733), .C1(new_n1189), .C2(new_n737), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1163), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1162), .A2(new_n1192), .ZN(G375));
  NAND2_X1  g0993(.A1(new_n1086), .A2(new_n1032), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n731), .B1(new_n203), .B2(new_n808), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n355), .B1(new_n741), .B2(new_n472), .C1(new_n756), .C2(new_n450), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n761), .A2(new_n271), .B1(new_n429), .B2(new_n752), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(G283), .C2(new_n765), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1013), .B1(new_n975), .B2(new_n446), .C1(new_n974), .C2(new_n968), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n968), .A2(new_n819), .B1(new_n739), .B2(new_n248), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n742), .A2(G128), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n756), .B2(new_n826), .ZN(new_n1203));
  NOR4_X1   g1003(.A1(new_n1201), .A2(new_n1203), .A3(new_n355), .A4(new_n1166), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1118), .A2(new_n975), .B1(new_n985), .B2(new_n764), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G150), .B2(new_n753), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1198), .A2(new_n1200), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1195), .B1(new_n737), .B2(new_n1207), .C1(new_n908), .C2(new_n733), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1194), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1086), .A2(new_n1098), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1080), .A2(new_n1097), .A3(new_n1085), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n946), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1209), .A2(new_n1212), .ZN(G381));
  AOI21_X1  g1013(.A(new_n1191), .B1(new_n1153), .B2(new_n1161), .ZN(new_n1214));
  INV_X1    g1014(.A(G378), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(G384), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G396), .A2(G393), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1062), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  OR4_X1    g1019(.A1(G387), .A2(new_n1216), .A3(G381), .A4(new_n1219), .ZN(G407));
  OAI211_X1 g1020(.A(G407), .B(G213), .C1(G343), .C2(new_n1216), .ZN(G409));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n657), .A2(G213), .A3(G2897), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT60), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1211), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1101), .A2(KEYINPUT60), .A3(new_n1097), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n1210), .A3(new_n679), .A4(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1228), .A2(G384), .A3(new_n1209), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G384), .B1(new_n1228), .B2(new_n1209), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1224), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1211), .A2(new_n1225), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n679), .B1(new_n1101), .B2(new_n1097), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT60), .B1(new_n1101), .B2(new_n1097), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1194), .A2(new_n1208), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1217), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1228), .A2(new_n1209), .A3(G384), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1223), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1231), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G375), .A2(G378), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT125), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1158), .A2(KEYINPUT125), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n915), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n946), .B(new_n1128), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1103), .A2(new_n1126), .A3(new_n1190), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1248), .A2(new_n1249), .B1(G213), .B2(new_n657), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1240), .B1(new_n1241), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1222), .B1(new_n1251), .B2(KEYINPUT61), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n657), .A2(G213), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1032), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1249), .A2(new_n1255), .A3(new_n1246), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1253), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1253), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1241), .A2(new_n1250), .A3(new_n1258), .A4(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(new_n1261), .A3(new_n1263), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1229), .A2(new_n1230), .A3(new_n1224), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1223), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT61), .B1(new_n1267), .B2(new_n1257), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT126), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1252), .A2(new_n1264), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G387), .A2(new_n1062), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G393), .B(new_n793), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n964), .A2(G390), .A3(new_n1000), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1272), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G390), .B1(new_n964), .B2(new_n1000), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n999), .B(new_n1062), .C1(new_n948), .C2(new_n963), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1275), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1274), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1270), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1241), .A2(new_n1250), .A3(KEYINPUT63), .A4(new_n1258), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1284), .A2(new_n1274), .A3(new_n1278), .A4(new_n1268), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1280), .A2(new_n1285), .ZN(G405));
  NAND2_X1  g1086(.A1(new_n1241), .A2(new_n1216), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1287), .B(new_n1259), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(new_n1279), .ZN(G402));
endmodule


