//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  AND2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G155gat), .B(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT2), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n206), .B1(new_n205), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT29), .ZN(new_n214));
  NOR2_X1   g013(.A1(G197gat), .A2(G204gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(G197gat), .A2(G204gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G211gat), .A2(G218gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  OAI22_X1  g018(.A1(new_n215), .A2(new_n217), .B1(new_n219), .B2(KEYINPUT22), .ZN(new_n220));
  NOR2_X1   g019(.A1(G211gat), .A2(G218gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT72), .ZN(new_n222));
  NOR3_X1   g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G197gat), .ZN(new_n225));
  INV_X1    g024(.A(G204gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n227), .A2(new_n216), .B1(new_n228), .B2(new_n218), .ZN(new_n229));
  INV_X1    g028(.A(G211gat), .ZN(new_n230));
  INV_X1    g029(.A(G218gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(KEYINPUT72), .A3(new_n218), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n214), .B1(new_n224), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT83), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT3), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n223), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n229), .A2(new_n233), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT29), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT83), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n213), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n204), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT2), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT76), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT76), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT2), .ZN(new_n247));
  NAND2_X1  g046(.A1(G141gat), .A2(G148gat), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n243), .A2(new_n245), .A3(new_n247), .A4(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n206), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n214), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT73), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT73), .B1(new_n238), .B2(new_n239), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G228gat), .ZN(new_n260));
  INV_X1    g059(.A(G233gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n202), .B1(new_n242), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n213), .ZN(new_n265));
  INV_X1    g064(.A(new_n241), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n252), .B1(new_n240), .B2(KEYINPUT83), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n262), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(new_n224), .B2(new_n234), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n256), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n269), .B1(new_n272), .B2(new_n255), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(KEYINPUT84), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n259), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n220), .B1(new_n219), .B2(new_n221), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n229), .A2(new_n218), .A3(new_n232), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n214), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n213), .B1(new_n278), .B2(new_n252), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n269), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G22gat), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n264), .A2(new_n274), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT85), .ZN(new_n283));
  XOR2_X1   g082(.A(G78gat), .B(G106gat), .Z(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT31), .B(G50gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n264), .A2(new_n274), .A3(new_n280), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G22gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n282), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n287), .B(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G1gat), .B(G29gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT0), .ZN(new_n293));
  XNOR2_X1  g092(.A(G57gat), .B(G85gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  OAI21_X1  g094(.A(KEYINPUT3), .B1(new_n210), .B2(new_n212), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n254), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298));
  INV_X1    g097(.A(G134gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(G127gat), .ZN(new_n300));
  INV_X1    g099(.A(G127gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G134gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n306));
  OAI21_X1  g105(.A(G120gat), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n308));
  INV_X1    g107(.A(G120gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(new_n304), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n303), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G113gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(new_n309), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n298), .B1(G113gat), .B2(G120gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n299), .ZN(new_n317));
  NAND2_X1  g116(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(G127gat), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n299), .A2(G127gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(new_n322), .B2(KEYINPUT70), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n311), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT77), .B1(new_n297), .B2(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n328), .A2(new_n329), .A3(new_n301), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT70), .B1(new_n330), .B2(new_n320), .ZN(new_n331));
  INV_X1    g130(.A(new_n315), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n325), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n311), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n254), .A4(new_n296), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT5), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n333), .A2(new_n334), .A3(new_n213), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(KEYINPUT80), .A3(KEYINPUT4), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n344));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n213), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT80), .B1(new_n342), .B2(KEYINPUT4), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n338), .B(new_n341), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT81), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n342), .A2(KEYINPUT4), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(new_n343), .A3(new_n345), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n338), .A4(new_n341), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n335), .A2(new_n265), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n339), .B1(new_n357), .B2(new_n342), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n359));
  OR3_X1    g158(.A1(new_n358), .A2(KEYINPUT79), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n342), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n340), .B1(new_n361), .B2(KEYINPUT4), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n344), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n338), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT79), .B1(new_n358), .B2(new_n359), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n295), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT23), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT25), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(G169gat), .B2(G176gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n370), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G190gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT66), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT66), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G190gat), .ZN(new_n380));
  INV_X1    g179(.A(G183gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT65), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT65), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G183gat), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n378), .A2(new_n380), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT24), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n381), .A2(new_n377), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(new_n391), .A3(new_n389), .ZN(new_n392));
  NAND2_X1  g191(.A1(G169gat), .A2(G176gat), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n392), .A2(new_n372), .A3(new_n369), .A4(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT25), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n376), .A2(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT28), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n378), .A2(new_n380), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT27), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n399), .B1(new_n382), .B2(new_n384), .ZN(new_n400));
  NOR2_X1   g199(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n386), .ZN(new_n403));
  AND2_X1   g202(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n378), .B(new_n380), .C1(new_n404), .C2(new_n401), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n405), .B2(KEYINPUT28), .ZN(new_n406));
  INV_X1    g205(.A(G169gat), .ZN(new_n407));
  INV_X1    g206(.A(G176gat), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT26), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n407), .B(new_n408), .C1(new_n409), .C2(KEYINPUT67), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(KEYINPUT67), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n368), .A2(KEYINPUT67), .A3(new_n409), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n393), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n402), .A2(new_n406), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT68), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT68), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n402), .A2(new_n406), .A3(new_n417), .A4(new_n414), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n396), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G226gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(new_n261), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(KEYINPUT29), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n376), .A2(new_n390), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n394), .A2(new_n395), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n427), .A2(new_n415), .A3(new_n421), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n272), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n416), .A2(new_n418), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n427), .A3(new_n421), .ZN(new_n431));
  INV_X1    g230(.A(new_n272), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n415), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n422), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G8gat), .B(G36gat), .Z(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT74), .ZN(new_n437));
  XNOR2_X1  g236(.A(G64gat), .B(G92gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n429), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n430), .A2(new_n427), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n428), .B1(new_n442), .B2(new_n422), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n435), .B1(new_n443), .B2(new_n432), .ZN(new_n444));
  INV_X1    g243(.A(new_n439), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT75), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n441), .B1(new_n447), .B2(KEYINPUT30), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(KEYINPUT75), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n367), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n338), .B1(new_n346), .B2(new_n347), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n340), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT39), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n357), .A2(new_n342), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(new_n339), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n454), .A3(new_n340), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n295), .A3(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT40), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n291), .B1(new_n451), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT37), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n445), .B1(new_n444), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT38), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n443), .A2(new_n432), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n431), .A2(new_n434), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n465), .B(KEYINPUT37), .C1(new_n432), .C2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n429), .A2(KEYINPUT37), .A3(new_n435), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n464), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n439), .B1(new_n429), .B2(new_n435), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n356), .A2(new_n295), .A3(new_n366), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT82), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n356), .A2(new_n366), .ZN(new_n476));
  INV_X1    g275(.A(new_n295), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT6), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n356), .A2(KEYINPUT82), .A3(new_n366), .A4(new_n295), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n367), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n472), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n461), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n480), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n478), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT75), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT30), .B1(new_n471), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n450), .A2(new_n488), .A3(new_n440), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n367), .B1(new_n474), .B2(new_n473), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n486), .B(new_n489), .C1(new_n490), .C2(KEYINPUT6), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n291), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n493));
  AOI211_X1 g292(.A(new_n396), .B(new_n326), .C1(new_n416), .C2(new_n418), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n335), .B1(new_n430), .B2(new_n427), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G227gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(new_n261), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT34), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT34), .ZN(new_n500));
  INV_X1    g299(.A(new_n498), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n500), .B(new_n501), .C1(new_n494), .C2(new_n495), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT33), .B1(new_n496), .B2(new_n498), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G43gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(G71gat), .B(G99gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n499), .B(new_n502), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n442), .A2(new_n326), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n419), .A2(new_n335), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(new_n498), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT33), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n506), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n508), .A2(new_n509), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n500), .B1(new_n513), .B2(new_n501), .ZN(new_n514));
  INV_X1    g313(.A(new_n502), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(KEYINPUT32), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n507), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n507), .B2(new_n516), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n493), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n507), .A2(new_n516), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n517), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n516), .A3(new_n518), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(KEYINPUT36), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n484), .A2(new_n492), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT35), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT85), .ZN(new_n529));
  AND4_X1   g328(.A1(new_n529), .A2(new_n289), .A3(new_n282), .A4(new_n286), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n283), .A2(new_n286), .B1(new_n289), .B2(new_n282), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(new_n523), .A3(new_n489), .A4(new_n524), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n533), .A2(KEYINPUT86), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n479), .A2(new_n482), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n528), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n519), .A2(new_n520), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n537), .A2(new_n538), .A3(new_n532), .A4(new_n489), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n486), .B1(new_n490), .B2(KEYINPUT6), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n539), .A2(KEYINPUT35), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n527), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT87), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT35), .B1(new_n539), .B2(new_n540), .ZN(new_n545));
  AND4_X1   g344(.A1(new_n532), .A2(new_n523), .A3(new_n489), .A4(new_n524), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n546), .A2(new_n535), .A3(new_n538), .A4(new_n528), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(KEYINPUT87), .A3(new_n527), .ZN(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G22gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT16), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(G1gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(G1gat), .B2(new_n550), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G8gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n556));
  NAND2_X1  g355(.A1(G29gat), .A2(G36gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT88), .ZN(new_n560));
  NOR2_X1   g359(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n561));
  INV_X1    g360(.A(G36gat), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(KEYINPUT88), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n558), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(G43gat), .A2(G50gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(G43gat), .A2(G50gat), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT15), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n556), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n559), .A2(new_n560), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n561), .A2(new_n562), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n571), .A3(new_n564), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n557), .ZN(new_n573));
  INV_X1    g372(.A(new_n568), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(KEYINPUT89), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT91), .B(G50gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(G43gat), .ZN(new_n578));
  OR2_X1    g377(.A1(KEYINPUT90), .A2(G43gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(KEYINPUT90), .A2(G43gat), .ZN(new_n580));
  AOI21_X1  g379(.A(G50gat), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n576), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n558), .B1(new_n571), .B2(new_n559), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n583), .A2(new_n568), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n569), .A2(new_n575), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n555), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT92), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n587), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n582), .A2(new_n584), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT89), .B1(new_n573), .B2(new_n574), .ZN(new_n591));
  AOI211_X1 g390(.A(new_n556), .B(new_n568), .C1(new_n572), .C2(new_n557), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(KEYINPUT92), .A3(KEYINPUT17), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n554), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n586), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n585), .A2(new_n588), .A3(new_n587), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT17), .B1(new_n593), .B2(KEYINPUT92), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n555), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT93), .ZN(new_n601));
  NAND2_X1  g400(.A1(G229gat), .A2(G233gat), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n597), .A2(new_n601), .A3(KEYINPUT18), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n593), .B(new_n554), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n602), .B(KEYINPUT13), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G113gat), .B(G141gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G197gat), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT11), .B(G169gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n603), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT18), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT94), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(KEYINPUT94), .A3(new_n614), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n612), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n615), .A2(new_n606), .A3(new_n603), .ZN(new_n620));
  INV_X1    g419(.A(new_n611), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT95), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n619), .A2(new_n622), .A3(KEYINPUT95), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT21), .ZN(new_n628));
  INV_X1    g427(.A(G64gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(G57gat), .ZN(new_n630));
  INV_X1    g429(.A(G57gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT97), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(G57gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n630), .B1(new_n635), .B2(new_n629), .ZN(new_n636));
  NAND2_X1  g435(.A1(G71gat), .A2(G78gat), .ZN(new_n637));
  OR2_X1    g436(.A1(G71gat), .A2(G78gat), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT9), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT96), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n631), .A2(G64gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n630), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT9), .ZN(new_n645));
  XOR2_X1   g444(.A(G71gat), .B(G78gat), .Z(new_n646));
  AOI21_X1  g445(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n639), .B1(new_n630), .B2(new_n643), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n638), .A2(new_n637), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT96), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n641), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n555), .B1(new_n628), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n628), .ZN(new_n656));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  XNOR2_X1  g457(.A(G127gat), .B(G155gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT98), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G183gat), .B(G211gat), .Z(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n655), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n661), .A2(new_n662), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n654), .A3(new_n663), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G190gat), .B(G218gat), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n671));
  INV_X1    g470(.A(G92gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT100), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(G92gat), .ZN(new_n675));
  INV_X1    g474(.A(G85gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(G85gat), .A2(G92gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT7), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT7), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(G85gat), .A3(G92gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(G99gat), .ZN(new_n683));
  INV_X1    g482(.A(G106gat), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT8), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n677), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(G99gat), .B(G106gat), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n677), .A2(new_n682), .A3(new_n687), .A4(new_n685), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n598), .B2(new_n599), .ZN(new_n692));
  INV_X1    g491(.A(new_n691), .ZN(new_n693));
  AND2_X1   g492(.A1(G232gat), .A2(G233gat), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n593), .A2(new_n693), .B1(KEYINPUT41), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n671), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n693), .B1(new_n589), .B2(new_n594), .ZN(new_n697));
  INV_X1    g496(.A(new_n695), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n697), .A2(KEYINPUT101), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n670), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT101), .B1(new_n697), .B2(new_n698), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n692), .A2(new_n671), .A3(new_n695), .ZN(new_n702));
  INV_X1    g501(.A(new_n670), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n700), .A2(KEYINPUT99), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n694), .A2(KEYINPUT41), .ZN(new_n706));
  XNOR2_X1  g505(.A(G134gat), .B(G162gat), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n706), .B(new_n707), .Z(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n700), .A2(KEYINPUT99), .A3(new_n704), .A4(new_n708), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n669), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(G230gat), .A2(G233gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(G57gat), .B(G64gat), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n646), .B(new_n642), .C1(new_n639), .C2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT96), .B1(new_n648), .B2(new_n649), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n719), .A2(new_n641), .A3(new_n690), .A4(new_n689), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT10), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n651), .A2(new_n691), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(KEYINPUT102), .A3(new_n720), .ZN(new_n724));
  OR3_X1    g523(.A1(new_n651), .A2(new_n691), .A3(KEYINPUT102), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n722), .B1(new_n726), .B2(new_n721), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n715), .B1(new_n727), .B2(KEYINPUT103), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT10), .B1(new_n724), .B2(new_n725), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n729), .A2(new_n730), .A3(new_n722), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n715), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n724), .A2(new_n725), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(G120gat), .B(G148gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(G176gat), .B(G204gat), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n735), .B(new_n736), .Z(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n734), .B1(new_n727), .B2(new_n733), .ZN(new_n741));
  INV_X1    g540(.A(new_n737), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n714), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n544), .A2(new_n549), .A3(new_n627), .A4(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n535), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(G1gat), .Z(G1324gat));
  AND3_X1   g547(.A1(new_n548), .A2(KEYINPUT87), .A3(new_n527), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT87), .B1(new_n548), .B2(new_n527), .ZN(new_n750));
  INV_X1    g549(.A(new_n627), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n489), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT16), .B(G8gat), .Z(new_n754));
  NAND4_X1  g553(.A1(new_n752), .A2(new_n753), .A3(new_n745), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G8gat), .B1(new_n746), .B2(new_n489), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT42), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n760), .B1(new_n755), .B2(new_n756), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n746), .A2(new_n489), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT42), .B1(new_n764), .B2(new_n754), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT104), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n762), .A2(new_n766), .ZN(G1325gat));
  OAI21_X1  g566(.A(G15gat), .B1(new_n746), .B2(new_n526), .ZN(new_n768));
  INV_X1    g567(.A(new_n537), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n769), .A2(G15gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n746), .B2(new_n770), .ZN(G1326gat));
  NOR2_X1   g570(.A1(new_n746), .A2(new_n532), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT43), .B(G22gat), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n772), .B(new_n773), .Z(G1327gat));
  NAND4_X1  g573(.A1(new_n544), .A2(KEYINPUT44), .A3(new_n549), .A4(new_n712), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n492), .A2(new_n776), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n461), .A2(new_n483), .B1(new_n525), .B2(new_n521), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n491), .A2(KEYINPUT106), .A3(new_n291), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n548), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n712), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n669), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n613), .A2(KEYINPUT94), .A3(new_n614), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT94), .B1(new_n613), .B2(new_n614), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n788), .A2(new_n612), .B1(new_n620), .B2(new_n621), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n785), .A2(new_n789), .A3(new_n744), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n775), .A2(new_n784), .A3(new_n540), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT107), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G29gat), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n791), .A2(KEYINPUT107), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n795));
  INV_X1    g594(.A(new_n744), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n669), .A2(new_n712), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT105), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n752), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n535), .A2(G29gat), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n795), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR4_X1   g601(.A1(new_n799), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n535), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n793), .A2(new_n794), .B1(new_n802), .B2(new_n803), .ZN(G1328gat));
  INV_X1    g603(.A(KEYINPUT46), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n489), .A2(G36gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n800), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT108), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n775), .A2(new_n784), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n753), .A3(new_n790), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G36gat), .ZN(new_n811));
  INV_X1    g610(.A(new_n806), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT46), .B1(new_n799), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT108), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n800), .A2(new_n814), .A3(new_n805), .A4(new_n806), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n808), .A2(new_n811), .A3(new_n813), .A4(new_n815), .ZN(G1329gat));
  OAI211_X1 g615(.A(new_n579), .B(new_n580), .C1(new_n799), .C2(new_n769), .ZN(new_n817));
  INV_X1    g616(.A(new_n526), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n579), .A2(new_n580), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n775), .A2(new_n784), .A3(new_n821), .A4(new_n790), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT47), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n817), .A2(new_n825), .A3(new_n822), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(G1330gat));
  OAI21_X1  g626(.A(new_n577), .B1(new_n799), .B2(new_n532), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n532), .A2(new_n577), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n775), .A2(new_n784), .A3(new_n790), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT48), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT48), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n833), .A3(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(G1331gat));
  NAND3_X1  g634(.A1(new_n713), .A2(new_n789), .A3(new_n744), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT109), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n837), .A2(KEYINPUT110), .A3(new_n781), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT110), .B1(new_n837), .B2(new_n781), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n540), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(new_n635), .ZN(G1332gat));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n489), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n837), .A2(new_n781), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n837), .A2(KEYINPUT110), .A3(new_n781), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n849), .A3(new_n844), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n845), .A2(new_n851), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n840), .A2(new_n843), .A3(new_n844), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n629), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n856), .ZN(G1333gat));
  INV_X1    g656(.A(KEYINPUT50), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n838), .A2(new_n839), .A3(new_n526), .ZN(new_n859));
  INV_X1    g658(.A(G71gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n769), .A2(G71gat), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n840), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n858), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n840), .A2(new_n862), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n865), .B(KEYINPUT50), .C1(new_n859), .C2(new_n860), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(G1334gat));
  NAND2_X1  g666(.A1(new_n840), .A2(new_n291), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g668(.A1(new_n785), .A2(new_n623), .A3(new_n796), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n809), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(G85gat), .B1(new_n871), .B2(new_n535), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n785), .A2(new_n623), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n781), .A2(new_n712), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n781), .A2(KEYINPUT51), .A3(new_n712), .A4(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n878), .A2(new_n676), .A3(new_n540), .A4(new_n744), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n872), .A2(new_n879), .ZN(G1336gat));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n876), .A2(new_n881), .A3(new_n877), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n874), .A2(KEYINPUT112), .A3(new_n875), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n796), .A2(new_n489), .A3(G92gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n775), .A2(new_n784), .A3(new_n753), .A4(new_n870), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n673), .A2(new_n675), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT52), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT52), .B1(new_n878), .B2(new_n884), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1337gat));
  OAI21_X1  g692(.A(G99gat), .B1(new_n871), .B2(new_n526), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n537), .A2(new_n744), .A3(new_n683), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n895), .B(KEYINPUT113), .Z(new_n896));
  NAND2_X1  g695(.A1(new_n878), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(G1338gat));
  NOR3_X1   g697(.A1(new_n796), .A2(G106gat), .A3(new_n532), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT114), .Z(new_n900));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n883), .A3(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n775), .A2(new_n784), .A3(new_n291), .A4(new_n870), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G106gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT53), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT53), .B1(new_n878), .B2(new_n899), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1339gat));
  INV_X1    g707(.A(KEYINPUT115), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n910), .B(new_n715), .C1(new_n729), .C2(new_n722), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n911), .B2(new_n742), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n909), .A3(new_n742), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n910), .B1(new_n727), .B2(new_n733), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n728), .B2(new_n731), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n915), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n914), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n917), .B(KEYINPUT55), .C1(new_n919), .C2(new_n912), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n917), .B1(new_n919), .B2(new_n912), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT55), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n739), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n623), .A2(new_n918), .A3(new_n922), .A4(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n602), .B1(new_n597), .B2(new_n601), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n604), .A2(new_n605), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n610), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n744), .A2(new_n619), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n712), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n925), .A2(new_n922), .A3(new_n918), .ZN(new_n932));
  INV_X1    g731(.A(new_n712), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n619), .A2(new_n929), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n669), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n713), .A2(new_n789), .A3(new_n796), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n535), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n546), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(new_n312), .A3(new_n751), .ZN(new_n940));
  INV_X1    g739(.A(new_n939), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n623), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n312), .B2(new_n942), .ZN(G1340gat));
  NOR2_X1   g742(.A1(new_n939), .A2(new_n796), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(new_n309), .ZN(G1341gat));
  NOR2_X1   g744(.A1(new_n939), .A2(new_n669), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(new_n301), .ZN(G1342gat));
  NOR2_X1   g746(.A1(new_n939), .A2(new_n933), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n317), .A2(new_n318), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n948), .A2(KEYINPUT56), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G134gat), .B1(new_n939), .B2(new_n933), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT56), .B1(new_n948), .B2(new_n950), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(G1343gat));
  AOI21_X1  g753(.A(new_n932), .B1(new_n625), .B2(new_n626), .ZN(new_n955));
  INV_X1    g754(.A(new_n930), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n933), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n935), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n785), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n937), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n291), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT57), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n526), .A2(new_n540), .A3(new_n489), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT117), .Z(new_n964));
  AOI21_X1  g763(.A(new_n532), .B1(new_n936), .B2(new_n937), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT57), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n962), .A2(new_n627), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G141gat), .ZN(new_n969));
  XOR2_X1   g768(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n970));
  NAND2_X1  g769(.A1(new_n526), .A2(new_n291), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n971), .A2(new_n753), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n938), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n751), .A2(G141gat), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT118), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n970), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n969), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n962), .A2(new_n623), .A3(new_n967), .ZN(new_n978));
  AOI22_X1  g777(.A1(new_n978), .A2(G141gat), .B1(new_n973), .B2(new_n975), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT58), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(G1344gat));
  INV_X1    g780(.A(G148gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n973), .A2(new_n982), .A3(new_n744), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT59), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G148gat), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n962), .A2(new_n967), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(new_n986), .B2(new_n744), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n714), .A2(new_n627), .A3(new_n744), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n966), .B(new_n291), .C1(new_n959), .C2(new_n988), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n930), .B1(new_n932), .B2(new_n789), .ZN(new_n990));
  AND4_X1   g789(.A1(new_n712), .A2(new_n925), .A3(new_n918), .A4(new_n922), .ZN(new_n991));
  INV_X1    g790(.A(new_n934), .ZN(new_n992));
  AOI22_X1  g791(.A1(new_n990), .A2(new_n933), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n937), .B1(new_n993), .B2(new_n785), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(new_n291), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(KEYINPUT57), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n964), .A2(new_n796), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n989), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n984), .B1(new_n998), .B2(G148gat), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n983), .B1(new_n987), .B2(new_n999), .ZN(G1345gat));
  NAND2_X1  g799(.A1(new_n962), .A2(new_n967), .ZN(new_n1001));
  OAI21_X1  g800(.A(G155gat), .B1(new_n1001), .B2(new_n669), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n973), .A2(new_n207), .A3(new_n785), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(G1346gat));
  NAND3_X1  g803(.A1(new_n973), .A2(new_n208), .A3(new_n712), .ZN(new_n1005));
  XNOR2_X1  g804(.A(new_n1005), .B(KEYINPUT120), .ZN(new_n1006));
  OAI21_X1  g805(.A(G162gat), .B1(new_n1001), .B2(new_n933), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(G1347gat));
  AOI21_X1  g807(.A(new_n540), .B1(new_n936), .B2(new_n937), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n769), .A2(new_n291), .A3(new_n489), .ZN(new_n1010));
  AND2_X1   g809(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1011), .A2(new_n407), .A3(new_n623), .ZN(new_n1012));
  XNOR2_X1  g811(.A(new_n1012), .B(KEYINPUT121), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n407), .B1(new_n1011), .B2(new_n627), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1014), .A2(KEYINPUT122), .ZN(new_n1015));
  OR2_X1    g814(.A1(new_n1014), .A2(KEYINPUT122), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(G1348gat));
  NAND2_X1  g816(.A1(new_n1011), .A2(new_n744), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(G176gat), .ZN(G1349gat));
  INV_X1    g818(.A(KEYINPUT125), .ZN(new_n1020));
  NAND4_X1  g819(.A1(new_n994), .A2(new_n535), .A3(new_n785), .A4(new_n1010), .ZN(new_n1021));
  AND2_X1   g820(.A1(new_n382), .A2(new_n384), .ZN(new_n1022));
  INV_X1    g821(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1023), .A2(KEYINPUT123), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g824(.A1(new_n404), .A2(new_n401), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1026), .B1(new_n1022), .B2(KEYINPUT123), .ZN(new_n1027));
  INV_X1    g826(.A(new_n1027), .ZN(new_n1028));
  NAND4_X1  g827(.A1(new_n1009), .A2(new_n785), .A3(new_n1010), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g828(.A(new_n1020), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g829(.A1(new_n1030), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1031));
  OR2_X1    g830(.A1(new_n1030), .A2(KEYINPUT124), .ZN(new_n1032));
  INV_X1    g831(.A(KEYINPUT60), .ZN(new_n1033));
  NAND2_X1  g832(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1034));
  AOI21_X1  g833(.A(new_n1033), .B1(new_n1034), .B2(KEYINPUT124), .ZN(new_n1035));
  AOI21_X1  g834(.A(new_n1031), .B1(new_n1032), .B2(new_n1035), .ZN(G1350gat));
  AOI21_X1  g835(.A(new_n377), .B1(new_n1011), .B2(new_n712), .ZN(new_n1037));
  OR2_X1    g836(.A1(new_n1037), .A2(KEYINPUT61), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n1037), .A2(KEYINPUT61), .ZN(new_n1039));
  NAND4_X1  g838(.A1(new_n1011), .A2(new_n378), .A3(new_n380), .A4(new_n712), .ZN(new_n1040));
  NAND3_X1  g839(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(G1351gat));
  NOR2_X1   g840(.A1(new_n971), .A2(new_n489), .ZN(new_n1042));
  AND2_X1   g841(.A1(new_n1009), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g842(.A(G197gat), .B1(new_n1043), .B2(new_n623), .ZN(new_n1044));
  AND2_X1   g843(.A1(new_n989), .A2(new_n996), .ZN(new_n1045));
  NOR3_X1   g844(.A1(new_n818), .A2(new_n540), .A3(new_n489), .ZN(new_n1046));
  OR2_X1    g845(.A1(new_n1046), .A2(KEYINPUT126), .ZN(new_n1047));
  NAND2_X1  g846(.A1(new_n1046), .A2(KEYINPUT126), .ZN(new_n1048));
  AND3_X1   g847(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g848(.A1(new_n751), .A2(new_n225), .ZN(new_n1050));
  AOI21_X1  g849(.A(new_n1044), .B1(new_n1049), .B2(new_n1050), .ZN(G1352gat));
  NAND4_X1  g850(.A1(new_n1045), .A2(new_n744), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1052));
  NAND2_X1  g851(.A1(new_n1052), .A2(G204gat), .ZN(new_n1053));
  NAND3_X1  g852(.A1(new_n1043), .A2(new_n226), .A3(new_n744), .ZN(new_n1054));
  NAND2_X1  g853(.A1(new_n1054), .A2(KEYINPUT62), .ZN(new_n1055));
  OR2_X1    g854(.A1(new_n1054), .A2(KEYINPUT62), .ZN(new_n1056));
  NAND3_X1  g855(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(G1353gat));
  NAND3_X1  g856(.A1(new_n1043), .A2(new_n230), .A3(new_n785), .ZN(new_n1058));
  NAND4_X1  g857(.A1(new_n989), .A2(new_n996), .A3(new_n785), .A4(new_n1046), .ZN(new_n1059));
  AND3_X1   g858(.A1(new_n1059), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1060));
  AOI21_X1  g859(.A(KEYINPUT63), .B1(new_n1059), .B2(G211gat), .ZN(new_n1061));
  OAI21_X1  g860(.A(new_n1058), .B1(new_n1060), .B2(new_n1061), .ZN(G1354gat));
  NAND3_X1  g861(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1063));
  OAI21_X1  g862(.A(G218gat), .B1(new_n1063), .B2(new_n933), .ZN(new_n1064));
  NAND3_X1  g863(.A1(new_n1043), .A2(new_n231), .A3(new_n712), .ZN(new_n1065));
  NAND2_X1  g864(.A1(new_n1064), .A2(new_n1065), .ZN(G1355gat));
endmodule


