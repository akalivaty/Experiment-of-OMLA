

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581;

  XOR2_X1 U323 ( .A(G78GAT), .B(G148GAT), .Z(n291) );
  XOR2_X1 U324 ( .A(n414), .B(n365), .Z(n292) );
  NAND2_X1 U325 ( .A1(n556), .A2(n569), .ZN(n496) );
  XNOR2_X1 U326 ( .A(n314), .B(KEYINPUT31), .ZN(n315) );
  XNOR2_X1 U327 ( .A(n387), .B(n315), .ZN(n319) );
  NOR2_X1 U328 ( .A1(n455), .A2(n575), .ZN(n456) );
  XNOR2_X1 U329 ( .A(n322), .B(n413), .ZN(n323) );
  XNOR2_X1 U330 ( .A(n324), .B(n323), .ZN(n325) );
  NOR2_X1 U331 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U332 ( .A1(n485), .A2(n459), .ZN(n460) );
  XOR2_X1 U333 ( .A(KEYINPUT41), .B(n502), .Z(n556) );
  XNOR2_X1 U334 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U335 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n448) );
  XOR2_X1 U336 ( .A(G141GAT), .B(G22GAT), .Z(n378) );
  XNOR2_X1 U337 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n293), .B(G8GAT), .ZN(n438) );
  XOR2_X1 U339 ( .A(n378), .B(n438), .Z(n295) );
  NAND2_X1 U340 ( .A1(G229GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U342 ( .A(n296), .B(KEYINPUT67), .Z(n300) );
  XOR2_X1 U343 ( .A(G29GAT), .B(KEYINPUT8), .Z(n298) );
  XNOR2_X1 U344 ( .A(KEYINPUT7), .B(KEYINPUT70), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n420) );
  XNOR2_X1 U346 ( .A(n420), .B(KEYINPUT30), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U348 ( .A(G197GAT), .B(G43GAT), .Z(n302) );
  XNOR2_X1 U349 ( .A(G50GAT), .B(G36GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U351 ( .A(n304), .B(n303), .Z(n312) );
  XOR2_X1 U352 ( .A(KEYINPUT68), .B(KEYINPUT66), .Z(n306) );
  XNOR2_X1 U353 ( .A(KEYINPUT69), .B(KEYINPUT72), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U355 ( .A(KEYINPUT29), .B(G113GAT), .Z(n308) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(G15GAT), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U359 ( .A(n312), .B(n311), .Z(n474) );
  INV_X1 U360 ( .A(n474), .ZN(n569) );
  XNOR2_X1 U361 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n291), .B(n313), .ZN(n387) );
  AND2_X1 U363 ( .A1(G230GAT), .A2(G233GAT), .ZN(n314) );
  XOR2_X1 U364 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n317) );
  XNOR2_X1 U365 ( .A(G176GAT), .B(KEYINPUT33), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n324) );
  XNOR2_X1 U368 ( .A(G99GAT), .B(G71GAT), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n320), .B(G120GAT), .ZN(n365) );
  XNOR2_X1 U370 ( .A(G204GAT), .B(G64GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n321), .B(KEYINPUT75), .ZN(n358) );
  XOR2_X1 U372 ( .A(n365), .B(n358), .Z(n322) );
  XOR2_X1 U373 ( .A(G85GAT), .B(G92GAT), .Z(n413) );
  XNOR2_X1 U374 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n429) );
  XNOR2_X1 U375 ( .A(n325), .B(n429), .ZN(n473) );
  NAND2_X1 U376 ( .A1(n569), .A2(n473), .ZN(n459) );
  XOR2_X1 U377 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n327) );
  XNOR2_X1 U378 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n332) );
  XNOR2_X1 U380 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n328), .B(KEYINPUT2), .ZN(n385) );
  XOR2_X1 U382 ( .A(G162GAT), .B(n385), .Z(n330) );
  XOR2_X1 U383 ( .A(G113GAT), .B(KEYINPUT0), .Z(n371) );
  XNOR2_X1 U384 ( .A(G29GAT), .B(n371), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n345) );
  XOR2_X1 U387 ( .A(G85GAT), .B(G148GAT), .Z(n334) );
  XNOR2_X1 U388 ( .A(G141GAT), .B(G134GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U390 ( .A(G57GAT), .B(G120GAT), .Z(n336) );
  XNOR2_X1 U391 ( .A(G1GAT), .B(G127GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U393 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U394 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n340) );
  NAND2_X1 U395 ( .A1(G225GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U397 ( .A(KEYINPUT89), .B(n341), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U399 ( .A(n345), .B(n344), .Z(n543) );
  INV_X1 U400 ( .A(n543), .ZN(n566) );
  XOR2_X1 U401 ( .A(G176GAT), .B(G183GAT), .Z(n347) );
  XNOR2_X1 U402 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U404 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n349) );
  XNOR2_X1 U405 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U407 ( .A(n351), .B(n350), .Z(n375) );
  XOR2_X1 U408 ( .A(KEYINPUT21), .B(G218GAT), .Z(n353) );
  XNOR2_X1 U409 ( .A(KEYINPUT86), .B(G211GAT), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U411 ( .A(G197GAT), .B(n354), .Z(n388) );
  XOR2_X1 U412 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n356) );
  XNOR2_X1 U413 ( .A(G8GAT), .B(G92GAT), .ZN(n355) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n388), .B(n357), .ZN(n362) );
  XOR2_X1 U416 ( .A(G36GAT), .B(KEYINPUT78), .Z(n417) );
  XOR2_X1 U417 ( .A(n417), .B(n358), .Z(n360) );
  NAND2_X1 U418 ( .A1(G226GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U421 ( .A(n375), .B(n363), .Z(n488) );
  XOR2_X1 U422 ( .A(KEYINPUT27), .B(n488), .Z(n398) );
  NOR2_X1 U423 ( .A1(n566), .A2(n398), .ZN(n364) );
  XOR2_X1 U424 ( .A(KEYINPUT94), .B(n364), .Z(n509) );
  XOR2_X1 U425 ( .A(G43GAT), .B(G134GAT), .Z(n414) );
  NAND2_X1 U426 ( .A1(G227GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n292), .B(n366), .ZN(n370) );
  XOR2_X1 U428 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n368) );
  XNOR2_X1 U429 ( .A(KEYINPUT82), .B(KEYINPUT81), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U431 ( .A(n370), .B(n369), .Z(n373) );
  XOR2_X1 U432 ( .A(G15GAT), .B(G127GAT), .Z(n430) );
  XNOR2_X1 U433 ( .A(n430), .B(n371), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U435 ( .A(n375), .B(n374), .Z(n549) );
  XOR2_X1 U436 ( .A(KEYINPUT85), .B(n549), .Z(n391) );
  XOR2_X1 U437 ( .A(G204GAT), .B(KEYINPUT24), .Z(n377) );
  XNOR2_X1 U438 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n382) );
  XOR2_X1 U440 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n380) );
  XOR2_X1 U441 ( .A(G50GAT), .B(G162GAT), .Z(n419) );
  XNOR2_X1 U442 ( .A(n378), .B(n419), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U444 ( .A(n382), .B(n381), .Z(n384) );
  NAND2_X1 U445 ( .A1(G228GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n384), .B(n383), .ZN(n386) );
  XOR2_X1 U447 ( .A(n386), .B(n385), .Z(n390) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n544) );
  XOR2_X1 U450 ( .A(n544), .B(KEYINPUT28), .Z(n469) );
  NAND2_X1 U451 ( .A1(n391), .A2(n469), .ZN(n392) );
  NOR2_X1 U452 ( .A1(n509), .A2(n392), .ZN(n403) );
  INV_X1 U453 ( .A(n488), .ZN(n540) );
  NOR2_X1 U454 ( .A1(n549), .A2(n540), .ZN(n393) );
  NOR2_X1 U455 ( .A1(n393), .A2(n544), .ZN(n394) );
  XOR2_X1 U456 ( .A(n394), .B(KEYINPUT25), .Z(n395) );
  XNOR2_X1 U457 ( .A(KEYINPUT96), .B(n395), .ZN(n400) );
  XOR2_X1 U458 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n397) );
  NAND2_X1 U459 ( .A1(n544), .A2(n549), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n397), .B(n396), .ZN(n568) );
  NOR2_X1 U461 ( .A1(n568), .A2(n398), .ZN(n399) );
  NOR2_X1 U462 ( .A1(n400), .A2(n399), .ZN(n401) );
  NOR2_X1 U463 ( .A1(n401), .A2(n543), .ZN(n402) );
  NOR2_X1 U464 ( .A1(n403), .A2(n402), .ZN(n455) );
  XOR2_X1 U465 ( .A(G106GAT), .B(G99GAT), .Z(n405) );
  NAND2_X1 U466 ( .A1(G232GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U468 ( .A(G190GAT), .B(n406), .ZN(n424) );
  XOR2_X1 U469 ( .A(KEYINPUT65), .B(KEYINPUT77), .Z(n408) );
  XNOR2_X1 U470 ( .A(G218GAT), .B(KEYINPUT76), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U472 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n410) );
  XNOR2_X1 U473 ( .A(KEYINPUT64), .B(KEYINPUT11), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U475 ( .A(n412), .B(n411), .Z(n416) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n418) );
  XOR2_X1 U478 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n560) );
  XOR2_X1 U482 ( .A(G155GAT), .B(G71GAT), .Z(n426) );
  XNOR2_X1 U483 ( .A(G22GAT), .B(G183GAT), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n442) );
  XOR2_X1 U485 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n428) );
  XNOR2_X1 U486 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n429), .B(G78GAT), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n430), .B(G211GAT), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U491 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U492 ( .A1(G231GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U494 ( .A(n437), .B(KEYINPUT14), .Z(n440) );
  XNOR2_X1 U495 ( .A(n438), .B(KEYINPUT15), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n575) );
  INV_X1 U498 ( .A(n575), .ZN(n443) );
  NOR2_X1 U499 ( .A1(n560), .A2(n443), .ZN(n444) );
  XOR2_X1 U500 ( .A(KEYINPUT16), .B(n444), .Z(n445) );
  NOR2_X1 U501 ( .A1(n455), .A2(n445), .ZN(n446) );
  XNOR2_X1 U502 ( .A(KEYINPUT97), .B(n446), .ZN(n475) );
  NOR2_X1 U503 ( .A1(n459), .A2(n475), .ZN(n453) );
  NAND2_X1 U504 ( .A1(n453), .A2(n543), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U506 ( .A(G1GAT), .B(n449), .Z(G1324GAT) );
  NAND2_X1 U507 ( .A1(n488), .A2(n453), .ZN(n450) );
  XNOR2_X1 U508 ( .A(G8GAT), .B(n450), .ZN(G1325GAT) );
  XOR2_X1 U509 ( .A(G15GAT), .B(KEYINPUT35), .Z(n452) );
  INV_X1 U510 ( .A(n549), .ZN(n510) );
  NAND2_X1 U511 ( .A1(n453), .A2(n510), .ZN(n451) );
  XNOR2_X1 U512 ( .A(n452), .B(n451), .ZN(G1326GAT) );
  INV_X1 U513 ( .A(n469), .ZN(n513) );
  NAND2_X1 U514 ( .A1(n513), .A2(n453), .ZN(n454) );
  XNOR2_X1 U515 ( .A(n454), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U516 ( .A(KEYINPUT36), .B(n560), .ZN(n577) );
  NAND2_X1 U517 ( .A1(n577), .A2(n456), .ZN(n457) );
  XOR2_X1 U518 ( .A(KEYINPUT100), .B(n457), .Z(n458) );
  XNOR2_X1 U519 ( .A(KEYINPUT37), .B(n458), .ZN(n485) );
  XOR2_X1 U520 ( .A(KEYINPUT38), .B(n460), .Z(n468) );
  NOR2_X1 U521 ( .A1(n566), .A2(n468), .ZN(n463) );
  XOR2_X1 U522 ( .A(G29GAT), .B(KEYINPUT99), .Z(n461) );
  XNOR2_X1 U523 ( .A(KEYINPUT39), .B(n461), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n463), .B(n462), .ZN(G1328GAT) );
  NOR2_X1 U525 ( .A1(n468), .A2(n540), .ZN(n464) );
  XOR2_X1 U526 ( .A(G36GAT), .B(n464), .Z(G1329GAT) );
  NOR2_X1 U527 ( .A1(n549), .A2(n468), .ZN(n466) );
  XNOR2_X1 U528 ( .A(KEYINPUT40), .B(KEYINPUT101), .ZN(n465) );
  XNOR2_X1 U529 ( .A(G43GAT), .B(n467), .ZN(G1330GAT) );
  XNOR2_X1 U530 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U533 ( .A(G50GAT), .B(n472), .ZN(G1331GAT) );
  XNOR2_X1 U534 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n477) );
  INV_X1 U535 ( .A(n473), .ZN(n502) );
  NAND2_X1 U536 ( .A1(n556), .A2(n474), .ZN(n484) );
  NOR2_X1 U537 ( .A1(n475), .A2(n484), .ZN(n481) );
  NAND2_X1 U538 ( .A1(n481), .A2(n543), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(G1332GAT) );
  NAND2_X1 U540 ( .A1(n481), .A2(n488), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n478), .B(KEYINPUT104), .ZN(n479) );
  XNOR2_X1 U542 ( .A(G64GAT), .B(n479), .ZN(G1333GAT) );
  NAND2_X1 U543 ( .A1(n510), .A2(n481), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n480), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U545 ( .A(G78GAT), .B(KEYINPUT43), .Z(n483) );
  NAND2_X1 U546 ( .A1(n481), .A2(n513), .ZN(n482) );
  XNOR2_X1 U547 ( .A(n483), .B(n482), .ZN(G1335GAT) );
  XOR2_X1 U548 ( .A(G85GAT), .B(KEYINPUT105), .Z(n487) );
  NOR2_X1 U549 ( .A1(n485), .A2(n484), .ZN(n492) );
  NAND2_X1 U550 ( .A1(n492), .A2(n543), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(G1336GAT) );
  NAND2_X1 U552 ( .A1(n492), .A2(n488), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n489), .B(KEYINPUT106), .ZN(n490) );
  XNOR2_X1 U554 ( .A(G92GAT), .B(n490), .ZN(G1337GAT) );
  NAND2_X1 U555 ( .A1(n510), .A2(n492), .ZN(n491) );
  XNOR2_X1 U556 ( .A(n491), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n494) );
  NAND2_X1 U558 ( .A1(n492), .A2(n513), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U560 ( .A(G106GAT), .B(n495), .ZN(G1339GAT) );
  XNOR2_X1 U561 ( .A(KEYINPUT109), .B(KEYINPUT48), .ZN(n508) );
  XNOR2_X1 U562 ( .A(n496), .B(KEYINPUT46), .ZN(n498) );
  NOR2_X1 U563 ( .A1(n560), .A2(n575), .ZN(n497) );
  AND2_X1 U564 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n499), .B(KEYINPUT47), .ZN(n506) );
  XOR2_X1 U566 ( .A(KEYINPUT45), .B(KEYINPUT108), .Z(n501) );
  NAND2_X1 U567 ( .A1(n575), .A2(n577), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n501), .B(n500), .ZN(n504) );
  NOR2_X1 U569 ( .A1(n569), .A2(n502), .ZN(n503) );
  NAND2_X1 U570 ( .A1(n504), .A2(n503), .ZN(n505) );
  NAND2_X1 U571 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n541) );
  NOR2_X1 U573 ( .A1(n509), .A2(n541), .ZN(n523) );
  NAND2_X1 U574 ( .A1(n523), .A2(n510), .ZN(n511) );
  XNOR2_X1 U575 ( .A(KEYINPUT110), .B(n511), .ZN(n512) );
  NOR2_X1 U576 ( .A1(n513), .A2(n512), .ZN(n520) );
  NAND2_X1 U577 ( .A1(n520), .A2(n569), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n514), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n516) );
  NAND2_X1 U580 ( .A1(n520), .A2(n556), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U582 ( .A(G120GAT), .B(n517), .Z(G1341GAT) );
  NAND2_X1 U583 ( .A1(n575), .A2(n520), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(KEYINPUT50), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G127GAT), .B(n519), .ZN(G1342GAT) );
  XOR2_X1 U586 ( .A(G134GAT), .B(KEYINPUT51), .Z(n522) );
  NAND2_X1 U587 ( .A1(n520), .A2(n560), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(G1343GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n526) );
  INV_X1 U590 ( .A(n523), .ZN(n524) );
  NOR2_X1 U591 ( .A1(n568), .A2(n524), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n536), .A2(n569), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G141GAT), .B(n527), .ZN(G1344GAT) );
  NAND2_X1 U595 ( .A1(n536), .A2(n556), .ZN(n533) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(KEYINPUT53), .Z(n529) );
  XNOR2_X1 U597 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n528) );
  XNOR2_X1 U598 ( .A(n529), .B(n528), .ZN(n531) );
  XOR2_X1 U599 ( .A(G148GAT), .B(KEYINPUT52), .Z(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(G1345GAT) );
  XOR2_X1 U602 ( .A(G155GAT), .B(KEYINPUT117), .Z(n535) );
  NAND2_X1 U603 ( .A1(n536), .A2(n575), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(G1346GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n538) );
  NAND2_X1 U606 ( .A1(n536), .A2(n560), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U608 ( .A(G162GAT), .B(n539), .ZN(G1347GAT) );
  XNOR2_X1 U609 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n552) );
  NOR2_X1 U610 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n542), .B(KEYINPUT54), .ZN(n565) );
  NOR2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  AND2_X1 U613 ( .A1(n565), .A2(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U616 ( .A(KEYINPUT121), .B(n550), .Z(n561) );
  NAND2_X1 U617 ( .A1(n569), .A2(n561), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n554) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U622 ( .A(KEYINPUT56), .B(n555), .Z(n558) );
  NAND2_X1 U623 ( .A1(n561), .A2(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  NAND2_X1 U625 ( .A1(n575), .A2(n561), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(n564), .ZN(G1351GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  NAND2_X1 U632 ( .A1(n565), .A2(n566), .ZN(n567) );
  NOR2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n578), .A2(n569), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n578), .A2(n502), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n578), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n580) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(G218GAT), .B(n581), .Z(G1355GAT) );
endmodule

