//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  AOI21_X1  g001(.A(KEYINPUT13), .B1(new_n187), .B2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G128), .B(G143), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G122), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G116), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G122), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n196), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n196), .B2(new_n199), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n192), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(new_n194), .B(KEYINPUT88), .ZN(new_n203));
  XNOR2_X1  g017(.A(new_n199), .B(KEYINPUT14), .ZN(new_n204));
  OAI21_X1  g018(.A(G107), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n196), .A2(new_n197), .A3(new_n199), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n191), .B(new_n189), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n208), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT9), .B(G234), .Z(new_n210));
  XNOR2_X1  g024(.A(new_n210), .B(KEYINPUT73), .ZN(new_n211));
  INV_X1    g025(.A(G953), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(G217), .A3(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n209), .A2(new_n213), .ZN(new_n215));
  AOI21_X1  g029(.A(G902), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G478), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n216), .A2(new_n218), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n212), .A2(G952), .ZN(new_n222));
  INV_X1    g036(.A(G234), .ZN(new_n223));
  INV_X1    g037(.A(G237), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  AOI211_X1 g041(.A(new_n227), .B(new_n212), .C1(G234), .C2(G237), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT21), .B(G898), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G475), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT16), .ZN(new_n233));
  INV_X1    g047(.A(G140), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(G125), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(G125), .ZN(new_n238));
  INV_X1    g052(.A(G125), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G140), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT16), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT68), .A4(G125), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n237), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n237), .A2(new_n241), .A3(G146), .A4(new_n242), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n224), .A2(new_n212), .A3(G214), .ZN(new_n248));
  INV_X1    g062(.A(G143), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G237), .A2(G953), .ZN(new_n251));
  AOI21_X1  g065(.A(G143), .B1(new_n251), .B2(G214), .ZN(new_n252));
  OAI21_X1  g066(.A(G131), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n248), .A2(new_n249), .ZN(new_n254));
  INV_X1    g068(.A(G131), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n251), .A2(G143), .A3(G214), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n255), .B1(new_n254), .B2(new_n256), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT86), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT17), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n259), .B2(KEYINPUT17), .ZN(new_n262));
  OAI221_X1 g076(.A(new_n247), .B1(KEYINPUT17), .B2(new_n258), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G113), .B(G122), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT85), .B(G104), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n250), .A2(new_n252), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT18), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n268), .B(KEYINPUT81), .C1(new_n269), .C2(new_n255), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT81), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n254), .A2(new_n256), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n257), .B(new_n271), .C1(new_n272), .C2(KEYINPUT18), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n238), .A2(new_n240), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT80), .B1(new_n275), .B2(G146), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(G146), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(KEYINPUT80), .A3(G146), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n278), .A2(new_n279), .B1(KEYINPUT18), .B2(new_n259), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n263), .A2(new_n267), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n267), .B1(new_n263), .B2(new_n281), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n232), .B1(new_n285), .B2(new_n227), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT20), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n250), .A2(new_n252), .A3(G131), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT82), .B1(new_n289), .B2(new_n259), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT82), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n253), .A2(new_n291), .A3(new_n257), .ZN(new_n292));
  INV_X1    g106(.A(new_n275), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT83), .B(KEYINPUT19), .Z(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT83), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n275), .B1(new_n296), .B2(KEYINPUT19), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n297), .A3(new_n244), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n290), .A2(new_n246), .A3(new_n292), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n281), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT84), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n281), .A2(new_n299), .A3(KEYINPUT84), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n266), .A3(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n304), .A2(KEYINPUT87), .A3(new_n282), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT87), .B1(new_n304), .B2(new_n282), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(G475), .A2(G902), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n288), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n288), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(new_n304), .B2(new_n282), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n231), .B(new_n287), .C1(new_n309), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n313));
  XNOR2_X1  g127(.A(G110), .B(G122), .ZN(new_n314));
  INV_X1    g128(.A(G104), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT3), .B1(new_n315), .B2(G107), .ZN(new_n316));
  AOI21_X1  g130(.A(G101), .B1(new_n315), .B2(G107), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n197), .A3(G104), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT74), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n316), .A2(new_n317), .A3(new_n319), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n315), .A2(G107), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n316), .A2(new_n319), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n325), .B1(new_n327), .B2(G101), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G113), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT2), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT2), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G113), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n198), .A2(G119), .ZN(new_n334));
  INV_X1    g148(.A(G119), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G116), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n331), .B(new_n333), .C1(new_n334), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n333), .ZN(new_n338));
  XNOR2_X1  g152(.A(G116), .B(G119), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n327), .A2(new_n325), .A3(G101), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n329), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G101), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n197), .A2(G104), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(new_n326), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n321), .B2(new_n323), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(KEYINPUT5), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n330), .B1(new_n334), .B2(new_n349), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n348), .A2(new_n350), .B1(new_n339), .B2(new_n338), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n314), .B1(new_n343), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n313), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n314), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n341), .A2(new_n342), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n324), .B2(new_n328), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n347), .A2(new_n351), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n343), .A2(new_n352), .A3(new_n314), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT6), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n360), .A2(new_n361), .A3(new_n313), .A4(KEYINPUT6), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n244), .A2(G143), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n249), .A2(G146), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT0), .B(G128), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT64), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n249), .B2(G146), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n244), .A2(KEYINPUT64), .A3(G143), .ZN(new_n374));
  NAND2_X1  g188(.A1(KEYINPUT0), .A2(G128), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n373), .A2(new_n374), .A3(new_n376), .A4(new_n368), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n377), .A2(KEYINPUT65), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(KEYINPUT65), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n371), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n366), .B1(new_n380), .B2(new_n239), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n373), .A2(new_n374), .A3(new_n382), .A4(new_n368), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n187), .B1(new_n367), .B2(KEYINPUT1), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n369), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G125), .ZN(new_n386));
  INV_X1    g200(.A(new_n371), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n377), .A2(KEYINPUT65), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n377), .A2(KEYINPUT65), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n386), .B1(new_n390), .B2(G125), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n381), .B1(new_n391), .B2(new_n366), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(G224), .A3(new_n212), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n212), .A2(G224), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n381), .B(new_n394), .C1(new_n391), .C2(new_n366), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n365), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G210), .B1(G237), .B2(G902), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT79), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n394), .A2(KEYINPUT7), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n391), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n314), .B(KEYINPUT8), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n347), .A2(new_n351), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n359), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n361), .A3(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n381), .B(new_n401), .C1(new_n391), .C2(new_n366), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n227), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n397), .A2(new_n400), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n400), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n363), .A2(new_n364), .B1(new_n393), .B2(new_n395), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(new_n409), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G214), .B1(G237), .B2(G902), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n211), .A2(new_n227), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n417), .A2(G221), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(KEYINPUT76), .B(G469), .Z(new_n420));
  INV_X1    g234(.A(KEYINPUT11), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n189), .B2(G137), .ZN(new_n422));
  INV_X1    g236(.A(G137), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT11), .A3(G134), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n189), .A2(G137), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G131), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n422), .A2(new_n424), .A3(new_n255), .A4(new_n425), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n373), .A2(new_n374), .A3(new_n368), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT75), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n431), .B(KEYINPUT1), .C1(new_n249), .C2(G146), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G128), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n431), .B1(new_n367), .B2(KEYINPUT1), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n383), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n347), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n347), .A2(new_n385), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n429), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT12), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n347), .A2(new_n436), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT10), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n385), .A2(KEYINPUT10), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n441), .A2(new_n442), .B1(new_n443), .B2(new_n347), .ZN(new_n444));
  INV_X1    g258(.A(new_n429), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n380), .A2(new_n329), .A3(new_n342), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT12), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n448), .B(new_n429), .C1(new_n437), .C2(new_n438), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G140), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n212), .A2(G227), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n440), .A2(new_n447), .A3(new_n449), .A4(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n441), .A2(new_n442), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n443), .A2(new_n347), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n446), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n429), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n453), .B1(new_n459), .B2(new_n447), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n227), .B(new_n420), .C1(new_n455), .C2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n440), .A2(new_n447), .A3(new_n449), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n452), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n447), .A3(new_n453), .ZN(new_n464));
  AOI21_X1  g278(.A(G902), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G469), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n415), .A2(new_n416), .A3(new_n419), .A4(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n312), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n429), .B(new_n387), .C1(new_n388), .C2(new_n389), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT30), .ZN(new_n471));
  INV_X1    g285(.A(new_n425), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n189), .A2(G137), .ZN(new_n473));
  OAI21_X1  g287(.A(G131), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n385), .A2(new_n428), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n470), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n471), .B1(new_n470), .B2(new_n475), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n341), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n341), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n470), .A2(new_n480), .A3(new_n475), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n251), .A2(G210), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT27), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT26), .B(G101), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n479), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n470), .A2(new_n480), .A3(new_n475), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n480), .B1(new_n470), .B2(new_n475), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT28), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT28), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n485), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n486), .B1(new_n492), .B2(KEYINPUT31), .ZN(new_n493));
  INV_X1    g307(.A(new_n478), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n476), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n487), .B1(new_n495), .B2(new_n341), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT31), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n485), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT66), .ZN(new_n500));
  NOR2_X1   g314(.A1(G472), .A2(G902), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT66), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n493), .A2(new_n502), .A3(new_n498), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n500), .A2(KEYINPUT32), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n489), .A2(new_n485), .A3(new_n491), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT29), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n496), .ZN(new_n508));
  INV_X1    g322(.A(new_n485), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n227), .B1(new_n505), .B2(new_n506), .ZN(new_n511));
  OAI21_X1  g325(.A(G472), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n493), .A2(new_n502), .A3(new_n498), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n502), .B1(new_n493), .B2(new_n498), .ZN(new_n514));
  INV_X1    g328(.A(new_n501), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n504), .B(new_n512), .C1(new_n516), .C2(KEYINPUT32), .ZN(new_n517));
  INV_X1    g331(.A(G217), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(G234), .B2(new_n227), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n335), .A2(G128), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n335), .A2(G128), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n520), .B(new_n521), .C1(new_n522), .C2(KEYINPUT23), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G110), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT24), .B(G110), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT67), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n187), .B2(G119), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n335), .A2(KEYINPUT67), .A3(G128), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n187), .A2(G119), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n524), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n247), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n525), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n523), .A2(G110), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n530), .A2(KEYINPUT69), .A3(new_n525), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT70), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n293), .A2(new_n244), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n246), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n539), .B1(new_n538), .B2(new_n541), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n532), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT72), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n532), .B(KEYINPUT72), .C1(new_n543), .C2(new_n544), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n212), .A2(G221), .A3(G234), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT71), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT22), .B(G137), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n547), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n545), .A2(new_n546), .A3(new_n552), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT25), .B1(new_n556), .B2(new_n227), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT25), .ZN(new_n558));
  AOI211_X1 g372(.A(new_n558), .B(G902), .C1(new_n554), .C2(new_n555), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n519), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n519), .A2(G902), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n469), .A2(new_n517), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(G101), .ZN(G3));
  AND4_X1   g379(.A1(new_n560), .A2(new_n562), .A3(new_n419), .A4(new_n467), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n500), .A2(new_n227), .A3(new_n503), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n516), .B1(G472), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n216), .A2(new_n217), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n217), .A2(new_n227), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n214), .A2(new_n215), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT33), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT90), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n575), .B1(new_n215), .B2(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n574), .B(new_n577), .Z(new_n578));
  AOI21_X1  g392(.A(new_n573), .B1(new_n578), .B2(G478), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT87), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n281), .A2(KEYINPUT84), .A3(new_n299), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT84), .B1(new_n281), .B2(new_n299), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n581), .A2(new_n582), .A3(new_n267), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n583), .B2(new_n283), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n304), .A2(KEYINPUT87), .A3(new_n282), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n308), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n311), .B1(new_n586), .B2(KEYINPUT20), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n579), .B1(new_n587), .B2(new_n286), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT89), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n399), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n399), .A2(new_n589), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n397), .A2(new_n410), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(KEYINPUT89), .B(new_n398), .C1(new_n413), .C2(new_n409), .ZN(new_n594));
  INV_X1    g408(.A(new_n230), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n593), .A2(new_n594), .A3(new_n595), .A4(new_n416), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n569), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT34), .B(G104), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G6));
  NAND2_X1  g414(.A1(new_n586), .A2(KEYINPUT20), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n584), .A2(new_n288), .A3(new_n308), .A4(new_n585), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n286), .B1(new_n219), .B2(new_n220), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n596), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n569), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT35), .B(G107), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G9));
  NOR2_X1   g423(.A1(new_n553), .A2(KEYINPUT36), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n545), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n561), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n560), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n469), .A2(new_n568), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT37), .B(G110), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT91), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n614), .B(new_n616), .ZN(G12));
  INV_X1    g431(.A(G900), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n226), .B1(new_n228), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n601), .B2(new_n602), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n620), .A2(KEYINPUT92), .A3(new_n604), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT92), .B1(new_n620), .B2(new_n604), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n560), .A2(new_n612), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n504), .A2(new_n512), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT32), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n624), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n593), .A2(new_n594), .A3(new_n416), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n467), .A2(new_n419), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n623), .A2(new_n629), .A3(KEYINPUT93), .A4(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT93), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n517), .A2(new_n613), .A3(new_n632), .ZN(new_n635));
  INV_X1    g449(.A(new_n619), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n603), .A2(new_n604), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT92), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n620), .A2(KEYINPUT92), .A3(new_n604), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n634), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  XNOR2_X1  g458(.A(new_n415), .B(KEYINPUT38), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n287), .B1(new_n309), .B2(new_n311), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n221), .A4(new_n416), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n516), .A2(KEYINPUT32), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n496), .A2(new_n509), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n487), .A2(new_n488), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n227), .B1(new_n651), .B2(new_n485), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n504), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n624), .B1(new_n648), .B2(new_n654), .ZN(new_n655));
  OR3_X1    g469(.A1(new_n647), .A2(new_n655), .A3(KEYINPUT94), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT94), .B1(new_n647), .B2(new_n655), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n619), .B(KEYINPUT39), .Z(new_n658));
  NAND3_X1  g472(.A1(new_n467), .A2(new_n419), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT40), .Z(new_n660));
  NAND3_X1  g474(.A1(new_n656), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G143), .ZN(G45));
  NAND3_X1  g476(.A1(new_n646), .A2(new_n579), .A3(new_n636), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n629), .A2(new_n632), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  INV_X1    g480(.A(new_n447), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n445), .B1(new_n444), .B2(new_n446), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n452), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(G902), .B1(new_n669), .B2(new_n454), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n461), .B(new_n419), .C1(new_n466), .C2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n597), .A2(new_n517), .A3(new_n563), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT41), .B(G113), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G15));
  NAND4_X1  g489(.A1(new_n606), .A2(new_n517), .A3(new_n563), .A4(new_n672), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G116), .ZN(G18));
  NOR4_X1   g491(.A1(new_n587), .A2(new_n286), .A3(new_n221), .A4(new_n230), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n630), .A2(new_n671), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n517), .A2(new_n678), .A3(new_n613), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  OAI211_X1 g495(.A(new_n221), .B(new_n595), .C1(new_n587), .C2(new_n286), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n515), .B1(new_n493), .B2(new_n498), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n567), .B2(G472), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n683), .A2(new_n563), .A3(new_n685), .A4(new_n679), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G122), .ZN(G24));
  NAND2_X1  g501(.A1(new_n567), .A2(G472), .ZN(new_n688));
  INV_X1    g502(.A(new_n684), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n624), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n664), .A3(new_n679), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT95), .B(G125), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G27));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n411), .A2(new_n414), .A3(new_n416), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT96), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n462), .A2(new_n697), .A3(new_n452), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n464), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n697), .B1(new_n462), .B2(new_n452), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n466), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n466), .A2(new_n227), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n461), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n419), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n696), .B1(new_n705), .B2(KEYINPUT97), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n702), .B1(new_n670), .B2(new_n420), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n463), .A2(KEYINPUT96), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(G469), .A3(new_n464), .A4(new_n698), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n418), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT97), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n517), .A2(new_n563), .A3(new_n706), .A4(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n695), .B1(new_n713), .B2(new_n663), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n560), .A2(new_n562), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n625), .B2(new_n628), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n705), .A2(KEYINPUT97), .ZN(new_n717));
  INV_X1    g531(.A(new_n696), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n717), .A2(new_n712), .A3(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n719), .A3(KEYINPUT42), .A4(new_n664), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G131), .ZN(G33));
  INV_X1    g536(.A(KEYINPUT98), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n621), .B2(new_n622), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n639), .A2(KEYINPUT98), .A3(new_n640), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n716), .A4(new_n719), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G134), .ZN(G36));
  AOI21_X1  g541(.A(KEYINPUT45), .B1(new_n463), .B2(new_n464), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n466), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n708), .A2(KEYINPUT45), .A3(new_n464), .A4(new_n698), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n703), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n461), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n419), .B(new_n658), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT99), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n287), .B(new_n579), .C1(new_n309), .C2(new_n311), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(KEYINPUT101), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n740), .B1(new_n742), .B2(KEYINPUT100), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n646), .A2(new_n579), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n740), .A2(KEYINPUT100), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n744), .A2(KEYINPUT101), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n568), .A2(new_n624), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n743), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n739), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n749), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n696), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G137), .ZN(G39));
  OAI21_X1  g569(.A(new_n419), .B1(new_n735), .B2(new_n736), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(KEYINPUT47), .B(new_n419), .C1(new_n735), .C2(new_n736), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR4_X1   g574(.A1(new_n663), .A2(new_n517), .A3(new_n563), .A4(new_n696), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G140), .ZN(G42));
  NOR2_X1   g577(.A1(G952), .A2(G953), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n665), .A2(new_n692), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n646), .A2(new_n221), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n630), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n636), .A3(new_n710), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(new_n655), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n765), .A2(new_n769), .A3(new_n643), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n765), .A2(new_n769), .A3(new_n643), .A4(KEYINPUT52), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n714), .A2(new_n720), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n691), .A2(new_n719), .A3(new_n664), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n631), .A2(new_n696), .A3(new_n286), .A4(new_n221), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n629), .A2(new_n620), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n726), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n287), .B(new_n221), .C1(new_n309), .C2(new_n311), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n415), .A2(new_n595), .A3(new_n416), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n566), .A3(new_n568), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(new_n680), .A3(new_n686), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n588), .A2(KEYINPUT104), .ZN(new_n786));
  INV_X1    g600(.A(new_n782), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT104), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n579), .B(new_n788), .C1(new_n587), .C2(new_n286), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT105), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT105), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n786), .A2(new_n792), .A3(new_n787), .A4(new_n789), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n569), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n785), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n673), .A2(new_n676), .A3(new_n564), .A4(new_n614), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT106), .B1(new_n780), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n721), .A2(new_n726), .A3(new_n776), .A4(new_n778), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n673), .A2(new_n564), .A3(new_n614), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n785), .A3(new_n794), .A4(new_n676), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT106), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n774), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT107), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n799), .A2(new_n801), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n774), .A2(KEYINPUT53), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n806), .A2(new_n807), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n780), .A2(new_n797), .A3(KEYINPUT106), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n802), .B1(new_n799), .B2(new_n801), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n812), .A2(new_n813), .B1(new_n772), .B2(new_n773), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n808), .B(new_n810), .C1(new_n814), .C2(KEYINPUT53), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT107), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n812), .A2(new_n813), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(KEYINPUT53), .A3(new_n774), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n808), .B1(new_n806), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n811), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n743), .A2(new_n746), .A3(new_n226), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n696), .A2(new_n671), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n821), .A2(new_n716), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n824));
  NOR2_X1   g638(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n648), .A2(new_n654), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n563), .A3(new_n226), .A4(new_n822), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT112), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n646), .A3(new_n579), .ZN(new_n830));
  INV_X1    g644(.A(new_n679), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n690), .A2(new_n715), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n821), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n830), .B(new_n222), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n826), .B(new_n834), .C1(new_n823), .C2(new_n824), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n821), .A2(new_n822), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n836), .A2(new_n624), .A3(new_n690), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n829), .A2(new_n744), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n829), .A2(KEYINPUT113), .A3(new_n744), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n461), .B1(new_n466), .B2(new_n670), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT103), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n844), .A2(KEYINPUT108), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(KEYINPUT108), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n845), .A2(new_n846), .A3(new_n419), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n760), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n696), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n645), .A2(new_n416), .A3(new_n671), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT109), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n850), .B(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT50), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT111), .B1(new_n853), .B2(KEYINPUT110), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n853), .A2(KEYINPUT111), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n832), .B(new_n821), .C1(new_n849), .C2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n854), .B1(new_n833), .B2(new_n852), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n842), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n842), .A2(new_n857), .A3(KEYINPUT51), .A4(new_n858), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n835), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n764), .B1(new_n820), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n563), .A2(new_n416), .A3(new_n419), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT102), .Z(new_n867));
  NOR2_X1   g681(.A1(new_n645), .A2(new_n741), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n844), .B(KEYINPUT49), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n867), .A2(new_n827), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT115), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n817), .A2(KEYINPUT53), .A3(new_n774), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT53), .B1(new_n817), .B2(new_n774), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(KEYINPUT107), .A3(new_n815), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n863), .B1(new_n877), .B2(new_n811), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n873), .B(new_n870), .C1(new_n878), .C2(new_n764), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n872), .A2(new_n879), .ZN(G75));
  NOR2_X1   g694(.A1(new_n212), .A2(G952), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n774), .A2(KEYINPUT53), .A3(new_n809), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n875), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n227), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n885), .B2(G210), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n396), .B(KEYINPUT117), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n365), .B(KEYINPUT116), .Z(new_n889));
  XOR2_X1   g703(.A(new_n888), .B(new_n889), .Z(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n882), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n886), .B2(new_n891), .ZN(G51));
  OAI21_X1  g707(.A(KEYINPUT54), .B1(new_n875), .B2(new_n883), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n895), .A3(new_n815), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n806), .A2(new_n810), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n702), .B(KEYINPUT57), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(new_n460), .B2(new_n455), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n885), .A2(new_n730), .A3(new_n729), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n881), .B1(new_n901), .B2(new_n902), .ZN(G54));
  NAND3_X1  g717(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n904));
  INV_X1    g718(.A(new_n307), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n881), .ZN(G60));
  XNOR2_X1  g722(.A(new_n578), .B(KEYINPUT119), .ZN(new_n909));
  INV_X1    g723(.A(new_n820), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n572), .B(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n909), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AND4_X1   g727(.A1(new_n898), .A2(new_n896), .A3(new_n909), .A4(new_n912), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n881), .A3(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT60), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n897), .A2(new_n611), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n884), .A2(new_n917), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n919), .B(new_n882), .C1(new_n920), .C2(new_n556), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(KEYINPUT121), .A3(KEYINPUT61), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT61), .B1(new_n921), .B2(KEYINPUT121), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(G66));
  INV_X1    g739(.A(new_n229), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n212), .B1(new_n926), .B2(G224), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n801), .B2(new_n212), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n889), .B1(G898), .B2(new_n212), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n928), .B(new_n929), .Z(G69));
  NAND2_X1  g744(.A1(G900), .A2(G953), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n762), .A2(new_n721), .A3(new_n726), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n665), .A2(new_n692), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n642), .B2(new_n633), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n739), .A2(new_n716), .A3(new_n767), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n932), .A2(new_n754), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n931), .B1(new_n936), .B2(G953), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n295), .A2(new_n297), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT122), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n495), .B(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n659), .A2(new_n696), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n786), .A2(new_n789), .ZN(new_n942));
  INV_X1    g756(.A(new_n781), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n716), .B(new_n941), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n762), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n751), .B2(new_n753), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n934), .A2(new_n661), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n934), .A2(new_n661), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n946), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n940), .A2(G953), .ZN(new_n952));
  AOI22_X1  g766(.A1(new_n937), .A2(new_n940), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n212), .B1(G227), .B2(G900), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G72));
  NAND4_X1  g769(.A1(new_n946), .A2(new_n797), .A3(new_n948), .A4(new_n950), .ZN(new_n956));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n649), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT123), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n962), .A3(new_n649), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n958), .B1(new_n936), .B2(new_n801), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n508), .A2(new_n485), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT124), .Z(new_n967));
  AOI21_X1  g781(.A(new_n881), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n806), .A2(new_n818), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n970));
  INV_X1    g784(.A(new_n958), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n966), .A2(new_n649), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n970), .B1(new_n969), .B2(new_n972), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n964), .B(new_n968), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n975), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n973), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n980), .A2(KEYINPUT126), .A3(new_n964), .A4(new_n968), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(new_n981), .ZN(G57));
endmodule


