//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1197,
    new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT66), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n461), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n466), .A2(new_n467), .A3(G137), .A4(new_n468), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n461), .A2(new_n464), .A3(new_n468), .A4(new_n465), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT67), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n460), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n463), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n465), .A2(new_n476), .A3(new_n477), .A4(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n465), .A2(new_n476), .A3(G125), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT65), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n468), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n475), .A2(new_n484), .ZN(G160));
  MUX2_X1   g060(.A(G100), .B(G112), .S(G2105), .Z(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2104), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT68), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n461), .A2(new_n464), .A3(G2105), .A4(new_n465), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  INV_X1    g066(.A(new_n470), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n488), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT69), .ZN(G162));
  MUX2_X1   g070(.A(G102), .B(G114), .S(G2105), .Z(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2104), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n489), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n470), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n465), .A2(new_n476), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n500), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n499), .B1(new_n501), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n513), .A2(new_n519), .ZN(G166));
  INV_X1    g095(.A(new_n515), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  INV_X1    g097(.A(new_n517), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G51), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n510), .A2(KEYINPUT70), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n525), .A2(new_n530), .A3(G63), .A4(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n522), .A2(new_n524), .A3(new_n531), .A4(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND3_X1  g110(.A1(new_n525), .A2(new_n530), .A3(G64), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n512), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n515), .A2(new_n539), .B1(new_n517), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  NAND3_X1  g117(.A1(new_n525), .A2(new_n530), .A3(G56), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n512), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n515), .A2(new_n546), .B1(new_n517), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  OAI21_X1  g130(.A(KEYINPUT73), .B1(new_n526), .B2(new_n527), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n508), .A2(new_n557), .A3(new_n509), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G65), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT72), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n512), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n521), .A2(G91), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n514), .A2(KEYINPUT71), .A3(G53), .A4(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  INV_X1    g145(.A(G166), .ZN(G303));
  AOI22_X1  g146(.A1(G87), .A2(new_n521), .B1(new_n523), .B2(G49), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n525), .A2(new_n530), .ZN(new_n574));
  INV_X1    g149(.A(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n573), .B1(new_n576), .B2(G651), .ZN(new_n577));
  AOI21_X1  g152(.A(G74), .B1(new_n525), .B2(new_n530), .ZN(new_n578));
  NOR3_X1   g153(.A1(new_n578), .A2(KEYINPUT74), .A3(new_n512), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n572), .B1(new_n577), .B2(new_n579), .ZN(G288));
  NAND3_X1  g155(.A1(new_n514), .A2(G48), .A3(G543), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT75), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n512), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n521), .A2(G86), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n574), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n512), .B1(new_n589), .B2(KEYINPUT76), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(KEYINPUT76), .B2(new_n589), .ZN(new_n591));
  AOI22_X1  g166(.A1(G85), .A2(new_n521), .B1(new_n523), .B2(G47), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G290));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(G301), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n510), .A2(new_n514), .A3(G92), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT10), .Z(new_n597));
  NAND2_X1  g172(.A1(new_n523), .A2(G54), .ZN(new_n598));
  XNOR2_X1  g173(.A(KEYINPUT77), .B(G66), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n559), .A2(new_n599), .B1(G79), .B2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n598), .B1(new_n600), .B2(new_n512), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n597), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n595), .B1(new_n605), .B2(new_n594), .ZN(G284));
  AOI21_X1  g181(.A(new_n595), .B1(new_n605), .B2(new_n594), .ZN(G321));
  NOR2_X1   g182(.A1(G286), .A2(new_n594), .ZN(new_n608));
  INV_X1    g183(.A(G299), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n594), .ZN(G297));
  AOI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n594), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  INV_X1    g188(.A(new_n549), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(new_n597), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n601), .A2(new_n602), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n601), .A2(new_n602), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n619), .A2(G559), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n615), .B1(new_n620), .B2(G868), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(KEYINPUT80), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(KEYINPUT80), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n624), .B(new_n625), .C1(G111), .C2(new_n468), .ZN(new_n626));
  INV_X1    g201(.A(G123), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n489), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n492), .B2(G135), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n502), .A2(new_n473), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n634), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n631), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT81), .ZN(G156));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT15), .B(G2435), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2427), .ZN(new_n643));
  INV_X1    g218(.A(G2430), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n646), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(G401));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT82), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT17), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n660), .B1(new_n657), .B2(new_n659), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n658), .B2(new_n659), .ZN(new_n663));
  INV_X1    g238(.A(new_n659), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n664), .A2(new_n660), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n661), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT83), .Z(new_n669));
  AND2_X1   g244(.A1(new_n669), .A2(G2096), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(G2096), .ZN(new_n671));
  INV_X1    g246(.A(G2100), .ZN(new_n672));
  OR3_X1    g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n672), .B1(new_n670), .B2(new_n671), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT84), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT20), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n677), .A2(new_n679), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n682), .A3(new_n680), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n684), .B(new_n687), .C1(new_n682), .C2(new_n686), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n690), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  NOR2_X1   g270(.A1(G16), .A2(G23), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT87), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(G288), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT33), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G6), .B(G305), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT32), .B(G1981), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(KEYINPUT88), .B1(new_n705), .B2(G16), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n705), .A2(KEYINPUT88), .A3(G16), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n706), .B(new_n707), .C1(G166), .C2(new_n698), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1971), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n701), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n698), .A2(G24), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT86), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G290), .B2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G1986), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  MUX2_X1   g294(.A(G95), .B(G107), .S(G2105), .Z(new_n720));
  AOI22_X1  g295(.A1(new_n492), .A2(G131), .B1(G2104), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT85), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n490), .A2(new_n722), .A3(G119), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n490), .B2(G119), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G25), .B(new_n725), .S(G29), .Z(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT35), .B(G1991), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n718), .A2(new_n719), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n712), .A2(new_n713), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT89), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(KEYINPUT36), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n730), .B(new_n732), .Z(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G33), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n473), .A2(G103), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT25), .Z(new_n737));
  AOI22_X1  g312(.A1(new_n502), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n468), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G139), .B2(new_n492), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT93), .Z(new_n741));
  OAI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n734), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G2072), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n734), .A2(G26), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  INV_X1    g320(.A(G104), .ZN(new_n746));
  AND3_X1   g321(.A1(new_n746), .A2(new_n468), .A3(KEYINPUT90), .ZN(new_n747));
  AOI21_X1  g322(.A(KEYINPUT90), .B1(new_n746), .B2(new_n468), .ZN(new_n748));
  OAI221_X1 g323(.A(G2104), .B1(G116), .B2(new_n468), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G128), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(new_n489), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G140), .B2(new_n492), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(new_n734), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT91), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n753), .A2(KEYINPUT91), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n745), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT92), .B(G2067), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G2084), .ZN(new_n760));
  AND2_X1   g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  NOR2_X1   g336(.A1(KEYINPUT24), .A2(G34), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n734), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G160), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n734), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n743), .B(new_n759), .C1(new_n760), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n698), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT23), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n609), .B2(new_n698), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n765), .A2(new_n760), .ZN(new_n771));
  NOR2_X1   g346(.A1(G29), .A2(G32), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT26), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n775), .A2(new_n776), .B1(G105), .B2(new_n473), .ZN(new_n777));
  INV_X1    g352(.A(G129), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n489), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n492), .B2(G141), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n772), .B1(new_n780), .B2(G29), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT94), .Z(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT27), .B(G1996), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n771), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n770), .B(new_n784), .C1(new_n782), .C2(new_n783), .ZN(new_n785));
  NOR2_X1   g360(.A1(G16), .A2(G19), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n549), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1341), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n698), .A2(G5), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G171), .B2(new_n698), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G1961), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT31), .B(G11), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT30), .B(G28), .Z(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(G29), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n629), .B2(G29), .ZN(new_n795));
  INV_X1    g370(.A(G2078), .ZN(new_n796));
  NAND2_X1  g371(.A1(G164), .A2(G29), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G27), .B2(G29), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n791), .B1(KEYINPUT95), .B2(new_n795), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  AOI211_X1 g374(.A(new_n788), .B(new_n799), .C1(new_n796), .C2(new_n798), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n757), .A2(new_n758), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n698), .A2(G21), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G168), .B2(new_n698), .ZN(new_n803));
  INV_X1    g378(.A(G1966), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  AOI22_X1  g380(.A1(KEYINPUT95), .A2(new_n795), .B1(new_n790), .B2(G1961), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n801), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n785), .A2(new_n800), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G29), .A2(G35), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G162), .B2(G29), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(G2090), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(G2090), .ZN(new_n814));
  NOR2_X1   g389(.A1(G4), .A2(G16), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n605), .B2(G16), .ZN(new_n816));
  INV_X1    g391(.A(G1348), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n766), .A2(new_n808), .A3(new_n813), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n733), .A2(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  NAND2_X1  g397(.A1(new_n605), .A2(G559), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT38), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n549), .A2(KEYINPUT97), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT97), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n545), .B2(new_n548), .ZN(new_n827));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  INV_X1    g403(.A(G67), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n574), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G651), .ZN(new_n831));
  AOI22_X1  g406(.A1(G93), .A2(new_n521), .B1(new_n523), .B2(G55), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n825), .A2(new_n827), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n614), .A2(new_n834), .A3(new_n826), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n824), .B(new_n836), .Z(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n834), .A2(G860), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n840), .A2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(new_n741), .B(new_n780), .ZN(new_n844));
  INV_X1    g419(.A(G130), .ZN(new_n845));
  AND2_X1   g420(.A1(G118), .A2(G2105), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G106), .B2(new_n468), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n489), .A2(new_n845), .B1(new_n847), .B2(new_n460), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n492), .B2(G142), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n634), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n725), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n501), .A2(new_n504), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT98), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n490), .A2(G126), .B1(G2104), .B2(new_n496), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n501), .A2(new_n855), .A3(new_n504), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(new_n752), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n851), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n844), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(G162), .B(new_n764), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n630), .ZN(new_n862));
  AOI21_X1  g437(.A(G37), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n862), .B2(new_n860), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g440(.A1(new_n834), .A2(G868), .ZN(new_n866));
  XNOR2_X1  g441(.A(G303), .B(G305), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n869));
  NAND2_X1  g444(.A1(G290), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n591), .A2(KEYINPUT101), .A3(new_n592), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(G288), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(G288), .B1(new_n870), .B2(new_n871), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n876), .A2(new_n872), .A3(new_n867), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n620), .B(new_n836), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n605), .A2(G299), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n619), .A2(new_n609), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT41), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n605), .B2(G299), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n619), .A2(KEYINPUT99), .A3(new_n609), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n880), .A4(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n879), .A2(new_n883), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n883), .A2(new_n888), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(KEYINPUT100), .A3(new_n879), .ZN(new_n893));
  INV_X1    g468(.A(new_n882), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n879), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n896), .A2(KEYINPUT42), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(KEYINPUT42), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n878), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n896), .A2(KEYINPUT42), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n875), .A2(new_n877), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(KEYINPUT42), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n866), .B1(new_n904), .B2(G868), .ZN(G295));
  AOI21_X1  g480(.A(new_n866), .B1(new_n904), .B2(G868), .ZN(G331));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g482(.A1(G171), .A2(KEYINPUT102), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n538), .B2(new_n541), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(G168), .A3(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n910), .A2(G168), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OR3_X1    g488(.A1(new_n836), .A2(new_n913), .A3(KEYINPUT104), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n836), .A2(new_n913), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n833), .A2(new_n911), .A3(new_n835), .A4(new_n912), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT104), .A3(new_n916), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n885), .A2(new_n880), .A3(new_n887), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n914), .B(new_n917), .C1(new_n918), .C2(new_n886), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n836), .A2(KEYINPUT103), .A3(new_n913), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT103), .B1(new_n836), .B2(new_n913), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n916), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n894), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n919), .A2(new_n886), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n901), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n894), .B1(new_n914), .B2(new_n917), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n892), .B2(new_n923), .ZN(new_n928));
  AOI21_X1  g503(.A(G37), .B1(new_n928), .B2(new_n878), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n907), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n916), .ZN(new_n931));
  INV_X1    g506(.A(new_n922), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n932), .B2(new_n920), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n883), .A2(new_n888), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n901), .B1(new_n935), .B2(new_n927), .ZN(new_n936));
  INV_X1    g511(.A(new_n927), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n878), .B(new_n937), .C1(new_n934), .C2(new_n933), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  AND4_X1   g514(.A1(new_n907), .A2(new_n936), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT44), .B1(new_n930), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT43), .B1(new_n926), .B2(new_n929), .ZN(new_n943));
  AND4_X1   g518(.A1(KEYINPUT43), .A2(new_n936), .A3(new_n938), .A4(new_n939), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n941), .A2(new_n945), .ZN(G397));
  XNOR2_X1  g521(.A(new_n752), .B(G2067), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n780), .B(G1996), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n856), .A2(new_n854), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n855), .B1(new_n501), .B2(new_n504), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n470), .A2(new_n471), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n956), .A2(new_n467), .B1(G101), .B2(new_n473), .ZN(new_n957));
  INV_X1    g532(.A(new_n483), .ZN(new_n958));
  OAI21_X1  g533(.A(G2105), .B1(new_n958), .B2(new_n480), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n957), .A2(new_n959), .A3(G40), .A4(new_n472), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n949), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT105), .Z(new_n963));
  INV_X1    g538(.A(new_n961), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n725), .B(new_n727), .Z(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(G290), .B(G1986), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n966), .B1(new_n961), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT116), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n953), .B2(new_n960), .ZN(new_n970));
  INV_X1    g545(.A(G40), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n475), .A2(new_n484), .A3(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n972), .A2(new_n857), .A3(KEYINPUT116), .A4(new_n950), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G2067), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(new_n950), .C1(new_n951), .C2(new_n952), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n972), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n817), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n976), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n619), .ZN(new_n983));
  OAI211_X1 g558(.A(KEYINPUT45), .B(new_n950), .C1(new_n951), .C2(new_n952), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n954), .B1(G164), .B2(G1384), .ZN(new_n985));
  XOR2_X1   g560(.A(KEYINPUT56), .B(G2072), .Z(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT114), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n984), .A2(new_n972), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n852), .A2(new_n854), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n950), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n960), .B1(new_n992), .B2(new_n954), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(KEYINPUT115), .A3(new_n984), .A4(new_n987), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n977), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n953), .B2(new_n977), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n972), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT110), .B(G1956), .Z(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G65), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n556), .B2(new_n558), .ZN(new_n1003));
  INV_X1    g578(.A(new_n562), .ZN(new_n1004));
  OAI21_X1  g579(.A(G651), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n568), .A2(new_n1005), .A3(KEYINPUT57), .A4(new_n564), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT113), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1005), .A2(new_n1009), .A3(new_n564), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n568), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1009), .B1(new_n1005), .B2(new_n564), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT112), .B(new_n1008), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT111), .B1(new_n563), .B2(new_n565), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(new_n568), .A3(new_n1010), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT112), .B1(new_n1016), .B2(new_n1008), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1007), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n983), .B1(new_n1001), .B2(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1018), .A2(KEYINPUT117), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1018), .A2(KEYINPUT117), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1001), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT58), .B(G1341), .Z(new_n1025));
  NAND3_X1  g600(.A1(new_n970), .A2(new_n973), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1996), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n993), .A2(new_n1027), .A3(new_n984), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n549), .B1(KEYINPUT118), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT119), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(KEYINPUT59), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1029), .A2(new_n1037), .A3(new_n1032), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1036), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1037), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1041));
  AOI211_X1 g616(.A(KEYINPUT119), .B(new_n1031), .C1(new_n1026), .C2(new_n1028), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  AND4_X1   g619(.A1(KEYINPUT61), .A2(new_n995), .A3(new_n1018), .A4(new_n1000), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n990), .A2(new_n994), .B1(new_n998), .B2(new_n999), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT61), .B1(new_n1046), .B2(new_n1018), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1001), .A2(new_n1019), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n976), .A2(KEYINPUT60), .A3(new_n619), .A4(new_n981), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n976), .A2(KEYINPUT60), .A3(new_n981), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n605), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1056), .A2(new_n1057), .B1(KEYINPUT60), .B2(new_n982), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1024), .B1(new_n1050), .B2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT123), .B(G1961), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n980), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G164), .A2(G1384), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n960), .B1(new_n1062), .B2(KEYINPUT45), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(G2078), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n955), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n984), .A2(new_n796), .A3(new_n972), .A4(new_n985), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT124), .B1(new_n1068), .B2(new_n1064), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(KEYINPUT124), .A3(new_n1064), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1067), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT125), .B1(new_n1072), .B2(G301), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1071), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n1069), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1074), .B(G171), .C1(new_n1076), .C2(new_n1067), .ZN(new_n1077));
  OR3_X1    g652(.A1(new_n958), .A2(new_n480), .A3(KEYINPUT126), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT126), .B1(new_n958), .B2(new_n480), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n468), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1065), .A2(G40), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1080), .A2(new_n475), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(new_n955), .A3(new_n984), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1061), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G301), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1073), .A2(new_n1077), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G303), .A2(G8), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n980), .A2(G2090), .ZN(new_n1093));
  AOI21_X1  g668(.A(G1971), .B1(new_n993), .B2(new_n984), .ZN(new_n1094));
  OAI211_X1 g669(.A(G8), .B(new_n1092), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT106), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n984), .A2(new_n972), .A3(new_n985), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1098), .A2(G1971), .B1(G2090), .B2(new_n980), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1099), .A2(KEYINPUT106), .A3(G8), .A4(new_n1092), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(G1976), .B(new_n572), .C1(new_n577), .C2(new_n579), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1102), .B(G8), .C1(new_n953), .C2(new_n960), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n576), .A2(new_n573), .A3(G651), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT74), .B1(new_n578), .B2(new_n512), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1976), .B1(new_n1106), .B2(new_n572), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1103), .A2(KEYINPUT52), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT107), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1103), .B2(KEYINPUT52), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(G305), .A2(G1981), .ZN(new_n1112));
  INV_X1    g687(.A(G1981), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n582), .A2(new_n1113), .A3(new_n584), .A4(new_n585), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT108), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT49), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g692(.A(KEYINPUT108), .B(KEYINPUT49), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1118));
  OAI21_X1  g693(.A(G8), .B1(new_n953), .B2(new_n960), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NOR4_X1   g695(.A1(new_n1103), .A2(new_n1109), .A3(new_n1107), .A4(KEYINPUT52), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1111), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1092), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n997), .A2(new_n972), .ZN(new_n1124));
  INV_X1    g699(.A(G2090), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1094), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G8), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1123), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1101), .A2(new_n1122), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(G1966), .B1(new_n955), .B2(new_n1063), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n978), .A2(new_n760), .A3(new_n972), .A4(new_n979), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(G8), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT121), .B1(new_n1133), .B2(G168), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT45), .B1(new_n857), .B2(new_n950), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n972), .B1(new_n992), .B2(new_n954), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n804), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1131), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1138), .A2(new_n1139), .A3(G8), .A4(G286), .ZN(new_n1140));
  NAND2_X1  g715(.A1(G286), .A2(G8), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1141), .A2(KEYINPUT122), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(KEYINPUT51), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1133), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1143), .ZN(new_n1145));
  OAI211_X1 g720(.A(G8), .B(new_n1145), .C1(new_n1138), .C2(G286), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1134), .A2(new_n1140), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1129), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1072), .A2(G301), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1149), .B(KEYINPUT54), .C1(G301), .C2(new_n1085), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1089), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1059), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1138), .A2(G8), .A3(G168), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1153), .B1(new_n1129), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1092), .B1(new_n1099), .B2(G8), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1156), .A2(new_n1154), .A3(new_n1153), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(new_n1101), .A3(new_n1122), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1129), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1134), .A2(new_n1140), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1162), .A2(KEYINPUT62), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT62), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1160), .B(new_n1161), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1122), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1119), .B(KEYINPUT109), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1120), .A2(G1976), .A3(G288), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1114), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1159), .A2(new_n1166), .A3(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n968), .B1(new_n1152), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n725), .A2(new_n727), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n963), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n752), .A2(new_n975), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n964), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OR3_X1    g753(.A1(new_n964), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT46), .B1(new_n964), .B2(G1996), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n947), .A2(new_n780), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1179), .A2(new_n1180), .B1(new_n961), .B2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT47), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n964), .A2(G1986), .A3(G290), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT127), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT48), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1185), .A2(KEYINPUT48), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1187), .A2(new_n966), .ZN(new_n1188));
  AOI211_X1 g763(.A(new_n1178), .B(new_n1183), .C1(new_n1186), .C2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1174), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g765(.A1(new_n860), .A2(new_n862), .ZN(new_n1192));
  AND2_X1   g766(.A1(new_n1192), .A2(new_n863), .ZN(new_n1193));
  NOR2_X1   g767(.A1(G401), .A2(new_n458), .ZN(new_n1194));
  NAND4_X1  g768(.A1(new_n673), .A2(new_n694), .A3(new_n674), .A4(new_n1194), .ZN(new_n1195));
  NOR4_X1   g769(.A1(new_n1193), .A2(new_n943), .A3(new_n944), .A4(new_n1195), .ZN(G308));
  NOR2_X1   g770(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1197));
  NOR2_X1   g771(.A1(new_n943), .A2(new_n944), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n1198), .ZN(G225));
endmodule


