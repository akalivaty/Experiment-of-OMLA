//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT21), .ZN(new_n209));
  XOR2_X1   g008(.A(G57gat), .B(G64gat), .Z(new_n210));
  AOI22_X1  g009(.A1(new_n210), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212));
  XOR2_X1   g011(.A(new_n212), .B(KEYINPUT96), .Z(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(KEYINPUT9), .ZN(new_n215));
  INV_X1    g014(.A(G71gat), .ZN(new_n216));
  INV_X1    g015(.A(G78gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n208), .B1(new_n209), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G231gat), .A2(G233gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G127gat), .B(G155gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(G211gat), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n225), .B(new_n227), .Z(new_n228));
  NAND2_X1  g027(.A1(new_n220), .A2(new_n209), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n229), .B(new_n230), .Z(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n228), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(G134gat), .B(G162gat), .Z(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT97), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n235), .B(new_n236), .Z(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G50gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G43gat), .ZN(new_n240));
  INV_X1    g039(.A(G43gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G50gat), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT15), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT90), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT15), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n241), .A2(G50gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n239), .A2(G43gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n243), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G29gat), .ZN(new_n250));
  INV_X1    g049(.A(G36gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT14), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT14), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(G29gat), .B2(G36gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(G29gat), .A2(G36gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT15), .B1(new_n240), .B2(new_n242), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(KEYINPUT90), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT91), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n249), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n261));
  OAI211_X1 g060(.A(KEYINPUT90), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT15), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n257), .B2(KEYINPUT90), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT91), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n243), .A2(new_n256), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n260), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT92), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT17), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(KEYINPUT92), .A3(KEYINPUT17), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G99gat), .B(G106gat), .Z(new_n274));
  NAND2_X1  g073(.A1(G85gat), .A2(G92gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT7), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G99gat), .A2(G106gat), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n278), .A2(KEYINPUT8), .ZN(new_n279));
  NOR2_X1   g078(.A1(G85gat), .A2(G92gat), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT99), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n280), .B1(KEYINPUT8), .B2(new_n278), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT99), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI211_X1 g083(.A(new_n274), .B(new_n277), .C1(new_n281), .C2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n274), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n284), .ZN(new_n287));
  INV_X1    g086(.A(new_n277), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n273), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(new_n286), .A3(new_n288), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n282), .A2(new_n283), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n279), .A2(KEYINPUT99), .A3(new_n280), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n274), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n268), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G190gat), .B(G218gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n299), .B(KEYINPUT100), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n238), .B1(new_n302), .B2(KEYINPUT101), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n298), .A2(new_n301), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n303), .B(new_n304), .C1(KEYINPUT101), .C2(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n302), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n237), .B(KEYINPUT98), .Z(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G230gat), .ZN(new_n310));
  INV_X1    g109(.A(G233gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n220), .B1(new_n289), .B2(new_n285), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n211), .A2(new_n213), .B1(new_n218), .B2(new_n210), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n314), .A3(new_n292), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT10), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n296), .A2(KEYINPUT10), .A3(new_n314), .A4(new_n292), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n312), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(new_n315), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n312), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G176gat), .B(G204gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT102), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(G120gat), .ZN(new_n326));
  INV_X1    g125(.A(G148gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n320), .A2(new_n322), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n233), .A2(new_n309), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT103), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT75), .B(G155gat), .ZN(new_n336));
  INV_X1    g135(.A(G162gat), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT2), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT74), .B1(new_n327), .B2(G141gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n340));
  INV_X1    g139(.A(G141gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(G148gat), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n339), .B(new_n342), .C1(new_n341), .C2(G148gat), .ZN(new_n343));
  INV_X1    g142(.A(G155gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(new_n337), .ZN(new_n345));
  NOR2_X1   g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n338), .B(new_n343), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(KEYINPUT73), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT2), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n341), .A2(G148gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n327), .A2(G141gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n348), .B(new_n352), .C1(new_n344), .C2(new_n337), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  XOR2_X1   g154(.A(G211gat), .B(G218gat), .Z(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G197gat), .B(G204gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(G211gat), .A2(G218gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT22), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(new_n361), .A3(new_n358), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n354), .B1(new_n355), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT70), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n356), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n357), .A2(new_n368), .A3(new_n362), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n347), .A2(new_n355), .A3(new_n353), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(new_n364), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G228gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(new_n311), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT79), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n379));
  OAI221_X1 g178(.A(new_n379), .B1(new_n376), .B2(new_n311), .C1(new_n367), .C2(new_n374), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT3), .B1(new_n372), .B2(new_n364), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n381), .A2(new_n354), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n370), .A2(KEYINPUT71), .A3(new_n371), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT71), .B1(new_n370), .B2(new_n371), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n373), .A2(new_n364), .ZN(new_n386));
  AOI211_X1 g185(.A(new_n376), .B(new_n311), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n378), .A2(new_n380), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT80), .B(G22gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(G78gat), .B(G106gat), .Z(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT31), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(new_n239), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n394));
  OAI21_X1  g193(.A(G22gat), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n387), .A2(new_n382), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n396), .A2(new_n397), .A3(new_n394), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n390), .B(new_n393), .C1(new_n395), .C2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n393), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n388), .A2(new_n389), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n388), .A2(new_n389), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT69), .ZN(new_n405));
  INV_X1    g204(.A(G190gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n222), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G169gat), .ZN(new_n408));
  INV_X1    g207(.A(G176gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT26), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT27), .B(G183gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(KEYINPUT28), .A3(new_n406), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT28), .B1(new_n414), .B2(new_n406), .ZN(new_n417));
  OAI221_X1 g216(.A(new_n412), .B1(new_n413), .B2(new_n410), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n407), .A2(KEYINPUT24), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n222), .A2(new_n406), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n407), .A2(KEYINPUT24), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT23), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n410), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT25), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n423), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n422), .A2(new_n426), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  OR3_X1    g229(.A1(new_n407), .A2(KEYINPUT65), .A3(KEYINPUT24), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT24), .B1(new_n407), .B2(KEYINPUT65), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n420), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n426), .A2(KEYINPUT64), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT64), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n424), .B2(new_n425), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n433), .A2(new_n428), .A3(new_n434), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT25), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n430), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT1), .ZN(new_n440));
  XNOR2_X1  g239(.A(G127gat), .B(G134gat), .ZN(new_n441));
  XOR2_X1   g240(.A(KEYINPUT67), .B(G120gat), .Z(new_n442));
  INV_X1    g241(.A(G113gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT68), .B(G113gat), .ZN(new_n445));
  INV_X1    g244(.A(G120gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n440), .B(new_n441), .C1(new_n444), .C2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(G127gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(G134gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT66), .B(G134gat), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(new_n449), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n443), .A2(new_n446), .ZN(new_n453));
  NAND2_X1  g252(.A1(G113gat), .A2(G120gat), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n440), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G227gat), .A2(G233gat), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n448), .A2(new_n456), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n430), .A2(new_n460), .A3(new_n438), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT34), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n458), .A2(KEYINPUT34), .A3(new_n459), .A4(new_n461), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(G15gat), .B(G43gat), .Z(new_n467));
  XNOR2_X1  g266(.A(G71gat), .B(G99gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n459), .B1(new_n458), .B2(new_n461), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(KEYINPUT33), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT32), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n461), .ZN(new_n475));
  INV_X1    g274(.A(new_n459), .ZN(new_n476));
  AOI221_X4 g275(.A(new_n472), .B1(KEYINPUT33), .B2(new_n469), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n405), .B(new_n466), .C1(new_n474), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n466), .A2(new_n405), .ZN(new_n479));
  INV_X1    g278(.A(new_n461), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n460), .B1(new_n430), .B2(new_n438), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT32), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n483), .B(new_n469), .C1(KEYINPUT33), .C2(new_n470), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n471), .A2(new_n473), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n464), .A2(KEYINPUT69), .A3(new_n465), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n479), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n404), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n438), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n418), .A2(new_n429), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT72), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(G226gat), .A2(G233gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n430), .A2(new_n494), .A3(new_n438), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n493), .A2(KEYINPUT29), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n439), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n372), .ZN(new_n500));
  INV_X1    g299(.A(new_n495), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n494), .B1(new_n430), .B2(new_n438), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n430), .A2(new_n493), .A3(new_n438), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n504), .A3(new_n385), .ZN(new_n505));
  XOR2_X1   g304(.A(G8gat), .B(G36gat), .Z(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(G64gat), .ZN(new_n507));
  INV_X1    g306(.A(G92gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n500), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n500), .A2(new_n505), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n509), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n500), .A2(new_n505), .A3(KEYINPUT30), .A4(new_n510), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n347), .A2(new_n353), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT3), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(new_n457), .A3(new_n373), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n448), .A2(new_n456), .A3(new_n347), .A4(new_n353), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(KEYINPUT4), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n521), .ZN(new_n523));
  XOR2_X1   g322(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT5), .ZN(new_n527));
  NAND2_X1  g326(.A1(G225gat), .A2(G233gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT77), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n460), .A2(new_n530), .A3(new_n354), .A4(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT77), .B1(new_n521), .B2(KEYINPUT4), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n532), .B(new_n533), .C1(new_n523), .C2(new_n524), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n534), .A2(new_n528), .A3(new_n520), .ZN(new_n535));
  OR3_X1    g334(.A1(new_n460), .A2(new_n354), .A3(KEYINPUT78), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n457), .A2(new_n518), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(KEYINPUT78), .A3(new_n521), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT5), .B1(new_n539), .B2(new_n528), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n529), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT0), .B(G57gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G85gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(G1gat), .B(G29gat), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n543), .B(new_n544), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT6), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n529), .B(new_n545), .C1(new_n535), .C2(new_n540), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n541), .A2(KEYINPUT6), .A3(new_n546), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n517), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n489), .A2(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(KEYINPUT86), .A2(KEYINPUT35), .ZN(new_n555));
  NAND2_X1  g354(.A1(KEYINPUT86), .A2(KEYINPUT35), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n554), .A2(KEYINPUT87), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT35), .B1(new_n489), .B2(new_n553), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n559), .B1(new_n551), .B2(new_n550), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n399), .A2(new_n403), .B1(new_n478), .B2(new_n487), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n560), .A2(new_n561), .A3(new_n555), .A4(new_n556), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT87), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n550), .A2(new_n551), .A3(new_n511), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n514), .A2(KEYINPUT37), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT38), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n499), .A2(new_n372), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n385), .B1(new_n503), .B2(new_n504), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT37), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n568), .A2(new_n569), .A3(new_n509), .A4(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n514), .A2(KEYINPUT37), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT38), .B1(new_n574), .B2(new_n567), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n510), .A2(KEYINPUT38), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n566), .A2(new_n573), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT83), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(new_n526), .B2(new_n528), .ZN(new_n579));
  INV_X1    g378(.A(new_n528), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n522), .A2(KEYINPUT83), .A3(new_n580), .A4(new_n525), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n539), .A2(new_n528), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n579), .A2(KEYINPUT39), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n545), .ZN(new_n584));
  XOR2_X1   g383(.A(KEYINPUT84), .B(KEYINPUT39), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(new_n579), .B2(new_n581), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n588), .A2(KEYINPUT40), .B1(new_n541), .B2(new_n546), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT85), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(new_n588), .B2(KEYINPUT40), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT40), .ZN(new_n592));
  OAI211_X1 g391(.A(KEYINPUT85), .B(new_n592), .C1(new_n584), .C2(new_n587), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n589), .A2(new_n591), .A3(new_n559), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n594), .A3(new_n404), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n399), .A2(KEYINPUT82), .A3(new_n403), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT82), .B1(new_n399), .B2(new_n403), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n553), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n488), .B(KEYINPUT36), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n565), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n268), .A2(KEYINPUT92), .A3(KEYINPUT17), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT17), .B1(new_n268), .B2(KEYINPUT92), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n208), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT93), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n208), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n268), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n604), .A2(KEYINPUT18), .A3(new_n607), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n268), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n606), .B(KEYINPUT13), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n609), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n616), .B1(new_n273), .B2(new_n208), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n607), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT18), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G113gat), .B(G141gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G169gat), .B(G197gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n615), .A2(new_n620), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n614), .A2(KEYINPUT94), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n610), .A2(new_n629), .A3(new_n613), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n620), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT95), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n626), .B(KEYINPUT89), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n631), .B2(new_n634), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n627), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n335), .A2(new_n601), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n552), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g440(.A1(new_n638), .A2(new_n559), .ZN(new_n642));
  NAND2_X1  g441(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n643));
  OR2_X1    g442(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(KEYINPUT42), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(KEYINPUT42), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n647), .B(new_n648), .C1(new_n207), .C2(new_n642), .ZN(G1325gat));
  AOI21_X1  g448(.A(G15gat), .B1(new_n638), .B2(new_n488), .ZN(new_n650));
  INV_X1    g449(.A(new_n599), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n638), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n650), .B1(G15gat), .B2(new_n652), .ZN(G1326gat));
  NOR2_X1   g452(.A1(new_n596), .A2(new_n597), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT43), .B(G22gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1327gat));
  INV_X1    g457(.A(new_n309), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n565), .B2(new_n600), .ZN(new_n660));
  INV_X1    g459(.A(new_n233), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n332), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n660), .A2(new_n637), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n250), .A3(new_n639), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT45), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n601), .A2(new_n309), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n660), .B2(new_n669), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n610), .A2(new_n629), .A3(new_n613), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n629), .B1(new_n610), .B2(new_n613), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT18), .B1(new_n617), .B2(new_n607), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT95), .B1(new_n674), .B2(new_n633), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT104), .B1(new_n677), .B2(new_n627), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n679));
  INV_X1    g478(.A(new_n627), .ZN(new_n680));
  AOI211_X1 g479(.A(new_n679), .B(new_n680), .C1(new_n675), .C2(new_n676), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n670), .A2(new_n683), .A3(new_n662), .ZN(new_n684));
  OAI21_X1  g483(.A(G29gat), .B1(new_n684), .B2(new_n552), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n665), .A2(new_n685), .ZN(G1328gat));
  NAND3_X1  g485(.A1(new_n663), .A2(new_n251), .A3(new_n559), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT46), .Z(new_n688));
  OAI21_X1  g487(.A(G36gat), .B1(new_n684), .B2(new_n517), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1329gat));
  OAI21_X1  g489(.A(G43gat), .B1(new_n684), .B2(new_n599), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n663), .A2(new_n241), .A3(new_n488), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(KEYINPUT47), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT107), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n692), .B(KEYINPUT106), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n695), .A2(new_n691), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(KEYINPUT47), .B2(new_n696), .ZN(G1330gat));
  NAND3_X1  g496(.A1(new_n663), .A2(new_n239), .A3(new_n655), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n684), .A2(new_n404), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n699), .A2(KEYINPUT109), .ZN(new_n700));
  OAI21_X1  g499(.A(G50gat), .B1(new_n699), .B2(KEYINPUT109), .ZN(new_n701));
  OAI211_X1 g500(.A(KEYINPUT48), .B(new_n698), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G50gat), .B1(new_n684), .B2(new_n654), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n703), .A2(new_n698), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(G1331gat));
  NOR2_X1   g505(.A1(new_n233), .A2(new_n309), .ZN(new_n707));
  INV_X1    g506(.A(new_n332), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n683), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n601), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n710), .A2(KEYINPUT110), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(KEYINPUT110), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n639), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g515(.A1(new_n713), .A2(new_n517), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  AND2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n717), .B2(new_n718), .ZN(G1333gat));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n714), .A2(G71gat), .A3(new_n651), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724));
  INV_X1    g523(.A(new_n488), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n216), .B1(new_n713), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n724), .B1(new_n723), .B2(new_n726), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n722), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n729), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(KEYINPUT50), .A3(new_n727), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(G1334gat));
  NOR2_X1   g532(.A1(new_n713), .A2(new_n654), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(new_n217), .ZN(G1335gat));
  AOI21_X1  g534(.A(new_n669), .B1(new_n601), .B2(new_n309), .ZN(new_n736));
  AOI211_X1 g535(.A(new_n659), .B(new_n666), .C1(new_n565), .C2(new_n600), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n233), .B(new_n709), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT112), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n670), .A2(new_n740), .A3(new_n233), .A4(new_n709), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n552), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(G85gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n660), .A2(new_n233), .A3(new_n682), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n332), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n639), .A2(new_n743), .ZN(new_n748));
  OAI22_X1  g547(.A1(new_n742), .A2(new_n743), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT113), .ZN(G1336gat));
  NAND2_X1  g549(.A1(new_n739), .A2(new_n741), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n508), .B1(new_n751), .B2(new_n559), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n744), .A2(KEYINPUT114), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n745), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n744), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n332), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n559), .A2(new_n508), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT52), .B1(new_n752), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  OAI21_X1  g559(.A(G92gat), .B1(new_n738), .B2(new_n517), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n760), .B(new_n761), .C1(new_n747), .C2(new_n757), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(G1337gat));
  AOI21_X1  g562(.A(new_n599), .B1(new_n739), .B2(new_n741), .ZN(new_n764));
  INV_X1    g563(.A(G99gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n488), .A2(new_n765), .ZN(new_n766));
  OAI22_X1  g565(.A1(new_n764), .A2(new_n765), .B1(new_n747), .B2(new_n766), .ZN(G1338gat));
  NOR3_X1   g566(.A1(new_n404), .A2(G106gat), .A3(new_n708), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n746), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  OAI21_X1  g569(.A(G106gat), .B1(new_n738), .B2(new_n404), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n755), .A3(new_n768), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n654), .B1(new_n739), .B2(new_n741), .ZN(new_n774));
  INV_X1    g573(.A(G106gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n776), .A2(KEYINPUT115), .A3(KEYINPUT53), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT115), .B1(new_n776), .B2(KEYINPUT53), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n772), .B1(new_n777), .B2(new_n778), .ZN(G1339gat));
  NAND2_X1  g578(.A1(new_n682), .A2(new_n333), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n317), .A2(new_n318), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  INV_X1    g581(.A(new_n312), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n317), .A2(new_n318), .A3(new_n312), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT54), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n328), .B(new_n784), .C1(new_n786), .C2(new_n319), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n331), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n788), .B2(new_n787), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n617), .A2(new_n607), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n611), .A2(new_n612), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n625), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n627), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n309), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n678), .B2(new_n681), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n332), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n796), .B1(new_n799), .B2(new_n659), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n780), .B1(new_n800), .B2(new_n661), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(new_n654), .A3(new_n488), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n680), .B1(new_n675), .B2(new_n676), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n639), .A2(new_n517), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n801), .A2(new_n639), .A3(new_n517), .A4(new_n561), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n682), .A2(new_n445), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n805), .A2(new_n443), .B1(new_n806), .B2(new_n807), .ZN(G1340gat));
  NOR3_X1   g607(.A1(new_n802), .A2(new_n708), .A3(new_n804), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n708), .A2(new_n442), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n809), .A2(new_n446), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT116), .Z(G1341gat));
  OR4_X1    g611(.A1(new_n449), .A2(new_n802), .A3(new_n233), .A4(new_n804), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n449), .B1(new_n806), .B2(new_n233), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n814), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(G1342gat));
  NOR3_X1   g617(.A1(new_n806), .A2(new_n451), .A3(new_n659), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT56), .ZN(new_n820));
  INV_X1    g619(.A(G134gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n802), .A2(new_n659), .A3(new_n804), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(G1343gat));
  INV_X1    g622(.A(new_n790), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n637), .A2(new_n679), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n677), .A2(KEYINPUT104), .A3(new_n627), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n798), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n659), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n661), .B1(new_n829), .B2(new_n795), .ZN(new_n830));
  INV_X1    g629(.A(new_n780), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n404), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n651), .A2(new_n804), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(G141gat), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT58), .B1(new_n836), .B2(new_n637), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n832), .B2(new_n404), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841));
  XOR2_X1   g640(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n842));
  AND3_X1   g641(.A1(new_n787), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n841), .B1(new_n787), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n840), .B1(new_n845), .B2(new_n789), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n787), .A2(new_n842), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT119), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n787), .A2(new_n841), .A3(new_n842), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n789), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(KEYINPUT120), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n846), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n798), .B1(new_n803), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n796), .B1(new_n854), .B2(new_n659), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT121), .B1(new_n855), .B2(new_n661), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT120), .B1(new_n850), .B2(new_n851), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n840), .B(new_n789), .C1(new_n848), .C2(new_n849), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n828), .B1(new_n859), .B2(new_n637), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n795), .B1(new_n860), .B2(new_n309), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n233), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n856), .A2(new_n863), .A3(new_n780), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(KEYINPUT57), .A3(new_n655), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n864), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n655), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n839), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n869), .A2(new_n637), .A3(new_n834), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n837), .B1(new_n870), .B2(new_n341), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n683), .A3(new_n834), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n872), .A2(G141gat), .B1(new_n637), .B2(new_n836), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(G1344gat));
  INV_X1    g674(.A(new_n404), .ZN(new_n876));
  OAI211_X1 g675(.A(KEYINPUT57), .B(new_n876), .C1(new_n830), .C2(new_n831), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n801), .A2(KEYINPUT123), .A3(KEYINPUT57), .A4(new_n876), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n335), .A2(new_n803), .B1(new_n233), .B2(new_n861), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n838), .B1(new_n881), .B2(new_n654), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n834), .A2(new_n332), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n884), .A2(G148gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n833), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n869), .A2(new_n332), .A3(new_n834), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT59), .B1(new_n891), .B2(G148gat), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT124), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(G148gat), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n883), .B2(new_n885), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n897), .A2(G148gat), .B1(new_n833), .B2(new_n888), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n893), .A2(new_n900), .ZN(G1345gat));
  NAND3_X1  g700(.A1(new_n869), .A2(new_n661), .A3(new_n834), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n835), .A2(new_n233), .ZN(new_n903));
  MUX2_X1   g702(.A(new_n902), .B(new_n903), .S(new_n336), .Z(G1346gat));
  NAND4_X1  g703(.A1(new_n869), .A2(G162gat), .A3(new_n309), .A4(new_n834), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n337), .B1(new_n835), .B2(new_n659), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(G1347gat));
  AOI21_X1  g706(.A(KEYINPUT125), .B1(new_n561), .B2(new_n559), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n832), .A2(new_n639), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n561), .A2(KEYINPUT125), .A3(new_n559), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n408), .A3(new_n683), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n552), .A2(new_n559), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n802), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G169gat), .B1(new_n916), .B2(new_n803), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n917), .ZN(G1348gat));
  AOI21_X1  g717(.A(G176gat), .B1(new_n912), .B2(new_n332), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n916), .A2(new_n409), .A3(new_n708), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(G1349gat));
  OAI21_X1  g720(.A(G183gat), .B1(new_n916), .B2(new_n233), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n661), .A2(new_n414), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n911), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g724(.A1(new_n912), .A2(new_n406), .A3(new_n309), .ZN(new_n926));
  OAI21_X1  g725(.A(G190gat), .B1(new_n916), .B2(new_n659), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n927), .A2(KEYINPUT61), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(KEYINPUT61), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(G1351gat));
  NOR2_X1   g729(.A1(new_n651), .A2(new_n914), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n883), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n803), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n833), .A2(new_n931), .ZN(new_n935));
  OR3_X1    g734(.A1(new_n935), .A2(G197gat), .A3(new_n682), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n934), .B1(new_n933), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(new_n938), .ZN(G1352gat));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n940), .B1(new_n932), .B2(new_n708), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n883), .A2(KEYINPUT127), .A3(new_n332), .A4(new_n931), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(G204gat), .A3(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n935), .A2(G204gat), .A3(new_n708), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT62), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1353gat));
  OR3_X1    g745(.A1(new_n935), .A2(G211gat), .A3(new_n233), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n883), .A2(new_n661), .A3(new_n931), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1354gat));
  OAI21_X1  g750(.A(G218gat), .B1(new_n932), .B2(new_n659), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n659), .A2(G218gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n935), .B2(new_n953), .ZN(G1355gat));
endmodule


