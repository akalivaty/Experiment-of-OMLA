//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1112,
    new_n1113, new_n1114, new_n1115;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT64), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT65), .Z(G319));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(KEYINPUT66), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n470), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  OR2_X1    g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(G2104), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT68), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n465), .B1(new_n466), .B2(KEYINPUT67), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n475), .A2(G101), .B1(G137), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT72), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n476), .A2(new_n478), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(G2105), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n486), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(new_n472), .A3(new_n489), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT71), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(new_n494), .B2(G136), .ZN(G162));
  INV_X1    g070(.A(G102), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n474), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n487), .A2(G126), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(new_n466), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n497), .B1(new_n500), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  AOI211_X1 g079(.A(new_n503), .B(new_n504), .C1(new_n479), .C2(G138), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n477), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT3), .B1(new_n477), .B2(G2104), .ZN(new_n507));
  OAI211_X1 g082(.A(G138), .B(new_n472), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT73), .B1(new_n508), .B2(KEYINPUT4), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT4), .A2(G2105), .ZN(new_n511));
  NOR3_X1   g086(.A1(new_n462), .A2(new_n463), .A3(new_n461), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT66), .B1(new_n467), .B2(new_n468), .ZN(new_n513));
  OAI211_X1 g088(.A(G138), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT74), .ZN(new_n515));
  INV_X1    g090(.A(G138), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n516), .B1(new_n464), .B2(new_n469), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(new_n518), .A3(new_n511), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n502), .B1(new_n510), .B2(new_n520), .ZN(G164));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT6), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT75), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n522), .A2(KEYINPUT6), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT76), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT5), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n527), .B1(new_n531), .B2(KEYINPUT77), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n533), .A2(KEYINPUT5), .A3(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G62), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT78), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G75), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n527), .ZN(new_n540));
  INV_X1    g115(.A(new_n535), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n526), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n540), .A2(G651), .B1(G88), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n530), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(G166));
  NAND2_X1  g120(.A1(new_n542), .A2(G89), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n528), .A2(G51), .ZN(new_n547));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT7), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n535), .B(new_n551), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n552), .A2(G63), .A3(G651), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(G168));
  NAND2_X1  g129(.A1(new_n528), .A2(G52), .ZN(new_n555));
  INV_X1    g130(.A(G90), .ZN(new_n556));
  INV_X1    g131(.A(new_n542), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n552), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n522), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n558), .A2(new_n560), .ZN(G171));
  AND2_X1   g136(.A1(new_n542), .A2(G81), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n552), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n522), .ZN(new_n564));
  AOI211_X1 g139(.A(new_n562), .B(new_n564), .C1(G43), .C2(new_n528), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(new_n528), .A2(G53), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n542), .A2(G91), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n535), .A2(G65), .ZN(new_n575));
  AND2_X1   g150(.A1(G78), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n573), .A2(new_n574), .A3(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  OR2_X1    g155(.A1(new_n544), .A2(KEYINPUT80), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n544), .A2(KEYINPUT80), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G303));
  AOI22_X1  g158(.A1(G49), .A2(new_n528), .B1(new_n542), .B2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n552), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT81), .Z(G288));
  NAND2_X1  g162(.A1(new_n542), .A2(G86), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n528), .A2(G48), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n535), .A2(G61), .ZN(new_n590));
  AND2_X1   g165(.A1(G73), .A2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n588), .A2(new_n589), .A3(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n552), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n522), .ZN(new_n595));
  AOI22_X1  g170(.A1(G47), .A2(new_n528), .B1(new_n542), .B2(G85), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OR3_X1    g175(.A1(new_n557), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n541), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n528), .A2(G54), .B1(G651), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT10), .B1(new_n557), .B2(new_n600), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n601), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT82), .Z(new_n608));
  OAI21_X1  g183(.A(new_n599), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n599), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G299), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G280));
  XOR2_X1   g188(.A(G280), .B(KEYINPUT83), .Z(G297));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G860), .ZN(G148));
  NOR2_X1   g191(.A1(new_n565), .A2(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n608), .A2(new_n615), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT84), .Z(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n475), .A2(new_n470), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n490), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G123), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(KEYINPUT85), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(KEYINPUT85), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n630), .B(new_n631), .C1(G111), .C2(new_n472), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(new_n494), .B2(G135), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n626), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT86), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT87), .B(KEYINPUT16), .Z(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  AND2_X1   g225(.A1(new_n650), .A2(G14), .ZN(G401));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT88), .Z(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(new_n654), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n654), .B(KEYINPUT17), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n659), .B(new_n656), .C1(new_n653), .C2(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n653), .A2(new_n660), .A3(new_n655), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2096), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n625), .ZN(G227));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n676), .B(new_n677), .C1(new_n675), .C2(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n682), .B(new_n685), .ZN(G229));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G25), .ZN(new_n688));
  AOI22_X1  g263(.A1(new_n494), .A2(G131), .B1(G119), .B2(new_n627), .ZN(new_n689));
  OR2_X1    g264(.A1(G95), .A2(G2105), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n690), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT91), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT92), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n688), .B1(new_n694), .B2(new_n687), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT93), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT35), .B(G1991), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n698), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT94), .B(G16), .Z(new_n701));
  MUX2_X1   g276(.A(G290), .B(G24), .S(new_n701), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1986), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n701), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1971), .ZN(new_n706));
  MUX2_X1   g281(.A(G23), .B(new_n586), .S(G16), .Z(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT33), .B(G1976), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n707), .B(new_n708), .Z(new_n709));
  MUX2_X1   g284(.A(G6), .B(G305), .S(G16), .Z(new_n710));
  XOR2_X1   g285(.A(KEYINPUT32), .B(G1981), .Z(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  NOR3_X1   g287(.A1(new_n706), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT34), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n703), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n699), .A2(new_n700), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT95), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n713), .A2(new_n714), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(KEYINPUT95), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT96), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n722), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n720), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G35), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT101), .B1(new_n727), .B2(G29), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n727), .A2(KEYINPUT101), .A3(G29), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n728), .B(new_n729), .C1(G162), .C2(new_n687), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT29), .B(G2090), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n717), .A2(new_n723), .A3(new_n718), .A4(new_n719), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n701), .A2(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n565), .B2(new_n701), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1341), .Z(new_n736));
  NAND2_X1  g311(.A1(G299), .A2(G16), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n701), .A2(G20), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT102), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT23), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G1956), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G2078), .ZN(new_n744));
  NOR2_X1   g319(.A1(G164), .A2(new_n687), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G27), .B2(new_n687), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n736), .B(new_n743), .C1(new_n744), .C2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G4), .ZN(new_n748));
  MUX2_X1   g323(.A(new_n748), .B(new_n608), .S(G16), .Z(new_n749));
  INV_X1    g324(.A(G1348), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n747), .B(new_n751), .C1(new_n744), .C2(new_n746), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT100), .B(G11), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT31), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n634), .A2(G29), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT99), .ZN(new_n756));
  NAND2_X1  g331(.A1(G168), .A2(G16), .ZN(new_n757));
  OR2_X1    g332(.A1(G16), .A2(G21), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n756), .B2(new_n757), .ZN(new_n760));
  INV_X1    g335(.A(G1966), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G28), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n764), .A2(new_n765), .A3(new_n687), .ZN(new_n766));
  NOR2_X1   g341(.A1(G5), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G171), .B2(G16), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G1961), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(G1961), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n762), .A2(new_n766), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G2084), .ZN(new_n772));
  INV_X1    g347(.A(G34), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT24), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n773), .B2(KEYINPUT24), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT97), .Z(new_n776));
  AOI22_X1  g351(.A1(G160), .A2(G29), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n771), .B1(new_n772), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n752), .A2(new_n754), .A3(new_n755), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n687), .A2(G33), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n470), .A2(G127), .ZN(new_n782));
  NAND2_X1  g357(.A1(G115), .A2(G2104), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n472), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n494), .B2(G139), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n781), .B1(new_n789), .B2(new_n687), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G2072), .Z(new_n791));
  OR2_X1    g366(.A1(G29), .A2(G32), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT26), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n494), .B2(G141), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n475), .A2(G105), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n627), .A2(G129), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n792), .B1(new_n798), .B2(new_n687), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT27), .B(G1996), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n777), .A2(G2084), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n791), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT98), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n780), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n726), .A2(new_n732), .A3(new_n733), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n799), .A2(new_n800), .ZN(new_n806));
  AOI21_X1  g381(.A(KEYINPUT28), .B1(new_n687), .B2(G26), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n687), .A2(G26), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n627), .A2(G128), .ZN(new_n809));
  OR2_X1    g384(.A1(G104), .A2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n810), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n494), .B2(G140), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n808), .B1(new_n813), .B2(new_n687), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n807), .B1(new_n814), .B2(KEYINPUT28), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G2067), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n805), .A2(new_n806), .A3(new_n817), .ZN(G311));
  AND3_X1   g393(.A1(new_n726), .A2(new_n733), .A3(new_n804), .ZN(new_n819));
  INV_X1    g394(.A(new_n806), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n819), .A2(new_n820), .A3(new_n816), .A4(new_n732), .ZN(G150));
  AOI22_X1  g396(.A1(new_n552), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(new_n522), .ZN(new_n823));
  AOI22_X1  g398(.A1(G55), .A2(new_n528), .B1(new_n542), .B2(G93), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT104), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  MUX2_X1   g403(.A(new_n826), .B(new_n825), .S(new_n565), .Z(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n608), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n831), .B(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n828), .B1(new_n835), .B2(G860), .ZN(G145));
  INV_X1    g411(.A(KEYINPUT107), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n788), .B(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n789), .A2(new_n837), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n798), .B(new_n813), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT106), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n520), .A2(new_n510), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n841), .B1(new_n520), .B2(new_n510), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n501), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n840), .B(new_n844), .ZN(new_n845));
  MUX2_X1   g420(.A(new_n838), .B(new_n839), .S(new_n845), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n494), .A2(G142), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n627), .A2(G130), .ZN(new_n848));
  NOR2_X1   g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(new_n472), .B2(G118), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n623), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n694), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n846), .A2(new_n853), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n482), .B(new_n634), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G162), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  OR3_X1    g433(.A1(new_n854), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n854), .B2(new_n855), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g438(.A1(new_n826), .A2(new_n611), .ZN(new_n864));
  XNOR2_X1  g439(.A(G299), .B(new_n607), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT41), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n829), .B(new_n618), .ZN(new_n868));
  MUX2_X1   g443(.A(new_n866), .B(new_n867), .S(new_n868), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT42), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n586), .B(G305), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G290), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G166), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n870), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n864), .B1(new_n875), .B2(new_n611), .ZN(G295));
  OAI21_X1  g451(.A(new_n864), .B1(new_n875), .B2(new_n611), .ZN(G331));
  XOR2_X1   g452(.A(G171), .B(G168), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n829), .B(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n879), .A2(new_n865), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n866), .ZN(new_n881));
  OR3_X1    g456(.A1(new_n880), .A2(new_n881), .A3(new_n874), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n874), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n860), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT43), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n882), .A2(new_n886), .A3(new_n860), .A4(new_n883), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(KEYINPUT44), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n889), .A3(new_n887), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n884), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n892), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT109), .B(G1384), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n844), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n481), .A2(G40), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n894), .B1(new_n901), .B2(G1996), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n813), .B(G2067), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n900), .B1(new_n904), .B2(new_n798), .ZN(new_n905));
  INV_X1    g480(.A(G1996), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(KEYINPUT46), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT47), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n694), .A2(new_n698), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n798), .A2(G1996), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n798), .A2(G1996), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n903), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G2067), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(new_n915), .B2(new_n813), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n909), .B1(new_n901), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n694), .B(new_n697), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT111), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n900), .B1(new_n919), .B2(new_n913), .ZN(new_n920));
  OR2_X1    g495(.A1(G290), .A2(G1986), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n901), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n922), .B(KEYINPUT48), .Z(new_n923));
  AOI21_X1  g498(.A(new_n917), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT127), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT63), .ZN(new_n926));
  INV_X1    g501(.A(G8), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n581), .B2(new_n582), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT55), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI211_X1 g505(.A(KEYINPUT55), .B(new_n927), .C1(new_n581), .C2(new_n582), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT113), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n928), .A2(new_n929), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT113), .B1(new_n935), .B2(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n899), .ZN(new_n938));
  NOR2_X1   g513(.A1(G164), .A2(G1384), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n942));
  AND4_X1   g517(.A1(new_n518), .A2(new_n470), .A3(G138), .A4(new_n511), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n518), .B1(new_n517), .B2(new_n511), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n503), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n508), .A2(KEYINPUT73), .A3(KEYINPUT4), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT106), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n520), .A2(new_n510), .A3(new_n841), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n502), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n942), .B1(new_n952), .B2(G1384), .ZN(new_n953));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n844), .A2(KEYINPUT112), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n941), .B1(new_n956), .B2(new_n940), .ZN(new_n957));
  INV_X1    g532(.A(G2090), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n844), .A2(KEYINPUT45), .A3(new_n895), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n960), .A2(new_n938), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n897), .B1(G164), .B2(G1384), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1971), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n927), .B1(new_n959), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n937), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n965), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n953), .A2(new_n955), .A3(KEYINPUT50), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n899), .B1(new_n939), .B2(new_n940), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n969), .A2(new_n958), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(G8), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n935), .B2(new_n931), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n956), .A2(new_n938), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(G8), .ZN(new_n975));
  XNOR2_X1  g550(.A(G305), .B(G1981), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT49), .Z(new_n977));
  OR2_X1    g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1976), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n586), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT52), .B1(new_n975), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT52), .B1(G288), .B2(new_n979), .ZN(new_n982));
  INV_X1    g557(.A(new_n980), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n974), .A3(G8), .A4(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n967), .A2(new_n973), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT114), .B1(new_n957), .B2(new_n772), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT50), .B1(new_n953), .B2(new_n955), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n990));
  NOR4_X1   g565(.A1(new_n989), .A2(new_n990), .A3(G2084), .A4(new_n941), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n953), .A2(new_n955), .A3(new_n897), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n899), .B1(new_n939), .B2(KEYINPUT45), .ZN(new_n993));
  AOI21_X1  g568(.A(G1966), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n988), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n995), .A2(new_n927), .A3(G286), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n926), .B1(new_n987), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT115), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n966), .B1(new_n930), .B2(new_n932), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(new_n926), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n985), .B1(new_n937), .B2(new_n966), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1001), .A2(new_n1002), .A3(KEYINPUT116), .A4(new_n996), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n996), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1007), .B(new_n926), .C1(new_n987), .C2(new_n997), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n999), .A2(new_n1003), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G305), .A2(G1981), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G288), .A2(G1976), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n977), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(new_n975), .ZN(new_n1013));
  INV_X1    g588(.A(new_n967), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1014), .B2(new_n986), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G286), .A2(G8), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT123), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1017), .B(new_n1020), .C1(new_n995), .C2(new_n927), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT51), .B1(new_n995), .B2(new_n1020), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n956), .A2(new_n940), .ZN(new_n1023));
  INV_X1    g598(.A(new_n941), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n772), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n990), .ZN(new_n1026));
  INV_X1    g601(.A(new_n994), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n957), .A2(KEYINPUT114), .A3(new_n772), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1019), .B1(new_n1029), .B2(G8), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1021), .B1(new_n1022), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT124), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT124), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1021), .B(new_n1033), .C1(new_n1022), .C2(new_n1030), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n974), .A2(KEYINPUT119), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n956), .A2(new_n1037), .A3(new_n938), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n915), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n750), .B1(new_n989), .B2(new_n941), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1956), .B1(new_n969), .B2(new_n970), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT118), .B(G2072), .Z(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT56), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n961), .A2(new_n962), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G299), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT57), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1043), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1041), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1049), .B(KEYINPUT120), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1051), .A2(new_n608), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1039), .A2(KEYINPUT60), .A3(new_n1040), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(new_n608), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1049), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1046), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(new_n1042), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT61), .B1(new_n1059), .B2(new_n1050), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1050), .A2(KEYINPUT122), .A3(KEYINPUT61), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT122), .B1(new_n1050), .B2(KEYINPUT61), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT60), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1041), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(new_n608), .A3(new_n1055), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1061), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n961), .A2(new_n906), .A3(new_n962), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT58), .B(G1341), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n565), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT59), .B(new_n565), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1054), .B1(new_n1068), .B2(new_n1078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n957), .A2(G1961), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n992), .A2(new_n993), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n744), .A2(KEYINPUT53), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(KEYINPUT125), .ZN(new_n1084));
  INV_X1    g659(.A(new_n963), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT53), .B1(new_n1085), .B2(new_n744), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(G171), .B(KEYINPUT54), .Z(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n961), .A2(KEYINPUT53), .A3(new_n744), .A4(new_n898), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1086), .B1(KEYINPUT126), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1089), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1092), .A2(KEYINPUT126), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1093), .A2(new_n1080), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1035), .A2(new_n1079), .A3(new_n1090), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1032), .A2(new_n1098), .A3(new_n1034), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(G171), .A3(new_n1088), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1098), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n987), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1016), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT110), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n921), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(G290), .A2(G1986), .ZN(new_n1107));
  XOR2_X1   g682(.A(new_n1106), .B(new_n1107), .Z(new_n1108));
  OAI21_X1  g683(.A(new_n920), .B1(new_n901), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n925), .B1(new_n1104), .B2(new_n1109), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g685(.A(G229), .ZN(new_n1112));
  NOR2_X1   g686(.A1(G401), .A2(G227), .ZN(new_n1113));
  NAND4_X1  g687(.A1(new_n890), .A2(new_n1112), .A3(new_n891), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g688(.A1(new_n862), .A2(G319), .ZN(new_n1115));
  NOR2_X1   g689(.A1(new_n1114), .A2(new_n1115), .ZN(G308));
  OR2_X1    g690(.A1(new_n1114), .A2(new_n1115), .ZN(G225));
endmodule


