

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831;

  XNOR2_X1 U377 ( .A(n356), .B(n655), .ZN(n808) );
  XNOR2_X1 U378 ( .A(n633), .B(n551), .ZN(n636) );
  AND2_X1 U379 ( .A1(n489), .A2(n675), .ZN(n679) );
  INV_X1 U380 ( .A(n505), .ZN(n358) );
  NOR2_X1 U381 ( .A1(n668), .A2(n753), .ZN(n662) );
  BUF_X1 U382 ( .A(G143), .Z(n355) );
  XNOR2_X1 U383 ( .A(n502), .B(G122), .ZN(n607) );
  NOR2_X2 U384 ( .A1(n774), .A2(n772), .ZN(n499) );
  XNOR2_X2 U385 ( .A(n682), .B(n681), .ZN(n774) );
  NAND2_X1 U386 ( .A1(n405), .A2(n403), .ZN(n356) );
  XNOR2_X1 U387 ( .A(n357), .B(n687), .ZN(n694) );
  NAND2_X1 U388 ( .A1(n729), .A2(n685), .ZN(n357) );
  NAND2_X1 U389 ( .A1(n456), .A2(n454), .ZN(n453) );
  XNOR2_X2 U390 ( .A(n515), .B(n564), .ZN(n626) );
  XNOR2_X2 U391 ( .A(n670), .B(n498), .ZN(n471) );
  XNOR2_X2 U392 ( .A(n386), .B(n541), .ZN(n531) );
  NOR2_X2 U393 ( .A1(n676), .A2(n677), .ZN(n678) );
  XNOR2_X1 U394 ( .A(n597), .B(n596), .ZN(n799) );
  NOR2_X1 U395 ( .A1(G953), .A2(G237), .ZN(n608) );
  NAND2_X2 U396 ( .A1(n411), .A2(n410), .ZN(n705) );
  NOR2_X1 U397 ( .A1(n684), .A2(n683), .ZN(n729) );
  XNOR2_X1 U398 ( .A(n679), .B(KEYINPUT107), .ZN(n684) );
  NOR2_X1 U399 ( .A1(n772), .A2(n439), .ZN(n438) );
  BUF_X1 U400 ( .A(n756), .Z(n501) );
  INV_X1 U401 ( .A(KEYINPUT36), .ZN(n666) );
  INV_X1 U402 ( .A(KEYINPUT38), .ZN(n360) );
  INV_X2 U403 ( .A(G137), .ZN(n513) );
  NAND2_X2 U404 ( .A1(n705), .A2(n747), .ZN(n412) );
  AND2_X1 U405 ( .A1(n431), .A2(n430), .ZN(n391) );
  AND2_X1 U406 ( .A1(n421), .A2(n419), .ZN(n418) );
  AND2_X1 U407 ( .A1(n390), .A2(n389), .ZN(n387) );
  AND2_X1 U408 ( .A1(n451), .A2(n368), .ZN(n425) );
  NAND2_X1 U409 ( .A1(n667), .A2(n501), .ZN(n740) );
  OR2_X1 U410 ( .A1(n778), .A2(n448), .ZN(n456) );
  XNOR2_X1 U411 ( .A(n494), .B(n666), .ZN(n667) );
  AND2_X1 U412 ( .A1(n455), .A2(n640), .ZN(n454) );
  XNOR2_X1 U413 ( .A(n487), .B(n638), .ZN(n778) );
  NAND2_X1 U414 ( .A1(n358), .A2(n438), .ZN(n633) );
  NOR2_X1 U415 ( .A1(n649), .A2(n441), .ZN(n487) );
  XNOR2_X1 U416 ( .A(n544), .B(n606), .ZN(n505) );
  XNOR2_X1 U417 ( .A(n497), .B(KEYINPUT6), .ZN(n441) );
  NOR2_X1 U418 ( .A1(n683), .A2(n605), .ZN(n544) );
  XNOR2_X1 U419 ( .A(n672), .B(n495), .ZN(n731) );
  XNOR2_X1 U420 ( .A(n545), .B(n604), .ZN(n683) );
  XNOR2_X1 U421 ( .A(n569), .B(n813), .ZN(n794) );
  XNOR2_X1 U422 ( .A(n571), .B(KEYINPUT25), .ZN(n572) );
  XNOR2_X1 U423 ( .A(n543), .B(G101), .ZN(n576) );
  XNOR2_X1 U424 ( .A(G116), .B(G107), .ZN(n503) );
  XOR2_X1 U425 ( .A(G146), .B(G125), .Z(n590) );
  INV_X1 U426 ( .A(KEYINPUT22), .ZN(n551) );
  BUF_X1 U427 ( .A(n393), .Z(n359) );
  NOR2_X2 U428 ( .A1(G902), .A2(n792), .ZN(n629) );
  XNOR2_X1 U429 ( .A(n665), .B(n360), .ZN(n680) );
  INV_X1 U430 ( .A(n665), .ZN(n698) );
  NAND2_X1 U431 ( .A1(n359), .A2(n434), .ZN(n361) );
  NAND2_X1 U432 ( .A1(n393), .A2(n434), .ZN(n691) );
  BUF_X1 U433 ( .A(n704), .Z(n362) );
  XNOR2_X2 U434 ( .A(n816), .B(G146), .ZN(n577) );
  XNOR2_X2 U435 ( .A(n588), .B(n369), .ZN(n816) );
  NAND2_X1 U436 ( .A1(n536), .A2(n535), .ZN(n410) );
  OR2_X1 U437 ( .A1(n366), .A2(n540), .ZN(n535) );
  NAND2_X1 U438 ( .A1(n415), .A2(n413), .ZN(n419) );
  NAND2_X1 U439 ( .A1(n423), .A2(n422), .ZN(n421) );
  XNOR2_X1 U440 ( .A(n802), .B(n426), .ZN(n598) );
  INV_X1 U441 ( .A(n576), .ZN(n426) );
  INV_X1 U442 ( .A(KEYINPUT64), .ZN(n493) );
  NOR2_X1 U443 ( .A1(n467), .A2(n798), .ZN(n466) );
  NOR2_X1 U444 ( .A1(n548), .A2(G475), .ZN(n467) );
  NAND2_X1 U445 ( .A1(n482), .A2(n365), .ZN(n480) );
  OR2_X1 U446 ( .A1(n710), .A2(G210), .ZN(n481) );
  NAND2_X1 U447 ( .A1(n538), .A2(n432), .ZN(n747) );
  INV_X1 U448 ( .A(KEYINPUT2), .ZN(n433) );
  INV_X1 U449 ( .A(KEYINPUT102), .ZN(n496) );
  INV_X1 U450 ( .A(n425), .ZN(n423) );
  INV_X1 U451 ( .A(KEYINPUT85), .ZN(n527) );
  AND2_X1 U452 ( .A1(n743), .A2(KEYINPUT85), .ZN(n530) );
  AND2_X1 U453 ( .A1(n526), .A2(n742), .ZN(n525) );
  NAND2_X1 U454 ( .A1(n528), .A2(n527), .ZN(n526) );
  INV_X1 U455 ( .A(n743), .ZN(n528) );
  XNOR2_X1 U456 ( .A(n632), .B(n631), .ZN(n754) );
  XOR2_X1 U457 ( .A(G104), .B(G110), .Z(n555) );
  NOR2_X1 U458 ( .A1(n366), .A2(n539), .ZN(n537) );
  NAND2_X1 U459 ( .A1(n404), .A2(n398), .ZN(n397) );
  AND2_X1 U460 ( .A1(n653), .A2(n642), .ZN(n404) );
  NAND2_X1 U461 ( .A1(n401), .A2(n400), .ZN(n399) );
  NAND2_X1 U462 ( .A1(n402), .A2(n420), .ZN(n400) );
  NAND2_X1 U463 ( .A1(n395), .A2(n402), .ZN(n401) );
  INV_X1 U464 ( .A(KEYINPUT66), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n406), .B(KEYINPUT72), .ZN(n405) );
  NAND2_X1 U466 ( .A1(n370), .A2(n425), .ZN(n416) );
  INV_X1 U467 ( .A(KEYINPUT30), .ZN(n498) );
  OR2_X1 U468 ( .A1(n574), .A2(G902), .ZN(n575) );
  XNOR2_X1 U469 ( .A(n675), .B(KEYINPUT1), .ZN(n756) );
  XNOR2_X1 U470 ( .A(n577), .B(n384), .ZN(n714) );
  XNOR2_X1 U471 ( .A(n579), .B(n385), .ZN(n384) );
  XNOR2_X1 U472 ( .A(n446), .B(n442), .ZN(n579) );
  XNOR2_X1 U473 ( .A(n565), .B(n566), .ZN(n512) );
  XNOR2_X1 U474 ( .A(n567), .B(n511), .ZN(n510) );
  XNOR2_X1 U475 ( .A(KEYINPUT81), .B(KEYINPUT23), .ZN(n511) );
  XNOR2_X1 U476 ( .A(G134), .B(G122), .ZN(n621) );
  AND2_X1 U477 ( .A1(n459), .A2(n546), .ZN(n458) );
  NOR2_X1 U478 ( .A1(n710), .A2(n712), .ZN(n473) );
  AND2_X1 U479 ( .A1(n479), .A2(n712), .ZN(n475) );
  NAND2_X1 U480 ( .A1(n480), .A2(n484), .ZN(n472) );
  NOR2_X1 U481 ( .A1(n363), .A2(KEYINPUT44), .ZN(n414) );
  AND2_X1 U482 ( .A1(n694), .A2(n693), .ZN(n390) );
  XNOR2_X1 U483 ( .A(n740), .B(KEYINPUT88), .ZN(n389) );
  INV_X1 U484 ( .A(KEYINPUT67), .ZN(n543) );
  AND2_X1 U485 ( .A1(n420), .A2(KEYINPUT68), .ZN(n417) );
  XOR2_X1 U486 ( .A(KEYINPUT18), .B(KEYINPUT78), .Z(n593) );
  XNOR2_X1 U487 ( .A(n590), .B(n589), .ZN(n591) );
  NAND2_X1 U488 ( .A1(n358), .A2(n457), .ZN(n448) );
  XOR2_X1 U489 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n610) );
  XNOR2_X1 U490 ( .A(G113), .B(n355), .ZN(n612) );
  XOR2_X1 U491 ( .A(G140), .B(G131), .Z(n613) );
  XNOR2_X1 U492 ( .A(n578), .B(n447), .ZN(n446) );
  XNOR2_X1 U493 ( .A(G137), .B(KEYINPUT76), .ZN(n578) );
  NAND2_X1 U494 ( .A1(n608), .A2(G210), .ZN(n447) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n442) );
  XNOR2_X1 U496 ( .A(G116), .B(KEYINPUT97), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n445), .B(KEYINPUT5), .ZN(n444) );
  INV_X1 U498 ( .A(KEYINPUT98), .ZN(n445) );
  INV_X1 U499 ( .A(G104), .ZN(n502) );
  AND2_X1 U500 ( .A1(n710), .A2(G210), .ZN(n483) );
  NAND2_X1 U501 ( .A1(n523), .A2(n527), .ZN(n522) );
  NAND2_X1 U502 ( .A1(G234), .A2(G237), .ZN(n582) );
  XOR2_X1 U503 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n583) );
  INV_X1 U504 ( .A(KEYINPUT109), .ZN(n681) );
  NAND2_X1 U505 ( .A1(n680), .A2(n769), .ZN(n682) );
  OR2_X1 U506 ( .A1(G237), .A2(G902), .ZN(n601) );
  XOR2_X1 U507 ( .A(G902), .B(KEYINPUT15), .Z(n703) );
  INV_X1 U508 ( .A(n754), .ZN(n439) );
  INV_X1 U509 ( .A(KEYINPUT3), .ZN(n549) );
  XNOR2_X1 U510 ( .A(G110), .B(KEYINPUT16), .ZN(n596) );
  XNOR2_X1 U511 ( .A(n607), .B(n503), .ZN(n597) );
  XNOR2_X1 U512 ( .A(n557), .B(n556), .ZN(n561) );
  NOR2_X1 U513 ( .A1(n399), .A2(n397), .ZN(n403) );
  XNOR2_X1 U514 ( .A(n499), .B(KEYINPUT41), .ZN(n768) );
  NAND2_X1 U515 ( .A1(n520), .A2(n521), .ZN(n434) );
  XNOR2_X1 U516 ( .A(n678), .B(KEYINPUT28), .ZN(n489) );
  BUF_X1 U517 ( .A(n818), .Z(n492) );
  XNOR2_X1 U518 ( .A(n514), .B(n509), .ZN(n569) );
  XNOR2_X1 U519 ( .A(n512), .B(n510), .ZN(n509) );
  XOR2_X1 U520 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n624) );
  INV_X1 U521 ( .A(KEYINPUT105), .ZN(n495) );
  XNOR2_X1 U522 ( .A(n508), .B(n507), .ZN(n828) );
  INV_X1 U523 ( .A(KEYINPUT103), .ZN(n507) );
  NOR2_X1 U524 ( .A1(n501), .A2(n364), .ZN(n408) );
  XNOR2_X1 U525 ( .A(n491), .B(n490), .ZN(n720) );
  INV_X1 U526 ( .A(KEYINPUT99), .ZN(n490) );
  AND2_X1 U527 ( .A1(n648), .A2(n521), .ZN(n491) );
  NOR2_X1 U528 ( .A1(n501), .A2(n409), .ZN(n407) );
  INV_X1 U529 ( .A(n441), .ZN(n409) );
  AND2_X1 U530 ( .A1(n465), .A2(n464), .ZN(n463) );
  AND2_X1 U531 ( .A1(n472), .A2(n478), .ZN(n477) );
  NAND2_X1 U532 ( .A1(n476), .A2(n475), .ZN(n474) );
  AND2_X1 U533 ( .A1(n452), .A2(n450), .ZN(n363) );
  NAND2_X1 U534 ( .A1(n677), .A2(n550), .ZN(n364) );
  AND2_X1 U535 ( .A1(n481), .A2(n547), .ZN(n365) );
  AND2_X1 U536 ( .A1(KEYINPUT2), .A2(n703), .ZN(n366) );
  AND2_X1 U537 ( .A1(n466), .A2(KEYINPUT60), .ZN(n367) );
  INV_X1 U538 ( .A(G953), .ZN(n746) );
  OR2_X1 U539 ( .A1(n452), .A2(n450), .ZN(n368) );
  XOR2_X1 U540 ( .A(G131), .B(G134), .Z(n369) );
  XNOR2_X1 U541 ( .A(n602), .B(KEYINPUT93), .ZN(n603) );
  AND2_X1 U542 ( .A1(n424), .A2(n417), .ZN(n370) );
  AND2_X1 U543 ( .A1(n747), .A2(n469), .ZN(n371) );
  AND2_X1 U544 ( .A1(n747), .A2(n483), .ZN(n372) );
  AND2_X1 U545 ( .A1(n747), .A2(G469), .ZN(n373) );
  AND2_X1 U546 ( .A1(n468), .A2(n367), .ZN(n374) );
  NOR2_X1 U547 ( .A1(n668), .A2(KEYINPUT77), .ZN(n375) );
  BUF_X1 U548 ( .A(n753), .Z(n500) );
  INV_X1 U549 ( .A(KEYINPUT34), .ZN(n457) );
  INV_X1 U550 ( .A(n710), .ZN(n711) );
  XNOR2_X1 U551 ( .A(KEYINPUT87), .B(KEYINPUT46), .ZN(n376) );
  XOR2_X1 U552 ( .A(n563), .B(n562), .Z(n377) );
  INV_X1 U553 ( .A(KEYINPUT68), .ZN(n422) );
  INV_X1 U554 ( .A(KEYINPUT44), .ZN(n420) );
  OR2_X1 U555 ( .A1(n539), .A2(n540), .ZN(n378) );
  INV_X1 U556 ( .A(KEYINPUT82), .ZN(n540) );
  INV_X1 U557 ( .A(n470), .ZN(n469) );
  AND2_X1 U558 ( .A1(n790), .A2(n546), .ZN(n379) );
  AND2_X1 U559 ( .A1(KEYINPUT66), .A2(KEYINPUT44), .ZN(n380) );
  XOR2_X1 U560 ( .A(KEYINPUT89), .B(KEYINPUT63), .Z(n381) );
  NOR2_X1 U561 ( .A1(n492), .A2(G952), .ZN(n798) );
  INV_X1 U562 ( .A(n798), .ZN(n547) );
  INV_X1 U563 ( .A(n712), .ZN(n484) );
  INV_X1 U564 ( .A(KEYINPUT60), .ZN(n546) );
  INV_X1 U565 ( .A(n412), .ZN(n382) );
  INV_X1 U566 ( .A(n412), .ZN(n436) );
  NAND2_X1 U567 ( .A1(n636), .A2(n407), .ZN(n644) );
  NAND2_X1 U568 ( .A1(n636), .A2(n408), .ZN(n508) );
  BUF_X1 U569 ( .A(n731), .Z(n383) );
  BUF_X1 U570 ( .A(n763), .Z(n497) );
  NAND2_X1 U571 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U572 ( .A1(n391), .A2(n392), .ZN(n388) );
  OR2_X2 U573 ( .A1(n714), .A2(G902), .ZN(n542) );
  INV_X1 U574 ( .A(n598), .ZN(n385) );
  NAND2_X1 U575 ( .A1(n429), .A2(n428), .ZN(n392) );
  AND2_X2 U576 ( .A1(n516), .A2(n519), .ZN(n393) );
  NAND2_X1 U577 ( .A1(n647), .A2(n646), .ZN(n645) );
  XNOR2_X2 U578 ( .A(n629), .B(G478), .ZN(n647) );
  XNOR2_X1 U579 ( .A(n628), .B(n627), .ZN(n792) );
  XNOR2_X1 U580 ( .A(n394), .B(n671), .ZN(n700) );
  NAND2_X1 U581 ( .A1(n691), .A2(n770), .ZN(n394) );
  NAND2_X1 U582 ( .A1(n396), .A2(n395), .ZN(n406) );
  INV_X1 U583 ( .A(n643), .ZN(n395) );
  NAND2_X1 U584 ( .A1(n418), .A2(n416), .ZN(n396) );
  NAND2_X1 U585 ( .A1(n643), .A2(n380), .ZN(n398) );
  AND2_X2 U586 ( .A1(n533), .A2(n532), .ZN(n411) );
  NAND2_X1 U587 ( .A1(n412), .A2(n711), .ZN(n479) );
  NAND2_X1 U588 ( .A1(n412), .A2(n466), .ZN(n460) );
  NAND2_X1 U589 ( .A1(n412), .A2(n473), .ZN(n478) );
  NAND2_X1 U590 ( .A1(n412), .A2(n379), .ZN(n464) );
  NAND2_X1 U591 ( .A1(n412), .A2(n790), .ZN(n461) );
  NAND2_X1 U592 ( .A1(n449), .A2(n363), .ZN(n424) );
  NOR2_X1 U593 ( .A1(n414), .A2(KEYINPUT68), .ZN(n413) );
  NAND2_X1 U594 ( .A1(n453), .A2(n420), .ZN(n415) );
  NAND2_X1 U595 ( .A1(n425), .A2(n424), .ZN(n829) );
  XNOR2_X2 U596 ( .A(n427), .B(n549), .ZN(n802) );
  XNOR2_X2 U597 ( .A(G119), .B(G113), .ZN(n427) );
  INV_X1 U598 ( .A(n825), .ZN(n428) );
  NOR2_X1 U599 ( .A1(n831), .A2(n376), .ZN(n429) );
  NAND2_X1 U600 ( .A1(n831), .A2(n376), .ZN(n430) );
  NAND2_X1 U601 ( .A1(n825), .A2(n376), .ZN(n431) );
  NOR2_X1 U602 ( .A1(n362), .A2(n433), .ZN(n432) );
  NAND2_X1 U603 ( .A1(n705), .A2(n371), .ZN(n468) );
  NAND2_X1 U604 ( .A1(n705), .A2(n372), .ZN(n482) );
  NAND2_X1 U605 ( .A1(n705), .A2(n373), .ZN(n706) );
  NAND2_X1 U606 ( .A1(n705), .A2(n435), .ZN(n716) );
  AND2_X1 U607 ( .A1(n747), .A2(G472), .ZN(n435) );
  NAND2_X1 U608 ( .A1(n382), .A2(G478), .ZN(n791) );
  NAND2_X1 U609 ( .A1(n436), .A2(G217), .ZN(n795) );
  XNOR2_X2 U610 ( .A(n437), .B(KEYINPUT42), .ZN(n831) );
  NOR2_X2 U611 ( .A1(n768), .A2(n684), .ZN(n437) );
  NAND2_X1 U612 ( .A1(n828), .A2(n830), .ZN(n643) );
  NAND2_X1 U613 ( .A1(n757), .A2(n675), .ZN(n669) );
  XNOR2_X1 U614 ( .A(n611), .B(n440), .ZN(n615) );
  XNOR2_X1 U615 ( .A(n609), .B(n610), .ZN(n440) );
  XNOR2_X2 U616 ( .A(n617), .B(n618), .ZN(n646) );
  OR2_X1 U617 ( .A1(n441), .A2(n676), .ZN(n663) );
  NAND2_X1 U618 ( .A1(n501), .A2(n441), .ZN(n580) );
  INV_X1 U619 ( .A(n453), .ZN(n449) );
  INV_X1 U620 ( .A(n641), .ZN(n450) );
  NAND2_X1 U621 ( .A1(n453), .A2(n641), .ZN(n451) );
  NAND2_X1 U622 ( .A1(n778), .A2(KEYINPUT34), .ZN(n452) );
  NAND2_X1 U623 ( .A1(n505), .A2(KEYINPUT34), .ZN(n455) );
  NAND2_X1 U624 ( .A1(n460), .A2(n458), .ZN(n465) );
  NAND2_X1 U625 ( .A1(n470), .A2(n466), .ZN(n459) );
  NAND2_X1 U626 ( .A1(n374), .A2(n461), .ZN(n462) );
  NAND2_X1 U627 ( .A1(n463), .A2(n462), .ZN(G60) );
  NAND2_X1 U628 ( .A1(n548), .A2(G475), .ZN(n470) );
  NAND2_X1 U629 ( .A1(n471), .A2(n518), .ZN(n517) );
  AND2_X1 U630 ( .A1(n471), .A2(n375), .ZN(n520) );
  NAND2_X1 U631 ( .A1(n477), .A2(n474), .ZN(G51) );
  INV_X1 U632 ( .A(n480), .ZN(n476) );
  BUF_X1 U633 ( .A(n768), .Z(n485) );
  XNOR2_X1 U634 ( .A(n486), .B(KEYINPUT123), .ZN(G54) );
  NAND2_X1 U635 ( .A1(n488), .A2(n547), .ZN(n486) );
  NOR2_X2 U636 ( .A1(n794), .A2(G902), .ZN(n573) );
  NOR2_X2 U637 ( .A1(G902), .A2(n789), .ZN(n617) );
  XNOR2_X1 U638 ( .A(n625), .B(n624), .ZN(n628) );
  NAND2_X1 U639 ( .A1(n753), .A2(n754), .ZN(n637) );
  XNOR2_X2 U640 ( .A(n573), .B(n572), .ZN(n753) );
  NAND2_X1 U641 ( .A1(n662), .A2(n754), .ZN(n676) );
  XNOR2_X1 U642 ( .A(n706), .B(n377), .ZN(n488) );
  XNOR2_X1 U643 ( .A(n814), .B(n553), .ZN(n557) );
  NAND2_X1 U644 ( .A1(n665), .A2(n769), .ZN(n545) );
  XNOR2_X2 U645 ( .A(n506), .B(n603), .ZN(n665) );
  NAND2_X1 U646 ( .A1(n517), .A2(KEYINPUT77), .ZN(n516) );
  NAND2_X1 U647 ( .A1(n818), .A2(G234), .ZN(n515) );
  XNOR2_X2 U648 ( .A(n493), .B(G953), .ZN(n818) );
  XNOR2_X2 U649 ( .A(n637), .B(KEYINPUT69), .ZN(n757) );
  NAND2_X1 U650 ( .A1(n695), .A2(n665), .ZN(n494) );
  XNOR2_X2 U651 ( .A(n645), .B(n496), .ZN(n672) );
  XNOR2_X2 U652 ( .A(n619), .B(n559), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(n591), .ZN(n595) );
  INV_X1 U654 ( .A(n503), .ZN(n620) );
  INV_X1 U655 ( .A(n703), .ZN(n539) );
  NAND2_X1 U656 ( .A1(n538), .A2(n537), .ZN(n536) );
  XNOR2_X1 U657 ( .A(n504), .B(n381), .ZN(G57) );
  NAND2_X1 U658 ( .A1(n717), .A2(n547), .ZN(n504) );
  OR2_X2 U659 ( .A1(n707), .A2(n703), .ZN(n506) );
  INV_X1 U660 ( .A(n808), .ZN(n538) );
  XNOR2_X2 U661 ( .A(n513), .B(G140), .ZN(n565) );
  NAND2_X1 U662 ( .A1(n626), .A2(G221), .ZN(n514) );
  INV_X1 U663 ( .A(n668), .ZN(n518) );
  NAND2_X1 U664 ( .A1(n669), .A2(KEYINPUT77), .ZN(n519) );
  INV_X1 U665 ( .A(n669), .ZN(n521) );
  NAND2_X2 U666 ( .A1(n524), .A2(n522), .ZN(n704) );
  INV_X1 U667 ( .A(n531), .ZN(n523) );
  AND2_X2 U668 ( .A1(n529), .A2(n525), .ZN(n524) );
  NAND2_X1 U669 ( .A1(n531), .A2(n530), .ZN(n529) );
  NAND2_X1 U670 ( .A1(n817), .A2(n540), .ZN(n532) );
  NAND2_X1 U671 ( .A1(n534), .A2(n538), .ZN(n533) );
  NOR2_X2 U672 ( .A1(n817), .A2(n378), .ZN(n534) );
  NOR2_X1 U673 ( .A1(n817), .A2(n808), .ZN(n748) );
  XNOR2_X2 U674 ( .A(n674), .B(n673), .ZN(n825) );
  XNOR2_X1 U675 ( .A(n616), .B(n813), .ZN(n789) );
  INV_X1 U676 ( .A(KEYINPUT48), .ZN(n541) );
  XNOR2_X2 U677 ( .A(n542), .B(G472), .ZN(n763) );
  INV_X1 U678 ( .A(n501), .ZN(n696) );
  NAND2_X1 U679 ( .A1(n757), .A2(n756), .ZN(n649) );
  INV_X1 U680 ( .A(n790), .ZN(n548) );
  INV_X1 U681 ( .A(n500), .ZN(n550) );
  INV_X2 U682 ( .A(G143), .ZN(n558) );
  XNOR2_X1 U683 ( .A(KEYINPUT59), .B(KEYINPUT91), .ZN(n552) );
  XOR2_X1 U684 ( .A(n576), .B(G107), .Z(n553) );
  XNOR2_X1 U685 ( .A(n615), .B(n614), .ZN(n616) );
  INV_X1 U686 ( .A(n647), .ZN(n639) );
  XNOR2_X1 U687 ( .A(n714), .B(n713), .ZN(n715) );
  XOR2_X1 U688 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n563) );
  XOR2_X1 U689 ( .A(KEYINPUT95), .B(n565), .Z(n814) );
  NAND2_X1 U690 ( .A1(G227), .A2(n818), .ZN(n554) );
  XNOR2_X1 U691 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X2 U692 ( .A(n558), .B(G128), .ZN(n619) );
  XNOR2_X1 U693 ( .A(KEYINPUT4), .B(KEYINPUT65), .ZN(n559) );
  INV_X1 U694 ( .A(n577), .ZN(n560) );
  XNOR2_X1 U695 ( .A(n560), .B(n561), .ZN(n574) );
  XNOR2_X1 U696 ( .A(n574), .B(KEYINPUT122), .ZN(n562) );
  INV_X1 U697 ( .A(KEYINPUT45), .ZN(n655) );
  XOR2_X1 U698 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n564) );
  XNOR2_X1 U699 ( .A(G119), .B(G128), .ZN(n566) );
  XNOR2_X1 U700 ( .A(G110), .B(KEYINPUT24), .ZN(n567) );
  XNOR2_X1 U701 ( .A(n590), .B(KEYINPUT10), .ZN(n568) );
  XNOR2_X1 U702 ( .A(n568), .B(KEYINPUT71), .ZN(n813) );
  NAND2_X1 U703 ( .A1(n539), .A2(G234), .ZN(n570) );
  XNOR2_X1 U704 ( .A(n570), .B(KEYINPUT20), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G217), .A2(n630), .ZN(n571) );
  XNOR2_X2 U706 ( .A(n575), .B(G469), .ZN(n675) );
  NOR2_X1 U707 ( .A1(n500), .A2(n580), .ZN(n581) );
  XNOR2_X1 U708 ( .A(KEYINPUT80), .B(n581), .ZN(n634) );
  INV_X1 U709 ( .A(KEYINPUT0), .ZN(n606) );
  XNOR2_X1 U710 ( .A(n583), .B(n582), .ZN(n584) );
  NAND2_X1 U711 ( .A1(G952), .A2(n584), .ZN(n784) );
  NOR2_X1 U712 ( .A1(G953), .A2(n784), .ZN(n661) );
  NAND2_X1 U713 ( .A1(G902), .A2(n584), .ZN(n656) );
  INV_X1 U714 ( .A(n656), .ZN(n585) );
  NOR2_X1 U715 ( .A1(G898), .A2(n746), .ZN(n804) );
  NAND2_X1 U716 ( .A1(n585), .A2(n804), .ZN(n586) );
  XOR2_X1 U717 ( .A(KEYINPUT94), .B(n586), .Z(n587) );
  NOR2_X1 U718 ( .A1(n661), .A2(n587), .ZN(n605) );
  INV_X1 U719 ( .A(KEYINPUT19), .ZN(n604) );
  NAND2_X1 U720 ( .A1(G214), .A2(n601), .ZN(n769) );
  XOR2_X1 U721 ( .A(KEYINPUT17), .B(KEYINPUT92), .Z(n589) );
  NAND2_X1 U722 ( .A1(G224), .A2(n818), .ZN(n592) );
  XNOR2_X1 U723 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U724 ( .A(n595), .B(n594), .ZN(n600) );
  XNOR2_X1 U725 ( .A(n799), .B(n598), .ZN(n599) );
  XNOR2_X1 U726 ( .A(n599), .B(n600), .ZN(n707) );
  NAND2_X1 U727 ( .A1(n601), .A2(G210), .ZN(n602) );
  XNOR2_X1 U728 ( .A(KEYINPUT13), .B(G475), .ZN(n618) );
  XNOR2_X1 U729 ( .A(n607), .B(KEYINPUT100), .ZN(n611) );
  NAND2_X1 U730 ( .A1(G214), .A2(n608), .ZN(n609) );
  XNOR2_X1 U731 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U732 ( .A(n619), .B(KEYINPUT9), .ZN(n623) );
  XNOR2_X1 U733 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U734 ( .A(n622), .B(n623), .ZN(n625) );
  NAND2_X1 U735 ( .A1(G217), .A2(n626), .ZN(n627) );
  OR2_X1 U736 ( .A1(n646), .A2(n639), .ZN(n772) );
  XOR2_X1 U737 ( .A(KEYINPUT21), .B(KEYINPUT96), .Z(n632) );
  NAND2_X1 U738 ( .A1(n630), .A2(G221), .ZN(n631) );
  NAND2_X1 U739 ( .A1(n634), .A2(n636), .ZN(n635) );
  XNOR2_X1 U740 ( .A(n635), .B(KEYINPUT32), .ZN(n830) );
  INV_X1 U741 ( .A(n763), .ZN(n677) );
  XNOR2_X1 U742 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n641) );
  XNOR2_X1 U743 ( .A(KEYINPUT104), .B(KEYINPUT33), .ZN(n638) );
  NAND2_X1 U744 ( .A1(n646), .A2(n639), .ZN(n689) );
  XNOR2_X1 U745 ( .A(n689), .B(KEYINPUT79), .ZN(n640) );
  NAND2_X1 U746 ( .A1(n829), .A2(KEYINPUT44), .ZN(n642) );
  NOR2_X1 U747 ( .A1(n550), .A2(n644), .ZN(n718) );
  NOR2_X1 U748 ( .A1(n647), .A2(n646), .ZN(n735) );
  NOR2_X1 U749 ( .A1(n672), .A2(n735), .ZN(n773) );
  NOR2_X1 U750 ( .A1(n497), .A2(n505), .ZN(n648) );
  NOR2_X1 U751 ( .A1(n677), .A2(n649), .ZN(n765) );
  NAND2_X1 U752 ( .A1(n358), .A2(n765), .ZN(n650) );
  XNOR2_X1 U753 ( .A(n650), .B(KEYINPUT31), .ZN(n736) );
  NOR2_X1 U754 ( .A1(n720), .A2(n736), .ZN(n651) );
  NOR2_X1 U755 ( .A1(n773), .A2(n651), .ZN(n652) );
  NOR2_X1 U756 ( .A1(n718), .A2(n652), .ZN(n653) );
  NAND2_X1 U757 ( .A1(n769), .A2(n731), .ZN(n664) );
  NOR2_X1 U758 ( .A1(G900), .A2(n656), .ZN(n658) );
  INV_X1 U759 ( .A(n492), .ZN(n657) );
  NAND2_X1 U760 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U761 ( .A(KEYINPUT106), .B(n659), .Z(n660) );
  NOR2_X1 U762 ( .A1(n661), .A2(n660), .ZN(n668) );
  NOR2_X2 U763 ( .A1(n664), .A2(n663), .ZN(n695) );
  NAND2_X1 U764 ( .A1(n763), .A2(n769), .ZN(n670) );
  BUF_X1 U765 ( .A(n680), .Z(n770) );
  XOR2_X1 U766 ( .A(KEYINPUT39), .B(KEYINPUT73), .Z(n671) );
  NAND2_X1 U767 ( .A1(n700), .A2(n672), .ZN(n674) );
  XOR2_X1 U768 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n673) );
  INV_X1 U769 ( .A(KEYINPUT74), .ZN(n688) );
  NOR2_X1 U770 ( .A1(n688), .A2(KEYINPUT47), .ZN(n687) );
  INV_X1 U771 ( .A(n773), .ZN(n685) );
  NAND2_X1 U772 ( .A1(n688), .A2(KEYINPUT47), .ZN(n692) );
  NOR2_X1 U773 ( .A1(n698), .A2(n689), .ZN(n690) );
  NAND2_X1 U774 ( .A1(n361), .A2(n690), .ZN(n728) );
  AND2_X1 U775 ( .A1(n692), .A2(n728), .ZN(n693) );
  NAND2_X1 U776 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U777 ( .A(KEYINPUT43), .B(n697), .ZN(n699) );
  NAND2_X1 U778 ( .A1(n699), .A2(n698), .ZN(n743) );
  BUF_X1 U779 ( .A(n700), .Z(n701) );
  NAND2_X1 U780 ( .A1(n701), .A2(n735), .ZN(n742) );
  INV_X1 U781 ( .A(KEYINPUT83), .ZN(n702) );
  XNOR2_X2 U782 ( .A(n704), .B(n702), .ZN(n817) );
  XOR2_X1 U783 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n709) );
  XNOR2_X1 U784 ( .A(n707), .B(KEYINPUT55), .ZN(n708) );
  XNOR2_X1 U785 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U786 ( .A(KEYINPUT86), .B(KEYINPUT56), .ZN(n712) );
  XOR2_X1 U787 ( .A(KEYINPUT62), .B(KEYINPUT90), .Z(n713) );
  XNOR2_X1 U788 ( .A(n716), .B(n715), .ZN(n717) );
  XOR2_X1 U789 ( .A(G101), .B(n718), .Z(G3) );
  NAND2_X1 U790 ( .A1(n383), .A2(n720), .ZN(n719) );
  XNOR2_X1 U791 ( .A(n719), .B(G104), .ZN(G6) );
  XNOR2_X1 U792 ( .A(G107), .B(KEYINPUT27), .ZN(n724) );
  XOR2_X1 U793 ( .A(KEYINPUT110), .B(KEYINPUT26), .Z(n722) );
  NAND2_X1 U794 ( .A1(n720), .A2(n735), .ZN(n721) );
  XNOR2_X1 U795 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U796 ( .A(n724), .B(n723), .ZN(G9) );
  XOR2_X1 U797 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n726) );
  NAND2_X1 U798 ( .A1(n729), .A2(n735), .ZN(n725) );
  XNOR2_X1 U799 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U800 ( .A(G128), .B(n727), .ZN(G30) );
  XNOR2_X1 U801 ( .A(n355), .B(n728), .ZN(G45) );
  NAND2_X1 U802 ( .A1(n383), .A2(n729), .ZN(n730) );
  XNOR2_X1 U803 ( .A(n730), .B(G146), .ZN(G48) );
  XOR2_X1 U804 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n733) );
  NAND2_X1 U805 ( .A1(n736), .A2(n731), .ZN(n732) );
  XNOR2_X1 U806 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U807 ( .A(G113), .B(n734), .ZN(G15) );
  XOR2_X1 U808 ( .A(G116), .B(KEYINPUT115), .Z(n738) );
  NAND2_X1 U809 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U810 ( .A(n738), .B(n737), .ZN(G18) );
  XOR2_X1 U811 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n739) );
  XNOR2_X1 U812 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U813 ( .A(G125), .B(n741), .ZN(G27) );
  XNOR2_X1 U814 ( .A(G134), .B(n742), .ZN(G36) );
  XNOR2_X1 U815 ( .A(G140), .B(n743), .ZN(G42) );
  NOR2_X1 U816 ( .A1(n485), .A2(n778), .ZN(n744) );
  XOR2_X1 U817 ( .A(KEYINPUT120), .B(n744), .Z(n745) );
  NAND2_X1 U818 ( .A1(n746), .A2(n745), .ZN(n752) );
  INV_X1 U819 ( .A(n747), .ZN(n750) );
  NOR2_X1 U820 ( .A1(n748), .A2(KEYINPUT2), .ZN(n749) );
  NOR2_X1 U821 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U822 ( .A1(n752), .A2(n751), .ZN(n787) );
  NOR2_X1 U823 ( .A1(n754), .A2(n500), .ZN(n755) );
  XNOR2_X1 U824 ( .A(KEYINPUT49), .B(n755), .ZN(n761) );
  NOR2_X1 U825 ( .A1(n757), .A2(n501), .ZN(n759) );
  XNOR2_X1 U826 ( .A(KEYINPUT117), .B(KEYINPUT50), .ZN(n758) );
  XNOR2_X1 U827 ( .A(n759), .B(n758), .ZN(n760) );
  NAND2_X1 U828 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U829 ( .A1(n497), .A2(n762), .ZN(n764) );
  NOR2_X1 U830 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U831 ( .A(KEYINPUT51), .B(n766), .Z(n767) );
  NOR2_X1 U832 ( .A1(n485), .A2(n767), .ZN(n781) );
  NOR2_X1 U833 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U834 ( .A1(n772), .A2(n771), .ZN(n776) );
  NOR2_X1 U835 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U836 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U837 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U838 ( .A(n779), .B(KEYINPUT118), .ZN(n780) );
  NOR2_X1 U839 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U840 ( .A(KEYINPUT52), .B(n782), .ZN(n783) );
  NOR2_X1 U841 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U842 ( .A(n785), .B(KEYINPUT119), .ZN(n786) );
  NAND2_X1 U843 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U844 ( .A(KEYINPUT53), .B(n788), .Z(G75) );
  XNOR2_X1 U845 ( .A(n789), .B(n552), .ZN(n790) );
  XNOR2_X1 U846 ( .A(n791), .B(n792), .ZN(n793) );
  NOR2_X1 U847 ( .A1(n798), .A2(n793), .ZN(G63) );
  XNOR2_X1 U848 ( .A(n794), .B(KEYINPUT124), .ZN(n796) );
  XNOR2_X1 U849 ( .A(n795), .B(n796), .ZN(n797) );
  NOR2_X1 U850 ( .A1(n798), .A2(n797), .ZN(G66) );
  XNOR2_X1 U851 ( .A(G101), .B(n799), .ZN(n800) );
  XNOR2_X1 U852 ( .A(n800), .B(KEYINPUT125), .ZN(n801) );
  XOR2_X1 U853 ( .A(n802), .B(n801), .Z(n803) );
  NOR2_X1 U854 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U855 ( .A(KEYINPUT126), .B(n805), .Z(n812) );
  NAND2_X1 U856 ( .A1(G953), .A2(G224), .ZN(n806) );
  XNOR2_X1 U857 ( .A(KEYINPUT61), .B(n806), .ZN(n807) );
  NAND2_X1 U858 ( .A1(n807), .A2(G898), .ZN(n810) );
  OR2_X1 U859 ( .A1(n808), .A2(G953), .ZN(n809) );
  NAND2_X1 U860 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U861 ( .A(n812), .B(n811), .Z(G69) );
  XOR2_X1 U862 ( .A(n814), .B(n813), .Z(n815) );
  XNOR2_X1 U863 ( .A(n816), .B(n815), .ZN(n820) );
  XNOR2_X1 U864 ( .A(n817), .B(n820), .ZN(n819) );
  NAND2_X1 U865 ( .A1(n819), .A2(n492), .ZN(n824) );
  XNOR2_X1 U866 ( .A(G227), .B(n820), .ZN(n821) );
  NAND2_X1 U867 ( .A1(n821), .A2(G900), .ZN(n822) );
  NAND2_X1 U868 ( .A1(n822), .A2(G953), .ZN(n823) );
  NAND2_X1 U869 ( .A1(n824), .A2(n823), .ZN(G72) );
  XNOR2_X1 U870 ( .A(n825), .B(G131), .ZN(n826) );
  XNOR2_X1 U871 ( .A(n826), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U872 ( .A(G110), .B(KEYINPUT111), .Z(n827) );
  XNOR2_X1 U873 ( .A(n828), .B(n827), .ZN(G12) );
  XOR2_X1 U874 ( .A(n829), .B(G122), .Z(G24) );
  XNOR2_X1 U875 ( .A(n830), .B(G119), .ZN(G21) );
  XOR2_X1 U876 ( .A(n831), .B(G137), .Z(G39) );
endmodule

