//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n445, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G259));
  XOR2_X1   g021(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n457), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n473), .A2(new_n475), .A3(G125), .ZN(new_n476));
  INV_X1    g051(.A(G113), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT69), .B1(new_n477), .B2(new_n465), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(G113), .A3(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(G2105), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT70), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n473), .A2(new_n475), .A3(G125), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(new_n478), .A3(new_n480), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n485), .A2(new_n486), .A3(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n472), .B1(new_n483), .B2(new_n487), .ZN(G160));
  INV_X1    g063(.A(new_n470), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n468), .A2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(G124), .B2(new_n494), .ZN(G162));
  NAND4_X1  g070(.A1(new_n473), .A2(new_n475), .A3(G138), .A4(new_n469), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n468), .A2(new_n498), .A3(G138), .A4(new_n469), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n473), .A2(new_n475), .A3(G126), .A4(G2105), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n500), .A2(KEYINPUT71), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT71), .B1(new_n500), .B2(new_n504), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT72), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(new_n521), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n520), .A2(new_n527), .ZN(G166));
  NAND4_X1  g103(.A1(new_n515), .A2(G63), .A3(G651), .A4(new_n516), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n530), .B2(new_n522), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT73), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n517), .A2(new_n521), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n532), .A2(new_n533), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n531), .A2(KEYINPUT73), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n523), .A2(G51), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n540), .B1(new_n541), .B2(new_n529), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n535), .B(new_n537), .C1(new_n539), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT74), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n538), .A2(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n519), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT75), .B(G52), .Z(new_n549));
  OAI22_X1  g124(.A1(new_n525), .A2(new_n548), .B1(new_n522), .B2(new_n549), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(G171));
  AOI22_X1  g128(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n519), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n523), .A2(G43), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n525), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(new_n523), .A2(G53), .ZN(new_n566));
  AND2_X1   g141(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n515), .A2(new_n516), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n534), .A2(G91), .B1(new_n572), .B2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n568), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  AND2_X1   g150(.A1(new_n538), .A2(new_n544), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  OAI21_X1  g152(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n517), .A2(G87), .A3(new_n521), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n523), .A2(G49), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND3_X1  g156(.A1(new_n515), .A2(G61), .A3(new_n516), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n515), .A2(G86), .A3(new_n516), .A4(new_n521), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n521), .A2(G48), .A3(G543), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n585), .A2(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n570), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT78), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  XNOR2_X1  g169(.A(KEYINPUT79), .B(G47), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n534), .A2(G85), .B1(new_n523), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n594), .A2(KEYINPUT80), .A3(new_n596), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G290));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n534), .A2(new_n602), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(KEYINPUT10), .B1(new_n525), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n523), .A2(G54), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n519), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G171), .B2(new_n612), .ZN(G284));
  OAI21_X1  g189(.A(new_n613), .B1(G171), .B2(new_n612), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  XOR2_X1   g191(.A(G299), .B(KEYINPUT81), .Z(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(G868), .B2(new_n617), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(G868), .B2(new_n617), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n610), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n610), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g199(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n625));
  XNOR2_X1  g200(.A(G323), .B(new_n625), .ZN(G282));
  NAND2_X1  g201(.A1(new_n468), .A2(new_n466), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n489), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n494), .A2(G123), .ZN(new_n632));
  OR2_X1    g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n633), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n630), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT15), .ZN(new_n642));
  INV_X1    g217(.A(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT14), .ZN(new_n645));
  XOR2_X1   g220(.A(G2443), .B(G2446), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n646), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n647), .B2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n639), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n657), .A2(new_n638), .A3(new_n653), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n658), .A3(G14), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT83), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n661));
  NAND4_X1  g236(.A1(new_n656), .A2(new_n658), .A3(new_n661), .A4(G14), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n665), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n667), .A2(new_n668), .ZN(new_n674));
  AOI21_X1  g249(.A(KEYINPUT18), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n672), .B(new_n675), .Z(G227));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n687), .B(new_n688), .C1(new_n686), .C2(new_n685), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  INV_X1    g267(.A(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n691), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(KEYINPUT97), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n698), .A2(KEYINPUT23), .A3(G20), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT23), .ZN(new_n700));
  INV_X1    g275(.A(G20), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(G16), .ZN(new_n702));
  INV_X1    g277(.A(G299), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n699), .B(new_n702), .C1(new_n703), .C2(new_n698), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1956), .ZN(new_n705));
  NOR2_X1   g280(.A1(G29), .A2(G35), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G162), .B2(G29), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT29), .B(G2090), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(G29), .A2(G33), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n466), .A2(G103), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT25), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n489), .A2(G139), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n712), .B(new_n713), .C1(new_n469), .C2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n710), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G2072), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G11), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(KEYINPUT31), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(KEYINPUT31), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n709), .A2(new_n719), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n705), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n716), .A2(G27), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G164), .B2(new_n716), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(G2078), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT30), .B(G28), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n717), .A2(new_n718), .B1(new_n716), .B2(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n635), .A2(new_n716), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n724), .A2(new_n727), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n698), .A2(G5), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G171), .B2(new_n698), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT95), .B(G1961), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n726), .A2(G2078), .ZN(new_n736));
  AOI22_X1  g311(.A1(G141), .A2(new_n489), .B1(new_n494), .B2(G129), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n466), .A2(G105), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT26), .Z(new_n740));
  NAND3_X1  g315(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G32), .B(new_n741), .S(G29), .Z(new_n742));
  XOR2_X1   g317(.A(KEYINPUT27), .B(G1996), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n731), .A2(new_n735), .A3(new_n736), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(G166), .A2(G16), .ZN(new_n746));
  OR2_X1    g321(.A1(G16), .A2(G22), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT87), .B(G1971), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n746), .B2(new_n747), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n698), .A2(G23), .ZN(new_n751));
  INV_X1    g326(.A(G288), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n698), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT33), .B(G1976), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT86), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n753), .A2(new_n756), .ZN(new_n758));
  OAI22_X1  g333(.A1(new_n749), .A2(new_n750), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  MUX2_X1   g334(.A(G6), .B(G305), .S(G16), .Z(new_n760));
  XOR2_X1   g335(.A(KEYINPUT32), .B(G1981), .Z(new_n761));
  XOR2_X1   g336(.A(new_n760), .B(new_n761), .Z(new_n762));
  OR3_X1    g337(.A1(new_n759), .A2(new_n762), .A3(KEYINPUT34), .ZN(new_n763));
  OAI21_X1  g338(.A(KEYINPUT34), .B1(new_n759), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n716), .A2(G25), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n489), .A2(G131), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n494), .A2(G119), .ZN(new_n767));
  OR2_X1    g342(.A1(G95), .A2(G2105), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n768), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n765), .B1(new_n771), .B2(new_n716), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT35), .B(G1991), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n772), .B(new_n774), .ZN(new_n775));
  AND3_X1   g350(.A1(new_n763), .A2(new_n764), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT84), .ZN(new_n777));
  INV_X1    g352(.A(G24), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G16), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G290), .B2(G16), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n779), .B1(new_n781), .B2(new_n777), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT85), .B(G1986), .Z(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT88), .B(KEYINPUT36), .Z(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n782), .A2(new_n784), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n776), .A2(new_n785), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n698), .A2(G4), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n610), .B2(new_n698), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(KEYINPUT89), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(KEYINPUT89), .ZN(new_n793));
  INV_X1    g368(.A(G1348), .ZN(new_n794));
  OR3_X1    g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n716), .A2(G26), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n489), .A2(G140), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n494), .A2(G128), .ZN(new_n798));
  OAI21_X1  g373(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n469), .A2(G116), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n796), .B1(new_n801), .B2(G29), .ZN(new_n802));
  MUX2_X1   g377(.A(new_n796), .B(new_n802), .S(KEYINPUT28), .Z(new_n803));
  INV_X1    g378(.A(G2067), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(G19), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT90), .B1(new_n806), .B2(G16), .ZN(new_n807));
  OR3_X1    g382(.A1(new_n806), .A2(KEYINPUT90), .A3(G16), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n807), .B(new_n808), .C1(new_n559), .C2(new_n698), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1341), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n794), .B1(new_n792), .B2(new_n793), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n795), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT91), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n795), .A2(new_n811), .A3(KEYINPUT91), .A4(new_n812), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND3_X1   g392(.A1(new_n745), .A2(new_n789), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n698), .A2(G21), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G168), .B2(new_n698), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT94), .B(G1966), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(G160), .A2(G29), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT24), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n716), .B1(new_n825), .B2(G34), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT92), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(G34), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n827), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n824), .A2(G2084), .A3(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT93), .Z(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n782), .B(new_n783), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n787), .B1(new_n835), .B2(new_n776), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n818), .A2(new_n823), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n824), .A2(new_n831), .ZN(new_n839));
  INV_X1    g414(.A(G2084), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT96), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n697), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n745), .A2(new_n789), .A3(new_n817), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n844), .A2(new_n833), .A3(new_n836), .ZN(new_n845));
  INV_X1    g420(.A(new_n842), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n845), .A2(KEYINPUT97), .A3(new_n846), .A4(new_n823), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(G311));
  OAI21_X1  g423(.A(KEYINPUT98), .B1(new_n838), .B2(new_n842), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n845), .A2(new_n850), .A3(new_n846), .A4(new_n823), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G150));
  AOI22_X1  g427(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(new_n519), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n523), .A2(G55), .ZN(new_n855));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n525), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n858));
  OR3_X1    g433(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n854), .B2(new_n857), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n559), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n559), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n854), .A2(new_n857), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n610), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT39), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n867), .B(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(G860), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT101), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n863), .A2(G860), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(G145));
  XOR2_X1   g450(.A(new_n770), .B(new_n628), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n489), .A2(G142), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT103), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n494), .A2(G130), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n469), .A2(G118), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n878), .B(new_n879), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n876), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n715), .B(new_n741), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n502), .A2(new_n503), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(new_n497), .B2(new_n499), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n801), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n886), .B(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n885), .B(new_n890), .Z(new_n891));
  XNOR2_X1  g466(.A(G162), .B(KEYINPUT102), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n635), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(G160), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n890), .B(new_n883), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(KEYINPUT104), .B(G37), .Z(new_n898));
  AND3_X1   g473(.A1(new_n895), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(KEYINPUT40), .Z(G395));
  NOR2_X1   g475(.A1(new_n863), .A2(G868), .ZN(new_n901));
  XNOR2_X1  g476(.A(G166), .B(G288), .ZN(new_n902));
  INV_X1    g477(.A(new_n600), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT80), .B1(new_n594), .B2(new_n596), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(G166), .B(new_n752), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(new_n599), .A3(new_n600), .ZN(new_n907));
  XOR2_X1   g482(.A(G305), .B(KEYINPUT107), .Z(new_n908));
  AND3_X1   g483(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n908), .B1(new_n905), .B2(new_n907), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n911), .A2(KEYINPUT108), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n912), .A2(KEYINPUT42), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n865), .B(new_n622), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n703), .A2(new_n610), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  OAI21_X1  g491(.A(G299), .B1(new_n606), .B2(new_n609), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n914), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n915), .A2(new_n917), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT106), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n912), .A2(KEYINPUT42), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n913), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n925), .A2(new_n926), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n929), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n901), .B1(new_n931), .B2(G868), .ZN(G295));
  AOI21_X1  g507(.A(new_n901), .B1(new_n931), .B2(G868), .ZN(G331));
  NOR2_X1   g508(.A1(G286), .A2(G171), .ZN(new_n934));
  NOR2_X1   g509(.A1(G301), .A2(G168), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n865), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n865), .ZN(new_n937));
  NAND2_X1  g512(.A1(G286), .A2(G171), .ZN(new_n938));
  NAND2_X1  g513(.A1(G301), .A2(G168), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n936), .A2(new_n920), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n923), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n936), .B2(new_n940), .ZN(new_n943));
  OAI22_X1  g518(.A1(new_n941), .A2(new_n943), .B1(new_n909), .B2(new_n910), .ZN(new_n944));
  INV_X1    g519(.A(new_n940), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n937), .B1(new_n939), .B2(new_n938), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n924), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(KEYINPUT110), .A2(KEYINPUT41), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n918), .B2(new_n919), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT110), .B1(new_n942), .B2(new_n916), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n936), .A2(new_n949), .A3(new_n950), .A4(new_n940), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(new_n911), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n944), .A2(new_n952), .A3(new_n898), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT112), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n944), .A2(new_n952), .A3(new_n955), .A4(new_n898), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(KEYINPUT43), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n923), .B1(new_n945), .B2(new_n946), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n936), .A2(new_n920), .A3(new_n940), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n911), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(G37), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n944), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n963), .A2(KEYINPUT44), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n957), .A2(KEYINPUT113), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT113), .B1(new_n957), .B2(new_n964), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n944), .A2(new_n960), .A3(new_n962), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n944), .A2(new_n952), .A3(new_n961), .A4(new_n898), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n967), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI211_X1 g548(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n969), .C2(new_n970), .ZN(new_n974));
  OAI22_X1  g549(.A1(new_n965), .A2(new_n966), .B1(new_n973), .B2(new_n974), .ZN(G397));
  INV_X1    g550(.A(KEYINPUT125), .ZN(new_n976));
  NAND2_X1  g551(.A1(G286), .A2(G8), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT119), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n500), .A2(new_n504), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT71), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n505), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT50), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n888), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n985));
  INV_X1    g560(.A(new_n472), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n485), .A2(new_n486), .A3(G2105), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n486), .B1(new_n485), .B2(G2105), .ZN(new_n988));
  OAI211_X1 g563(.A(G40), .B(new_n986), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n984), .A2(new_n840), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  AOI21_X1  g567(.A(G1384), .B1(new_n500), .B2(new_n504), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n989), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n981), .A2(KEYINPUT45), .A3(new_n982), .A4(new_n505), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n821), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n978), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  NOR4_X1   g573(.A1(new_n506), .A2(new_n507), .A3(new_n992), .A4(G1384), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n992), .B1(new_n888), .B2(G1384), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(G160), .A3(G40), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n822), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n984), .A2(new_n840), .A3(new_n990), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(KEYINPUT119), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n977), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n998), .A2(G168), .A3(new_n1004), .ZN(new_n1006));
  INV_X1    g581(.A(G8), .ZN(new_n1007));
  NOR2_X1   g582(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1006), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1013));
  OAI21_X1  g588(.A(G8), .B1(new_n991), .B2(new_n997), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1005), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT62), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n976), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1006), .A2(new_n1011), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n1019), .C2(new_n1005), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n752), .A2(G1976), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT115), .B(G1976), .Z(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1025), .B(G8), .C1(new_n989), .C2(new_n994), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n483), .A2(new_n487), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1028), .A2(new_n993), .A3(G40), .A4(new_n986), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n1029), .B2(G8), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1022), .B(new_n1024), .C1(new_n1027), .C2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n585), .A2(new_n588), .A3(new_n693), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n519), .B1(new_n582), .B2(new_n583), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n586), .A2(new_n587), .ZN(new_n1034));
  OAI21_X1  g609(.A(G1981), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT116), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1032), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n989), .B2(new_n994), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT114), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1043), .A2(new_n1026), .B1(G1976), .B2(new_n752), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1031), .B(new_n1041), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G166), .A2(new_n1007), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT55), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n989), .B1(new_n983), .B2(new_n992), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n993), .A2(KEYINPUT45), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1971), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n984), .A2(new_n990), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G2090), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1049), .B(G8), .C1(new_n1052), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n981), .A2(new_n1056), .A3(new_n982), .A4(new_n505), .ZN(new_n1057));
  INV_X1    g632(.A(new_n989), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n994), .A2(KEYINPUT50), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(G2090), .ZN(new_n1061));
  OAI21_X1  g636(.A(G8), .B1(new_n1052), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1048), .B(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n983), .A2(new_n992), .ZN(new_n1066));
  INV_X1    g641(.A(G2078), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n1058), .A4(new_n1051), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  INV_X1    g644(.A(G1961), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1068), .A2(new_n1069), .B1(new_n1053), .B2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n995), .A2(KEYINPUT53), .A3(new_n1067), .A4(new_n996), .ZN(new_n1072));
  AOI21_X1  g647(.A(G301), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1047), .A2(new_n1055), .A3(new_n1065), .A4(new_n1073), .ZN(new_n1074));
  AOI211_X1 g649(.A(KEYINPUT124), .B(new_n1074), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1002), .A2(new_n1003), .A3(KEYINPUT119), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT119), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1077), .A2(new_n1078), .A3(G286), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1011), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1015), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1005), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1017), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1074), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1076), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1021), .B1(new_n1075), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT126), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n1088));
  NAND2_X1  g663(.A1(G299), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n568), .A2(new_n573), .A3(KEYINPUT57), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1050), .A2(new_n1051), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1956), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1060), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1091), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1029), .A2(G2067), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1053), .B2(new_n794), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(new_n611), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1093), .A2(new_n1091), .A3(new_n1095), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT117), .B(G1996), .Z(new_n1103));
  NAND4_X1  g678(.A1(new_n1066), .A2(new_n1058), .A3(new_n1051), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1029), .A2(new_n1106), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1105), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1102), .B1(new_n1110), .B2(new_n559), .ZN(new_n1111));
  NOR4_X1   g686(.A1(new_n1108), .A2(new_n1109), .A3(KEYINPUT59), .A4(new_n862), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1100), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1114), .B1(new_n1115), .B2(new_n1096), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n610), .B(new_n1097), .C1(new_n1053), .C2(new_n794), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT60), .B1(new_n1099), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1098), .A2(new_n1119), .A3(new_n610), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1091), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(KEYINPUT61), .A3(new_n1100), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1116), .A2(new_n1118), .A3(new_n1120), .A4(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1101), .B1(new_n1113), .B2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT122), .B(G2078), .Z(new_n1128));
  NAND4_X1  g703(.A1(new_n482), .A2(KEYINPUT53), .A3(G40), .A4(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1051), .A2(new_n1000), .A3(new_n986), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1071), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(G171), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1127), .B1(new_n1132), .B2(new_n1073), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1071), .A2(G301), .A3(new_n1072), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1131), .A2(G171), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1136), .A2(KEYINPUT54), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1047), .A2(new_n1055), .A3(new_n1065), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1016), .A2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1126), .A2(new_n1133), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1055), .A2(new_n1046), .ZN(new_n1143));
  INV_X1    g718(.A(G1976), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1041), .A2(new_n1144), .A3(new_n752), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1145), .A2(new_n1032), .B1(new_n1026), .B2(new_n1043), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1014), .A2(G286), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1140), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(G8), .B1(new_n1054), .B2(new_n1052), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1147), .B1(new_n1151), .B2(new_n1064), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1152), .A2(new_n1047), .A3(new_n1148), .A4(new_n1055), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1143), .B(new_n1146), .C1(new_n1150), .C2(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1142), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1021), .B(new_n1156), .C1(new_n1075), .C2(new_n1085), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1087), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n989), .A2(new_n1000), .ZN(new_n1159));
  INV_X1    g734(.A(G1996), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n741), .B(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n771), .A2(new_n774), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n801), .B(new_n804), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n773), .B2(new_n770), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(G1986), .B2(G290), .ZN(new_n1166));
  INV_X1    g741(.A(G290), .ZN(new_n1167));
  INV_X1    g742(.A(G1986), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1159), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1158), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1167), .A2(new_n1168), .A3(new_n1159), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT48), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1159), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n1174), .B2(new_n1165), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1163), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1159), .B1(new_n1176), .B2(new_n741), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT46), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1174), .B2(G1996), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1159), .A2(KEYINPUT46), .A3(new_n1160), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT47), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1183));
  OAI22_X1  g758(.A1(new_n1183), .A2(new_n1162), .B1(G2067), .B2(new_n801), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n1159), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1175), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1171), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g762(.A(G227), .ZN(new_n1189));
  NOR2_X1   g763(.A1(G229), .A2(new_n463), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n663), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g765(.A(new_n1191), .ZN(new_n1192));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n1193));
  AOI21_X1  g767(.A(new_n899), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n1191), .A2(KEYINPUT127), .ZN(new_n1195));
  AND3_X1   g769(.A1(new_n1194), .A2(new_n971), .A3(new_n1195), .ZN(G308));
  NAND3_X1  g770(.A1(new_n1194), .A2(new_n971), .A3(new_n1195), .ZN(G225));
endmodule


