//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT69), .B1(new_n187), .B2(G119), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT69), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n193), .A2(KEYINPUT68), .A3(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n194), .B1(new_n193), .B2(KEYINPUT68), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(G131), .B1(new_n199), .B2(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n205), .A3(new_n202), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n200), .A2(new_n205), .A3(KEYINPUT66), .A4(new_n202), .ZN(new_n209));
  AOI221_X4 g023(.A(KEYINPUT70), .B1(G131), .B2(new_n204), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(new_n209), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n204), .A2(G131), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT64), .A2(G146), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(G143), .A3(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT0), .B(G128), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT64), .A2(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT64), .A2(G146), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n221), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n221), .A2(G146), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n224), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n210), .A2(new_n214), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n219), .A2(new_n234), .A3(G128), .A4(new_n222), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT67), .B(G128), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n219), .B2(KEYINPUT1), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n217), .A2(new_n218), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n228), .B1(new_n238), .B2(new_n221), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n235), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n203), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n199), .A2(G137), .ZN(new_n242));
  OAI21_X1  g056(.A(G131), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n240), .A2(new_n212), .A3(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT30), .B1(new_n233), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n212), .A2(new_n213), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n223), .B2(new_n230), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n227), .A2(new_n229), .ZN(new_n249));
  INV_X1    g063(.A(new_n224), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(KEYINPUT65), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n246), .A2(new_n248), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n240), .A2(new_n212), .A3(new_n243), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n197), .B1(new_n245), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT71), .B(G237), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n256), .A2(new_n197), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n246), .A2(KEYINPUT70), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n212), .A2(new_n211), .A3(new_n213), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(new_n231), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT31), .B1(new_n258), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(new_n233), .B2(new_n265), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n254), .A2(new_n256), .ZN(new_n275));
  INV_X1    g089(.A(new_n197), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n266), .A2(new_n269), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n264), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n255), .B1(new_n269), .B2(new_n256), .ZN(new_n282));
  INV_X1    g096(.A(new_n257), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n270), .A4(new_n264), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n272), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(G472), .A2(G902), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT32), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n288), .ZN(new_n292));
  INV_X1    g106(.A(G472), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n264), .B(new_n274), .C1(new_n277), .C2(new_n278), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n210), .A2(new_n214), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n265), .B1(new_n296), .B2(new_n231), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n244), .B1(new_n296), .B2(new_n231), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n257), .B1(new_n298), .B2(new_n255), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n299), .B2(new_n276), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n294), .B(new_n295), .C1(new_n300), .C2(new_n264), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n297), .A2(KEYINPUT28), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n270), .B1(new_n298), .B2(new_n197), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n303), .B2(KEYINPUT28), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n280), .A2(new_n294), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI211_X1 g120(.A(KEYINPUT73), .B(new_n293), .C1(new_n301), .C2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n197), .B1(new_n269), .B2(new_n256), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT28), .B1(new_n310), .B2(new_n297), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n305), .A2(new_n311), .A3(new_n274), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n295), .A2(new_n294), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n264), .B1(new_n284), .B2(new_n270), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n309), .B(new_n312), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n308), .B1(new_n315), .B2(G472), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n291), .B(new_n292), .C1(new_n307), .C2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G217), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(G234), .B2(new_n309), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G125), .B(G140), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n321), .A2(KEYINPUT16), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G125), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(KEYINPUT16), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n216), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n325), .B1(new_n321), .B2(KEYINPUT16), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G146), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n236), .A2(KEYINPUT23), .A3(G119), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT75), .B1(new_n190), .B2(G128), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n332));
  INV_X1    g146(.A(G128), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(G119), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(G119), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n331), .B(new_n334), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G110), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n335), .B1(new_n236), .B2(G119), .ZN(new_n340));
  XOR2_X1   g154(.A(KEYINPUT24), .B(G110), .Z(new_n341));
  AOI21_X1  g155(.A(KEYINPUT74), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n341), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n329), .B(new_n339), .C1(new_n342), .C2(new_n345), .ZN(new_n346));
  OAI22_X1  g160(.A1(new_n338), .A2(G110), .B1(new_n340), .B2(new_n341), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n225), .A2(new_n226), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n327), .A2(G146), .B1(new_n349), .B2(new_n321), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n348), .B1(new_n347), .B2(new_n350), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n346), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT22), .B(G137), .ZN(new_n354));
  INV_X1    g168(.A(G953), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(G221), .A3(G234), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n354), .B(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n346), .B(new_n357), .C1(new_n351), .C2(new_n352), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n309), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n320), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n360), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n319), .A2(G902), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n365), .A2(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT9), .B(G234), .ZN(new_n371));
  OAI21_X1  g185(.A(G221), .B1(new_n371), .B2(G902), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n372), .B(KEYINPUT78), .Z(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G110), .B(G140), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n355), .A2(G227), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G104), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT3), .B1(new_n379), .B2(G107), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G104), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(G107), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n380), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n379), .A2(G107), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n382), .A2(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n234), .B1(G143), .B2(new_n216), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n333), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT1), .B1(new_n221), .B2(G146), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT80), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n394), .A2(new_n396), .B1(new_n219), .B2(new_n222), .ZN(new_n397));
  INV_X1    g211(.A(new_n235), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n391), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT10), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n240), .A2(KEYINPUT10), .A3(new_n391), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n380), .A2(new_n383), .A3(new_n385), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G101), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT4), .A3(new_n386), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT79), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n403), .A2(KEYINPUT79), .A3(new_n406), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n231), .B(new_n405), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n401), .A2(new_n402), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n378), .B1(new_n410), .B2(new_n296), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n267), .A2(new_n268), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n414), .A2(new_n401), .A3(new_n402), .A4(new_n409), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT82), .A3(new_n378), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n219), .A2(new_n222), .ZN(new_n417));
  INV_X1    g231(.A(new_n396), .ZN(new_n418));
  OAI21_X1  g232(.A(G128), .B1(new_n395), .B2(KEYINPUT80), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n390), .B1(new_n420), .B2(new_n235), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n390), .B(new_n235), .C1(new_n237), .C2(new_n239), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n267), .B(new_n268), .C1(new_n421), .C2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT12), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n425), .B1(new_n212), .B2(new_n213), .ZN(new_n427));
  OAI211_X1 g241(.A(KEYINPUT81), .B(new_n427), .C1(new_n423), .C2(new_n421), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n423), .B2(new_n421), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n426), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n413), .A2(new_n416), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n410), .A2(new_n296), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n410), .A2(new_n296), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n377), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI211_X1 g251(.A(G469), .B(G902), .C1(new_n433), .C2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n415), .A3(new_n378), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n424), .A2(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n436), .B1(new_n440), .B2(new_n428), .ZN(new_n441));
  OAI211_X1 g255(.A(G469), .B(new_n439), .C1(new_n441), .C2(new_n378), .ZN(new_n442));
  NAND2_X1  g256(.A1(G469), .A2(G902), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n374), .B1(new_n438), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n188), .A2(new_n191), .A3(KEYINPUT5), .A4(new_n192), .ZN(new_n446));
  INV_X1    g260(.A(G113), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n187), .A2(G119), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT5), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n193), .A2(new_n194), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n446), .A2(KEYINPUT83), .A3(new_n450), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n453), .A2(new_n391), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(new_n197), .ZN(new_n459));
  XNOR2_X1  g273(.A(G110), .B(G122), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n457), .B(new_n460), .C1(new_n458), .C2(new_n197), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(KEYINPUT6), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(new_n465), .A3(new_n461), .ZN(new_n466));
  INV_X1    g280(.A(G125), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n240), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n251), .A2(G125), .A3(new_n252), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n355), .A2(G224), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n464), .A2(new_n466), .A3(new_n472), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n446), .A2(KEYINPUT84), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n190), .A2(G116), .ZN(new_n475));
  OAI21_X1  g289(.A(G113), .B1(new_n475), .B2(KEYINPUT5), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n476), .B1(new_n446), .B2(KEYINPUT84), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT85), .B1(new_n478), .B2(new_n455), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT85), .ZN(new_n480));
  AOI211_X1 g294(.A(new_n480), .B(new_n454), .C1(new_n474), .C2(new_n477), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n391), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n460), .B(KEYINPUT8), .Z(new_n483));
  AND3_X1   g297(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n390), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n471), .A2(KEYINPUT7), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n468), .A2(new_n469), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT86), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n468), .B2(new_n469), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n487), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n234), .B1(new_n349), .B2(G143), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n249), .B1(new_n494), .B2(new_n236), .ZN(new_n495));
  AOI21_X1  g309(.A(G125), .B1(new_n495), .B2(new_n235), .ZN(new_n496));
  INV_X1    g310(.A(new_n469), .ZN(new_n497));
  OAI211_X1 g311(.A(KEYINPUT86), .B(new_n493), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n486), .A2(new_n492), .A3(new_n463), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n473), .A2(new_n499), .A3(new_n309), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n473), .A2(new_n499), .A3(new_n309), .A4(new_n501), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G214), .B1(G237), .B2(G902), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n445), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n236), .A2(G143), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n221), .A2(G128), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT13), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT90), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n510), .B2(new_n511), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n514), .B(G134), .C1(new_n513), .C2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(G116), .B(G122), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n382), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n509), .A2(new_n199), .A3(new_n510), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n509), .A2(new_n510), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G134), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n520), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT14), .ZN(new_n526));
  INV_X1    g340(.A(G122), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(G116), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n518), .B1(new_n528), .B2(new_n382), .ZN(new_n529));
  OR3_X1    g343(.A1(new_n518), .A2(new_n528), .A3(new_n382), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n371), .A2(new_n318), .A3(G953), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n522), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n532), .B1(new_n522), .B2(new_n531), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n309), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G478), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(KEYINPUT15), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n536), .B(new_n542), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT20), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT71), .B(G237), .Z(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(G214), .A3(new_n355), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(new_n221), .ZN(new_n548));
  AOI21_X1  g362(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n549));
  OAI21_X1  g363(.A(G131), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n221), .ZN(new_n552));
  INV_X1    g366(.A(G131), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(KEYINPUT17), .B(G131), .C1(new_n548), .C2(new_n549), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT89), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n329), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n556), .A2(new_n559), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(G113), .B(G122), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(new_n379), .ZN(new_n565));
  OAI211_X1 g379(.A(KEYINPUT18), .B(G131), .C1(new_n548), .C2(new_n549), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n349), .A2(new_n321), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n216), .B2(new_n321), .ZN(new_n568));
  NAND2_X1  g382(.A1(KEYINPUT18), .A2(G131), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n552), .A2(new_n554), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n566), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n563), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT88), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT87), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT19), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n321), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n576), .B1(new_n321), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n573), .B1(new_n578), .B2(new_n238), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n321), .A2(new_n577), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n580), .A2(KEYINPUT88), .A3(new_n349), .A4(new_n576), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n555), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n582), .B(new_n328), .C1(new_n583), .C2(new_n561), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n571), .ZN(new_n585));
  INV_X1    g399(.A(new_n565), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n572), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(G475), .A2(G902), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n545), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n589), .ZN(new_n591));
  AOI211_X1 g405(.A(KEYINPUT20), .B(new_n591), .C1(new_n572), .C2(new_n587), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n563), .A2(new_n571), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n586), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n594), .B2(new_n572), .ZN(new_n595));
  INV_X1    g409(.A(G475), .ZN(new_n596));
  OAI22_X1  g410(.A1(new_n590), .A2(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(G234), .A2(G237), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n598), .A2(G952), .A3(new_n355), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT21), .B(G898), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT92), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n598), .A2(G902), .A3(G953), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n544), .A2(new_n597), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n317), .A2(new_n370), .A3(new_n508), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  AND2_X1   g421(.A1(new_n442), .A2(new_n443), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n433), .A2(new_n437), .ZN(new_n609));
  INV_X1    g423(.A(G469), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n309), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n373), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n370), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n287), .A2(new_n309), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n615), .A2(G472), .B1(new_n288), .B2(new_n287), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n604), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT94), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n621), .B(new_n622), .C1(new_n534), .C2(new_n535), .ZN(new_n623));
  INV_X1    g437(.A(new_n535), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n624), .A2(new_n619), .A3(new_n620), .A4(new_n533), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n537), .A2(G902), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n536), .A2(new_n537), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n597), .A2(new_n618), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n506), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n309), .A2(new_n473), .A3(new_n499), .A4(new_n501), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(KEYINPUT93), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT93), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n503), .A2(new_n635), .A3(new_n504), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n617), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n597), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n618), .A3(new_n544), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n637), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n617), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  AND3_X1   g461(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT25), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT25), .B1(new_n361), .B2(new_n362), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n648), .A2(new_n649), .A3(new_n320), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n358), .A2(KEYINPUT36), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n353), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n353), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n652), .A2(new_n369), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT95), .B1(new_n650), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n363), .A2(new_n364), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n366), .A3(new_n319), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT95), .ZN(new_n658));
  INV_X1    g472(.A(new_n654), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n661), .A2(new_n508), .A3(new_n605), .A4(new_n616), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  AOI21_X1  g478(.A(new_n445), .B1(new_n655), .B2(new_n660), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n506), .B1(new_n504), .B2(new_n635), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n490), .B1(KEYINPUT86), .B2(new_n488), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n498), .A2(new_n463), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(G902), .B1(new_n669), .B2(new_n486), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n501), .B1(new_n670), .B2(new_n473), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n633), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n666), .B1(new_n672), .B2(new_n635), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n599), .B1(new_n603), .B2(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n597), .A2(new_n543), .A3(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n317), .A2(new_n665), .A3(new_n673), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XOR2_X1   g492(.A(new_n675), .B(KEYINPUT39), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n612), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT40), .Z(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT96), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(KEYINPUT96), .ZN(new_n683));
  INV_X1    g497(.A(new_n661), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n505), .B(KEYINPUT38), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n506), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n300), .A2(new_n280), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n309), .B1(new_n303), .B2(new_n264), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n291), .A2(new_n292), .A3(new_n689), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n590), .A2(new_n592), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n595), .A2(new_n596), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n543), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n682), .A2(new_n683), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G143), .ZN(G45));
  AOI22_X1  g511(.A1(new_n626), .A2(new_n627), .B1(new_n537), .B2(new_n536), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n642), .A2(new_n698), .A3(new_n675), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n317), .A2(new_n665), .A3(new_n673), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  NAND2_X1  g515(.A1(new_n609), .A2(new_n309), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(G469), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n374), .A3(new_n611), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n317), .A2(new_n370), .A3(new_n638), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  INV_X1    g522(.A(new_n370), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n307), .A2(new_n316), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n291), .A2(new_n292), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n644), .A3(new_n705), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NOR2_X1   g528(.A1(new_n704), .A2(new_n637), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n317), .A2(new_n605), .A3(new_n715), .A4(new_n661), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  XOR2_X1   g531(.A(KEYINPUT97), .B(G472), .Z(new_n718));
  OAI211_X1 g532(.A(new_n272), .B(new_n286), .C1(new_n264), .C2(new_n304), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n615), .A2(new_n718), .B1(new_n288), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n720), .A2(new_n370), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n637), .A2(new_n642), .A3(new_n543), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n618), .A3(new_n705), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT98), .B(G122), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G24));
  NAND4_X1  g539(.A1(new_n715), .A2(new_n661), .A3(new_n699), .A4(new_n720), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  INV_X1    g541(.A(KEYINPUT99), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n439), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n434), .A2(new_n415), .A3(KEYINPUT99), .A4(new_n378), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n729), .B(new_n730), .C1(new_n441), .C2(new_n378), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n610), .B1(new_n731), .B2(new_n309), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n374), .B1(new_n732), .B2(new_n438), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n672), .A2(new_n506), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT100), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n733), .A2(new_n734), .A3(KEYINPUT100), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n699), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n292), .B(KEYINPUT101), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n291), .B1(new_n307), .B2(new_n316), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n370), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT42), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n737), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n735), .ZN(new_n744));
  INV_X1    g558(.A(new_n699), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(KEYINPUT42), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n712), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n553), .ZN(G33));
  NAND3_X1  g563(.A1(new_n744), .A2(new_n712), .A3(new_n676), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  INV_X1    g565(.A(KEYINPUT103), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n698), .B1(new_n597), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n752), .B2(new_n597), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT43), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT43), .B1(new_n630), .B2(KEYINPUT102), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT102), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n698), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n642), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n761), .A2(new_n616), .A3(new_n684), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n734), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OR4_X1    g578(.A1(new_n763), .A2(new_n761), .A3(new_n616), .A4(new_n684), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT104), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n731), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n439), .B1(new_n441), .B2(new_n378), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n769), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(G469), .A3(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n443), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n443), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n611), .A3(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n777), .A2(new_n374), .A3(new_n679), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n764), .A2(KEYINPUT104), .A3(new_n765), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n768), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT105), .B(G137), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G39));
  NAND2_X1  g596(.A1(new_n777), .A2(new_n374), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n777), .A2(KEYINPUT47), .A3(new_n374), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n317), .A2(new_n745), .A3(new_n370), .A4(new_n734), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT106), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NAND3_X1  g605(.A1(new_n370), .A2(new_n374), .A3(new_n506), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n703), .A2(new_n611), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n792), .B1(KEYINPUT49), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(KEYINPUT49), .B2(new_n793), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n795), .A2(new_n690), .A3(new_n685), .A4(new_n754), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n698), .B1(new_n691), .B2(new_n692), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n672), .A2(new_n632), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT107), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .A4(new_n618), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT107), .B1(new_n631), .B2(new_n507), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n614), .A2(new_n801), .A3(new_n616), .A4(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n723), .A2(new_n803), .A3(new_n716), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n643), .A2(new_n507), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n614), .A2(new_n805), .A3(new_n616), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n606), .A2(new_n806), .A3(new_n662), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n804), .A2(new_n807), .A3(new_n706), .A4(new_n713), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n661), .A2(new_n720), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n744), .A2(new_n699), .A3(new_n809), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n734), .A2(new_n544), .A3(new_n597), .A4(new_n675), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n317), .A3(new_n665), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n750), .A3(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n808), .A2(new_n748), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT109), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n611), .B(new_n443), .C1(new_n610), .C2(new_n731), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n654), .B(new_n675), .C1(new_n365), .C2(new_n366), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n673), .A2(new_n816), .A3(new_n817), .A4(new_n374), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT108), .B1(new_n694), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n675), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n657), .A2(new_n659), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n733), .A2(new_n637), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT108), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(new_n823), .A3(new_n690), .A4(new_n693), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n677), .A2(new_n700), .A3(new_n726), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n825), .A2(new_n826), .A3(KEYINPUT52), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n677), .A2(new_n700), .A3(new_n726), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n819), .A2(new_n824), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n815), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT52), .B1(new_n825), .B2(new_n826), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n677), .A2(new_n700), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n830), .A3(new_n828), .A4(new_n726), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n835), .A3(KEYINPUT109), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n814), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT110), .B1(new_n827), .B2(new_n831), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n833), .A2(new_n835), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(KEYINPUT53), .A3(new_n814), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT54), .ZN(new_n846));
  INV_X1    g660(.A(new_n721), .ZN(new_n847));
  INV_X1    g661(.A(new_n599), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT111), .B1(new_n761), .B2(new_n848), .ZN(new_n849));
  AOI22_X1  g663(.A1(KEYINPUT43), .A2(new_n754), .B1(new_n759), .B2(new_n642), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n599), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n847), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n685), .A2(new_n506), .A3(new_n704), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n849), .A2(new_n852), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n704), .A2(new_n734), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n809), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n690), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n370), .A2(new_n861), .A3(new_n599), .A4(new_n859), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n642), .A3(new_n698), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n847), .B(new_n734), .C1(new_n849), .C2(new_n852), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n793), .B(KEYINPUT112), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n373), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT113), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n785), .A2(new_n786), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n864), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT51), .B1(new_n857), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n853), .A2(new_n715), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n862), .A2(new_n798), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(G952), .A3(new_n355), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n741), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n858), .A2(new_n875), .A3(new_n859), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n876), .A2(KEYINPUT48), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(KEYINPUT48), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n833), .A2(KEYINPUT109), .A3(new_n835), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT109), .B1(new_n833), .B2(new_n835), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n808), .A2(new_n748), .A3(new_n813), .A4(new_n838), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT54), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n833), .A2(new_n841), .A3(new_n835), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n841), .B1(new_n833), .B2(new_n835), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n814), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n838), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n867), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n865), .B1(new_n787), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n864), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n857), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AND4_X1   g710(.A1(new_n846), .A2(new_n881), .A3(new_n891), .A4(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(G952), .A2(G953), .ZN(new_n898));
  OAI211_X1 g712(.A(KEYINPUT114), .B(new_n797), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT114), .ZN(new_n900));
  INV_X1    g714(.A(new_n896), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n901), .A2(new_n871), .A3(new_n880), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n845), .A2(KEYINPUT54), .B1(new_n890), .B2(new_n886), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n900), .B1(new_n904), .B2(new_n796), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n899), .A2(new_n905), .ZN(G75));
  INV_X1    g720(.A(KEYINPUT116), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n889), .A2(new_n838), .B1(new_n884), .B2(new_n885), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n907), .B1(new_n908), .B2(new_n309), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT53), .B1(new_n843), .B2(new_n814), .ZN(new_n910));
  INV_X1    g724(.A(new_n748), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n712), .A2(new_n644), .A3(new_n705), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n606), .A2(new_n706), .A3(new_n806), .A4(new_n662), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n723), .A2(new_n803), .A3(new_n716), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n813), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n911), .A2(new_n915), .A3(new_n916), .A4(KEYINPUT53), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n917), .A2(new_n882), .A3(new_n883), .ZN(new_n918));
  OAI211_X1 g732(.A(KEYINPUT116), .B(G902), .C1(new_n910), .C2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n909), .A2(new_n502), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n464), .A2(new_n466), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(new_n472), .Z(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT55), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(KEYINPUT56), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n355), .A2(G952), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT117), .Z(new_n927));
  OAI211_X1 g741(.A(G210), .B(G902), .C1(new_n910), .C2(new_n918), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT56), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT115), .B1(new_n930), .B2(new_n923), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT115), .ZN(new_n932));
  INV_X1    g746(.A(new_n923), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n932), .B(new_n933), .C1(new_n928), .C2(new_n929), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n925), .B(new_n927), .C1(new_n931), .C2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(G51));
  INV_X1    g750(.A(KEYINPUT118), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n814), .A2(new_n832), .A3(KEYINPUT53), .A4(new_n836), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT54), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n937), .B1(new_n940), .B2(new_n910), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n886), .A2(new_n890), .A3(KEYINPUT118), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n941), .B(new_n942), .C1(new_n939), .C2(new_n908), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n443), .B(KEYINPUT57), .Z(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n609), .ZN(new_n946));
  INV_X1    g760(.A(new_n773), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n909), .A2(new_n947), .A3(new_n919), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n926), .B1(new_n946), .B2(new_n948), .ZN(G54));
  AND2_X1   g763(.A1(KEYINPUT58), .A2(G475), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n909), .A2(new_n919), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n572), .A3(new_n587), .ZN(new_n952));
  INV_X1    g766(.A(new_n926), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n909), .A2(new_n588), .A3(new_n919), .A4(new_n950), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G60));
  INV_X1    g769(.A(new_n626), .ZN(new_n956));
  NAND2_X1  g770(.A1(G478), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT59), .Z(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n903), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT119), .ZN(new_n960));
  INV_X1    g774(.A(new_n927), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n956), .A2(new_n958), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(new_n943), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT119), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n964), .B(new_n956), .C1(new_n903), .C2(new_n958), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n960), .A2(new_n963), .A3(new_n965), .ZN(G63));
  NAND2_X1  g780(.A1(new_n652), .A2(new_n653), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n318), .A2(new_n309), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n968), .B(new_n971), .C1(new_n910), .C2(new_n918), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT121), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n973), .A3(new_n927), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT61), .ZN(new_n975));
  INV_X1    g789(.A(new_n971), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n367), .B1(new_n908), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n977), .A2(new_n927), .A3(new_n972), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n975), .B(new_n978), .ZN(G66));
  AOI21_X1  g793(.A(new_n355), .B1(new_n601), .B2(G224), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT123), .Z(new_n981));
  XNOR2_X1  g795(.A(new_n915), .B(KEYINPUT122), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(G953), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n921), .B1(G898), .B2(new_n355), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT124), .Z(new_n985));
  XNOR2_X1  g799(.A(new_n983), .B(new_n985), .ZN(G69));
  AOI21_X1  g800(.A(new_n355), .B1(G227), .B2(G900), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n299), .B(new_n578), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n674), .B2(new_n355), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n778), .A2(new_n722), .A3(new_n875), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n790), .A2(new_n991), .A3(new_n911), .A4(new_n750), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n780), .A2(new_n829), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT125), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n780), .A2(KEYINPUT125), .A3(new_n829), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n990), .B1(new_n997), .B2(new_n355), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n696), .A2(new_n829), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n798), .B1(new_n544), .B2(new_n642), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n1002), .A2(new_n680), .A3(new_n734), .ZN(new_n1003));
  AOI22_X1  g817(.A1(new_n787), .A2(new_n789), .B1(new_n712), .B2(new_n1003), .ZN(new_n1004));
  AND4_X1   g818(.A1(new_n780), .A2(new_n1000), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n988), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n987), .B1(new_n998), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n987), .ZN(new_n1009));
  AOI211_X1 g823(.A(G953), .B(new_n992), .C1(new_n995), .C2(new_n996), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n1009), .B(new_n1006), .C1(new_n1010), .C2(new_n990), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1008), .A2(new_n1011), .ZN(G72));
  NAND2_X1  g826(.A1(new_n300), .A2(new_n280), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT126), .Z(new_n1014));
  NAND2_X1  g828(.A1(new_n995), .A2(new_n996), .ZN(new_n1015));
  INV_X1    g829(.A(new_n992), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1015), .A2(new_n982), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  AOI21_X1  g833(.A(new_n1014), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n687), .ZN(new_n1021));
  AND4_X1   g835(.A1(new_n1021), .A2(new_n845), .A3(new_n1019), .A4(new_n1013), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1019), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1023), .B1(new_n1005), .B2(new_n982), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n953), .B1(new_n1024), .B2(new_n1021), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n1020), .A2(new_n1022), .A3(new_n1025), .ZN(G57));
endmodule


