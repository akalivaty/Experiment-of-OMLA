//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1249, new_n1250, new_n1251;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G68), .B2(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G107), .ZN(new_n216));
  INV_X1    g0016(.A(G264), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  INV_X1    g0029(.A(G13), .ZN(new_n230));
  OAI21_X1  g0030(.A(KEYINPUT64), .B1(new_n203), .B2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(KEYINPUT64), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n232), .A2(G1), .A3(G13), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n235), .A2(new_n204), .ZN(new_n236));
  OAI21_X1  g0036(.A(G50), .B1(G58), .B2(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT65), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(new_n239));
  AOI211_X1 g0039(.A(new_n209), .B(new_n229), .C1(new_n236), .C2(new_n239), .ZN(G361));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n217), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT66), .ZN(new_n250));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  NOR2_X1   g0056(.A1(new_n230), .A2(G1), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n204), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n220), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n205), .A2(G33), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(new_n231), .A3(new_n233), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n203), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G50), .A3(new_n264), .ZN(new_n265));
  NOR3_X1   g0065(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT68), .B1(new_n266), .B2(new_n204), .ZN(new_n267));
  INV_X1    g0067(.A(G68), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n220), .A2(new_n225), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G20), .ZN(new_n273));
  OR2_X1    g0073(.A1(KEYINPUT8), .A2(G58), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT8), .A2(G58), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G150), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n267), .A2(new_n271), .A3(new_n276), .A4(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT69), .ZN(new_n280));
  AND3_X1   g0080(.A1(new_n279), .A2(new_n280), .A3(new_n262), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(new_n279), .B2(new_n262), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n260), .B(new_n265), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT70), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT9), .ZN(new_n285));
  AND3_X1   g0085(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n284), .B1(new_n283), .B2(new_n285), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n234), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n222), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n290), .A2(new_n292), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G222), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G223), .A2(G1698), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n289), .A2(new_n294), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT67), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n203), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n303), .B1(new_n308), .B2(new_n221), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G190), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n286), .A2(new_n287), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n283), .A2(new_n285), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(G200), .B1(new_n300), .B2(new_n309), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT71), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(KEYINPUT71), .B(G200), .C1(new_n300), .C2(new_n309), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n313), .A2(new_n314), .A3(new_n316), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n317), .ZN(new_n323));
  INV_X1    g0123(.A(new_n283), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(KEYINPUT9), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n283), .A2(new_n285), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT70), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n325), .A2(new_n327), .A3(new_n311), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT10), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G179), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n310), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G169), .B2(new_n310), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n324), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n273), .A2(G77), .B1(G20), .B2(new_n268), .ZN(new_n337));
  INV_X1    g0137(.A(new_n277), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n220), .B2(new_n338), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n339), .A2(new_n262), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n340), .A2(KEYINPUT11), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(KEYINPUT11), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n257), .A2(G20), .A3(new_n268), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT12), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n262), .B1(new_n203), .B2(G20), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G68), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n341), .A2(new_n342), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n226), .A2(G1698), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(G226), .B2(G1698), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n351), .B2(new_n293), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n303), .A2(KEYINPUT72), .ZN(new_n353));
  OR3_X1    g0153(.A1(new_n301), .A2(KEYINPUT72), .A3(new_n302), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n289), .A2(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n308), .A2(KEYINPUT73), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT73), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n305), .A2(new_n357), .A3(new_n307), .A4(new_n306), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(G238), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n361));
  NAND2_X1  g0161(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n355), .A2(new_n362), .A3(new_n359), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(G190), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n355), .A2(KEYINPUT13), .A3(new_n359), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(G200), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n348), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n366), .A2(new_n367), .A3(G169), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n361), .A2(G179), .A3(new_n363), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT14), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n366), .A2(new_n367), .A3(new_n374), .A4(G169), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n370), .B1(new_n376), .B2(new_n347), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n345), .A2(G77), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n259), .A2(new_n222), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n274), .A2(new_n275), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n380), .A2(new_n338), .B1(new_n204), .B2(new_n222), .ZN(new_n381));
  XOR2_X1   g0181(.A(KEYINPUT15), .B(G87), .Z(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n273), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n378), .B(new_n379), .C1(new_n263), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G238), .A2(G1698), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n295), .B(new_n385), .C1(new_n226), .C2(G1698), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n289), .B(new_n386), .C1(G107), .C2(new_n295), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G244), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n303), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n384), .B1(G190), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(G200), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n331), .A2(new_n336), .A3(new_n377), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G58), .A2(G68), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n397), .B(new_n398), .C1(G58), .C2(G68), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(G20), .B1(G159), .B2(new_n277), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n293), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n290), .A2(new_n292), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n403), .B1(new_n290), .B2(new_n292), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n204), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n402), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT16), .B(new_n400), .C1(new_n408), .C2(new_n268), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n399), .A2(G20), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n277), .A2(G159), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n407), .B1(new_n295), .B2(G20), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n268), .B1(new_n414), .B2(new_n401), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n410), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n409), .A2(new_n262), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n380), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n264), .ZN(new_n419));
  XOR2_X1   g0219(.A(new_n419), .B(KEYINPUT77), .Z(new_n420));
  NOR2_X1   g0220(.A1(new_n262), .A2(new_n259), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n420), .A2(new_n421), .B1(new_n380), .B2(new_n259), .ZN(new_n422));
  AND2_X1   g0222(.A1(G226), .A2(G1698), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n290), .A2(new_n292), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT78), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT78), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n290), .A2(new_n292), .A3(new_n423), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G87), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n290), .A2(new_n292), .A3(G223), .A4(new_n296), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n425), .A2(new_n427), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n289), .ZN(new_n431));
  INV_X1    g0231(.A(new_n303), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n388), .B2(G232), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G169), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n431), .A2(G179), .A3(new_n433), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n417), .A2(new_n422), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT18), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  INV_X1    g0239(.A(G190), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n431), .A2(new_n440), .A3(new_n433), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT79), .ZN(new_n442));
  INV_X1    g0242(.A(G200), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT79), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n431), .A2(new_n433), .A3(new_n445), .A4(new_n440), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n442), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(new_n417), .A3(new_n422), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT80), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT80), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n447), .A2(new_n450), .A3(new_n417), .A4(new_n422), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n439), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n448), .A2(KEYINPUT17), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n438), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n391), .A2(new_n332), .ZN(new_n455));
  INV_X1    g0255(.A(G169), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n390), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n384), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n395), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT5), .B(G41), .ZN(new_n461));
  INV_X1    g0261(.A(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G1), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G257), .A3(new_n307), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n461), .A2(G274), .A3(new_n463), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n465), .A2(KEYINPUT81), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT81), .B1(new_n465), .B2(new_n466), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n295), .A2(KEYINPUT4), .A3(G244), .A4(new_n296), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT4), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n293), .B2(new_n223), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n295), .A2(G250), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n296), .B1(new_n475), .B2(KEYINPUT4), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n289), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n469), .A2(G190), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n272), .A2(G1), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n262), .A2(new_n259), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G97), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n259), .A2(new_n212), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n216), .B1(new_n414), .B2(new_n401), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n338), .A2(new_n222), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT6), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n212), .A2(new_n216), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G97), .A2(G107), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n216), .A2(KEYINPUT6), .A3(G97), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n204), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n483), .A2(new_n484), .A3(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n481), .B(new_n482), .C1(new_n491), .C2(new_n263), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n443), .B1(new_n469), .B2(new_n477), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n478), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n469), .A2(G179), .A3(new_n477), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n456), .B1(new_n469), .B2(new_n477), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT82), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n492), .B(KEYINPUT82), .C1(new_n495), .C2(new_n496), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n494), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n290), .A2(new_n292), .A3(new_n204), .A4(G87), .ZN(new_n502));
  NOR2_X1   g0302(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n216), .A2(G20), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT23), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n505), .B(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  XOR2_X1   g0308(.A(KEYINPUT84), .B(KEYINPUT22), .Z(new_n509));
  NAND4_X1  g0309(.A1(new_n295), .A2(new_n509), .A3(new_n204), .A4(G87), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT24), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n508), .A2(new_n510), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n510), .A2(new_n512), .A3(new_n504), .A4(new_n507), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT24), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n262), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n480), .A2(G107), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n258), .A2(new_n505), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n519), .B(KEYINPUT25), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n464), .A2(new_n307), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G264), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n211), .A2(new_n296), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n213), .A2(G1698), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n290), .A2(new_n524), .A3(new_n292), .A4(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G294), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n272), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n289), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT85), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n523), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n289), .A2(new_n528), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n466), .B1(new_n532), .B2(KEYINPUT85), .ZN(new_n533));
  OAI21_X1  g0333(.A(G169), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n523), .A2(new_n532), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(G179), .A3(new_n466), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n521), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n523), .A2(new_n532), .A3(new_n466), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n443), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n532), .A2(KEYINPUT85), .B1(G264), .B2(new_n522), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n529), .A2(new_n530), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(new_n466), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n540), .B1(new_n543), .B2(G190), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n516), .A2(new_n262), .B1(G107), .B2(new_n480), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(new_n520), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n487), .A2(new_n210), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n349), .A2(new_n204), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(KEYINPUT19), .A3(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n290), .A2(new_n292), .A3(new_n204), .A4(G68), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n349), .A2(G20), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n549), .B(new_n550), .C1(KEYINPUT19), .C2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n382), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n552), .A2(new_n262), .B1(new_n259), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n479), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n421), .A2(new_n382), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n463), .A2(new_n302), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n211), .B1(new_n462), .B2(G1), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n307), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n223), .A2(G1698), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(G238), .B2(G1698), .ZN(new_n562));
  INV_X1    g0362(.A(G116), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n562), .A2(new_n293), .B1(new_n272), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n234), .A2(new_n288), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n456), .ZN(new_n568));
  INV_X1    g0368(.A(new_n560), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n289), .B2(new_n564), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n332), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n557), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n567), .A2(new_n440), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n480), .A2(G87), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n574), .B(new_n554), .C1(new_n443), .C2(new_n570), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n573), .B1(new_n575), .B2(KEYINPUT83), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n567), .A2(G200), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT83), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(new_n554), .A4(new_n574), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n572), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n538), .A2(new_n546), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n563), .A2(G20), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n471), .B(new_n204), .C1(G33), .C2(new_n212), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n262), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT20), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n258), .A2(new_n204), .A3(G116), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NOR4_X1   g0390(.A1(new_n262), .A2(new_n259), .A3(new_n563), .A4(new_n479), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n588), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G264), .A2(G1698), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n295), .B(new_n594), .C1(new_n213), .C2(G1698), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n289), .B(new_n595), .C1(G303), .C2(new_n295), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n522), .A2(G270), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n466), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(new_n332), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n589), .B(new_n591), .C1(new_n586), .C2(new_n587), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(G169), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n593), .A2(KEYINPUT21), .A3(G169), .A4(new_n598), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n598), .A2(new_n440), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n598), .A2(G200), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n602), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n600), .A2(new_n604), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n460), .A2(new_n501), .A3(new_n581), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT86), .ZN(G372));
  AND3_X1   g0411(.A1(new_n604), .A2(new_n605), .A3(new_n600), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n538), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n574), .A2(new_n554), .ZN(new_n614));
  XOR2_X1   g0414(.A(new_n614), .B(KEYINPUT87), .Z(new_n615));
  AOI21_X1  g0415(.A(new_n573), .B1(G200), .B2(new_n567), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n613), .A2(new_n501), .A3(new_n546), .A4(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n492), .ZN(new_n619));
  OR3_X1    g0419(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT88), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT88), .B1(new_n495), .B2(new_n496), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n572), .B1(new_n615), .B2(new_n616), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n572), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n499), .A2(new_n500), .A3(new_n580), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT26), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n618), .A2(new_n625), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n460), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g0430(.A(new_n630), .B(KEYINPUT89), .Z(new_n631));
  NOR2_X1   g0431(.A1(new_n452), .A2(new_n453), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n376), .A2(new_n347), .B1(new_n369), .B2(new_n459), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n438), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n335), .B1(new_n634), .B2(new_n331), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n631), .A2(new_n635), .ZN(G369));
  INV_X1    g0436(.A(new_n612), .ZN(new_n637));
  OR3_X1    g0437(.A1(new_n258), .A2(KEYINPUT27), .A3(G20), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT27), .B1(new_n258), .B2(G20), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(G213), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(G343), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n637), .A2(new_n593), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n642), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n609), .B1(new_n602), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G330), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n538), .A2(new_n546), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n521), .A2(new_n642), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n538), .B2(new_n644), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n521), .A2(new_n537), .A3(new_n644), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n612), .A2(new_n642), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n650), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(G399));
  INV_X1    g0458(.A(new_n207), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n547), .A2(G116), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G1), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n237), .B2(new_n661), .ZN(new_n664));
  XOR2_X1   g0464(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n665));
  XNOR2_X1  g0465(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n622), .A2(new_n624), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT26), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n627), .A2(KEYINPUT26), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n618), .A3(new_n626), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n644), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT29), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n629), .A2(new_n644), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n672), .B1(KEYINPUT29), .B2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n501), .A2(new_n581), .A3(new_n609), .A4(new_n644), .ZN(new_n675));
  INV_X1    g0475(.A(new_n468), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n465), .A2(KEYINPUT81), .A3(new_n466), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n477), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(new_n599), .A3(new_n535), .A4(new_n570), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT30), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n678), .A2(G179), .ZN(new_n682));
  AND4_X1   g0482(.A1(new_n539), .A2(new_n682), .A3(new_n567), .A4(new_n598), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n642), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n675), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT31), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n686), .B(new_n642), .C1(new_n681), .C2(new_n683), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n674), .B1(G330), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n666), .B1(new_n689), .B2(G1), .ZN(G364));
  NAND2_X1  g0490(.A1(new_n204), .A2(G13), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT91), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n203), .B1(new_n693), .B2(G45), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n660), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n646), .A2(G330), .ZN(new_n697));
  OR3_X1    g0497(.A1(new_n649), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(G13), .A2(G33), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G20), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n647), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n207), .A2(new_n295), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT92), .Z(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G355), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n252), .A2(new_n462), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n404), .A2(new_n405), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n659), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(G45), .B2(new_n238), .ZN(new_n709));
  OAI221_X1 g0509(.A(new_n705), .B1(G116), .B2(new_n207), .C1(new_n706), .C2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n235), .B1(G20), .B2(new_n456), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n701), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n443), .A2(G179), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n715), .A2(new_n204), .A3(new_n440), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G303), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n440), .A2(G20), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT93), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n721), .A2(G179), .A3(G200), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n204), .A2(new_n332), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G190), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n443), .ZN(new_n725));
  XOR2_X1   g0525(.A(KEYINPUT95), .B(G326), .Z(new_n726));
  AOI22_X1  g0526(.A1(new_n722), .A2(G329), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n332), .A2(new_n443), .A3(G190), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G311), .ZN(new_n731));
  INV_X1    g0531(.A(new_n723), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n732), .A2(G190), .A3(G200), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n727), .B1(new_n527), .B2(new_n730), .C1(new_n731), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n721), .A2(new_n715), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n719), .B(new_n735), .C1(G283), .C2(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n732), .A2(new_n443), .A3(G190), .ZN(new_n738));
  INV_X1    g0538(.A(G317), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT33), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n739), .A2(KEYINPUT33), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n724), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G322), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n737), .A2(new_n293), .A3(new_n742), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n717), .A2(new_n210), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n747), .A2(KEYINPUT94), .A3(new_n295), .ZN(new_n748));
  AOI21_X1  g0548(.A(KEYINPUT94), .B1(new_n747), .B2(new_n295), .ZN(new_n749));
  INV_X1    g0549(.A(new_n738), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n734), .A2(new_n222), .B1(new_n750), .B2(new_n268), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n736), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n216), .ZN(new_n754));
  INV_X1    g0554(.A(new_n743), .ZN(new_n755));
  INV_X1    g0555(.A(new_n725), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n225), .B1(new_n756), .B2(new_n220), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n729), .A2(G97), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n722), .A2(G159), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT32), .Z(new_n761));
  NAND4_X1  g0561(.A1(new_n752), .A2(new_n758), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n745), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n711), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n702), .A2(new_n713), .A3(new_n696), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n698), .A2(new_n765), .ZN(G396));
  NAND2_X1  g0566(.A1(new_n384), .A2(new_n642), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n394), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n458), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n459), .A2(new_n644), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n673), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n688), .A2(G330), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n773), .B(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(new_n660), .B2(new_n695), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n750), .A2(KEYINPUT96), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n750), .A2(KEYINPUT96), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G283), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n759), .B1(new_n210), .B2(new_n753), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n722), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n782), .A2(new_n731), .B1(new_n718), .B2(new_n756), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n293), .B1(new_n717), .B2(new_n216), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n785), .B1(new_n563), .B2(new_n734), .C1(new_n527), .C2(new_n755), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G159), .A2(new_n733), .B1(new_n743), .B2(G143), .ZN(new_n787));
  INV_X1    g0587(.A(G137), .ZN(new_n788));
  INV_X1    g0588(.A(G150), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n787), .B1(new_n788), .B2(new_n756), .C1(new_n789), .C2(new_n750), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT34), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n753), .A2(new_n268), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G50), .B2(new_n716), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(KEYINPUT97), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(new_n791), .B2(new_n790), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n722), .A2(G132), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n794), .A2(KEYINPUT97), .B1(G58), .B2(new_n729), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n796), .A2(new_n707), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n786), .B1(new_n792), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n711), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n711), .A2(new_n699), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n222), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n771), .A2(new_n699), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n801), .A2(new_n696), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n776), .A2(new_n805), .ZN(G384));
  INV_X1    g0606(.A(KEYINPUT40), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n417), .A2(new_n422), .ZN(new_n808));
  INV_X1    g0608(.A(new_n640), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n454), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n435), .A2(new_n436), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT37), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n814), .A2(new_n810), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n449), .B2(new_n451), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n417), .A2(new_n422), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n437), .B1(new_n818), .B2(new_n447), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n815), .B1(new_n819), .B2(new_n810), .ZN(new_n820));
  OAI21_X1  g0620(.A(KEYINPUT99), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n437), .A2(KEYINPUT37), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n450), .B1(new_n818), .B2(new_n447), .ZN(new_n823));
  INV_X1    g0623(.A(new_n451), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n810), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT99), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n814), .A2(new_n810), .A3(new_n448), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT37), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n812), .A2(new_n821), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT38), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n400), .B1(new_n408), .B2(new_n268), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n833), .A2(new_n410), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n409), .A2(new_n262), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n422), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n809), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n813), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(new_n823), .C2(new_n824), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n825), .ZN(new_n841));
  INV_X1    g0641(.A(new_n837), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n454), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n841), .A2(new_n843), .A3(KEYINPUT38), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n807), .B1(new_n832), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n376), .A2(new_n347), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(new_n369), .C1(new_n348), .C2(new_n644), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n347), .B(new_n642), .C1(new_n370), .C2(new_n376), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n771), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n685), .A2(new_n849), .A3(new_n687), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n841), .A2(new_n843), .A3(KEYINPUT38), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n841), .B2(new_n843), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n845), .A2(new_n850), .B1(new_n853), .B2(new_n807), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n688), .A2(new_n460), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n854), .B(new_n855), .Z(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(G330), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n846), .A2(new_n642), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT39), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n832), .A2(new_n859), .A3(new_n844), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT100), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT39), .B1(new_n851), .B2(new_n852), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n861), .B1(new_n860), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n438), .A2(new_n809), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n851), .A2(new_n852), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n847), .A2(new_n848), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n629), .A2(new_n644), .A3(new_n772), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(new_n770), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n866), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n857), .B(new_n872), .Z(new_n873));
  NAND2_X1  g0673(.A1(new_n674), .A2(new_n460), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n635), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n873), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n203), .B2(new_n693), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n488), .A2(new_n489), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n563), .B1(new_n879), .B2(KEYINPUT35), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n880), .B(new_n236), .C1(KEYINPUT35), .C2(new_n879), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT36), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n397), .A2(new_n398), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n883), .A2(new_n222), .A3(new_n237), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n268), .A2(G50), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT98), .ZN(new_n886));
  OAI211_X1 g0686(.A(G1), .B(new_n230), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n877), .A2(new_n882), .A3(new_n887), .ZN(G367));
  OAI21_X1  g0688(.A(new_n501), .B1(new_n619), .B2(new_n644), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n622), .A2(new_n642), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n657), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT42), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n499), .A2(new_n500), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n892), .B2(new_n538), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n644), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n615), .A2(new_n644), .ZN(new_n899));
  MUX2_X1   g0699(.A(new_n624), .B(new_n572), .S(new_n899), .Z(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT43), .Z(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT102), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n894), .A2(new_n905), .A3(new_n897), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT101), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n654), .A2(new_n892), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT103), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n660), .B(KEYINPUT41), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n657), .B1(new_n653), .B2(new_n656), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n649), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n689), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT104), .Z(new_n919));
  NAND2_X1  g0719(.A1(new_n657), .A2(new_n655), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n892), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT44), .Z(new_n922));
  NOR2_X1   g0722(.A1(new_n892), .A2(new_n920), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT45), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(new_n654), .Z(new_n926));
  OR2_X1    g0726(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n915), .B1(new_n927), .B2(new_n689), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n913), .B1(new_n911), .B2(new_n910), .C1(new_n928), .C2(new_n695), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n722), .A2(G137), .ZN(new_n930));
  AOI22_X1  g0730(.A1(G58), .A2(new_n716), .B1(new_n743), .B2(G150), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n729), .A2(G68), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n733), .A2(G50), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n930), .A2(new_n931), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(G143), .B2(new_n725), .ZN(new_n935));
  INV_X1    g0735(.A(new_n779), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(G159), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n736), .A2(G77), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n935), .A2(new_n937), .A3(new_n295), .A4(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT106), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n755), .A2(new_n718), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n779), .A2(new_n527), .B1(new_n731), .B2(new_n756), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n730), .A2(new_n216), .ZN(new_n943));
  INV_X1    g0743(.A(new_n707), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n716), .A2(G116), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT46), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n942), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n946), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT105), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n733), .A2(G283), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n722), .A2(G317), .B1(new_n736), .B2(G97), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n948), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n940), .B1(new_n941), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n711), .ZN(new_n957));
  INV_X1    g0757(.A(new_n701), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n900), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n708), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n712), .B1(new_n207), .B2(new_n553), .C1(new_n247), .C2(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n957), .A2(new_n696), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n929), .A2(new_n962), .ZN(G387));
  OAI211_X1 g0763(.A(new_n919), .B(new_n660), .C1(new_n689), .C2(new_n917), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n917), .A2(new_n695), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n944), .B1(new_n753), .B2(new_n563), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G303), .A2(new_n733), .B1(new_n743), .B2(G317), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n779), .B2(new_n731), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G322), .B2(new_n725), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT48), .Z(new_n970));
  OAI22_X1  g0770(.A1(new_n717), .A2(new_n527), .B1(new_n780), .B2(new_n730), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT109), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT49), .Z(new_n976));
  AOI211_X1 g0776(.A(new_n966), .B(new_n976), .C1(new_n722), .C2(new_n726), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n553), .A2(new_n730), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n380), .A2(new_n750), .B1(new_n734), .B2(new_n268), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n736), .A2(G97), .B1(G77), .B2(new_n716), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n980), .B(new_n707), .C1(new_n789), .C2(new_n782), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT108), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(G159), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n983), .B1(new_n982), .B2(new_n981), .C1(new_n984), .C2(new_n756), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n978), .B(new_n985), .C1(G50), .C2(new_n743), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n711), .B1(new_n977), .B2(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n653), .A2(new_n958), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n708), .B1(new_n244), .B2(new_n462), .ZN(new_n989));
  INV_X1    g0789(.A(new_n662), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n704), .A2(new_n990), .ZN(new_n991));
  AOI211_X1 g0791(.A(G45), .B(new_n990), .C1(G68), .C2(G77), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n380), .A2(G50), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT50), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n989), .A2(new_n991), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n207), .A2(G107), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n712), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n987), .A2(new_n696), .A3(new_n988), .A4(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n964), .A2(new_n965), .A3(new_n998), .ZN(G393));
  AOI22_X1  g0799(.A1(new_n936), .A2(G303), .B1(G283), .B2(new_n716), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n295), .B1(new_n722), .B2(G322), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(new_n527), .C2(new_n734), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n730), .A2(new_n563), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G311), .A2(new_n743), .B1(new_n725), .B2(G317), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT52), .ZN(new_n1005));
  NOR4_X1   g0805(.A1(new_n1002), .A2(new_n754), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT51), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n755), .A2(new_n984), .B1(new_n756), .B2(new_n789), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n936), .A2(G50), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n380), .B2(new_n734), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n717), .A2(new_n268), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n730), .A2(new_n222), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n944), .B1(new_n722), .B2(G143), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n210), .B2(new_n753), .C1(new_n1008), .C2(new_n1007), .ZN(new_n1014));
  NOR4_X1   g0814(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n711), .B1(new_n1006), .B2(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n712), .B1(new_n212), .B2(new_n207), .C1(new_n960), .C2(new_n255), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT110), .Z(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n696), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT111), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1016), .B(new_n1020), .C1(new_n891), .C2(new_n958), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n661), .B1(new_n919), .B2(new_n926), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1022), .B1(new_n927), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n926), .A2(new_n694), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(G390));
  NAND2_X1  g0826(.A1(new_n860), .A2(new_n862), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(KEYINPUT100), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n860), .A2(new_n862), .A3(new_n861), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n870), .A2(new_n858), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n685), .A2(G330), .A3(new_n687), .A4(new_n772), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(new_n868), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT112), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n858), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n832), .A2(new_n844), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n671), .B1(new_n458), .B2(new_n768), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n770), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1035), .B(new_n1036), .C1(new_n1039), .C2(new_n868), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n1031), .A2(new_n1034), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1034), .B1(new_n1031), .B2(new_n1040), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n855), .A2(G330), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n874), .A2(new_n635), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n869), .A2(new_n770), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1032), .A2(new_n868), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1046), .B1(new_n1047), .B2(new_n1033), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n771), .A2(KEYINPUT113), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n688), .A2(G330), .A3(new_n772), .A4(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1047), .A2(new_n1033), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1039), .B(new_n1050), .C1(new_n1051), .C2(new_n1049), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1045), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n661), .B1(new_n1043), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1053), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1043), .A2(new_n695), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1028), .A2(new_n699), .A3(new_n1029), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n716), .A2(G150), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1060), .B(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(G128), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(KEYINPUT54), .B(G143), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n295), .B1(new_n756), .B2(new_n1063), .C1(new_n734), .C2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G125), .B2(new_n722), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n984), .B2(new_n730), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1062), .B(new_n1067), .C1(G132), .C2(new_n743), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n220), .B2(new_n753), .C1(new_n788), .C2(new_n779), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT115), .Z(new_n1070));
  NOR2_X1   g0870(.A1(new_n779), .A2(new_n216), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n747), .B1(new_n753), .B2(new_n268), .C1(new_n527), .C2(new_n782), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1012), .B1(G116), .B2(new_n743), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n212), .B2(new_n734), .C1(new_n780), .C2(new_n756), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .A4(new_n295), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n711), .B1(new_n1070), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n802), .A2(new_n380), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1059), .A2(new_n696), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1057), .A2(new_n1058), .A3(new_n1078), .ZN(G378));
  INV_X1    g0879(.A(KEYINPUT57), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1045), .B1(new_n1043), .B2(new_n1053), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n324), .A2(new_n640), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT120), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n331), .B2(new_n336), .ZN(new_n1084));
  AOI211_X1 g0884(.A(KEYINPUT120), .B(new_n335), .C1(new_n322), .C2(new_n330), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n327), .A2(new_n311), .A3(new_n321), .A4(new_n328), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1087), .A2(KEYINPUT10), .A3(new_n315), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n314), .B1(new_n313), .B2(new_n325), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n336), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT120), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n331), .A2(new_n1083), .A3(new_n336), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1082), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1086), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1095), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n854), .A2(G330), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n853), .A2(new_n807), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n826), .B1(new_n825), .B2(new_n828), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT38), .B1(new_n1103), .B2(new_n812), .ZN(new_n1104));
  OAI211_X1 g0904(.A(KEYINPUT40), .B(new_n850), .C1(new_n1104), .C2(new_n851), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1100), .A2(new_n1105), .A3(G330), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1098), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1035), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n871), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1099), .B(new_n1108), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1098), .B1(new_n854), .B2(G330), .ZN(new_n1112));
  AND4_X1   g0912(.A1(G330), .A2(new_n1098), .A3(new_n1100), .A4(new_n1105), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n865), .B(new_n871), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1111), .A2(new_n1114), .A3(KEYINPUT121), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1108), .A2(new_n1099), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT121), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n865), .A4(new_n871), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1080), .B1(new_n1081), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1031), .A2(new_n1040), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1034), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1031), .A2(new_n1034), .A3(new_n1040), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n1053), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1045), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT122), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n872), .A2(new_n1128), .A3(new_n1099), .A4(new_n1108), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1111), .A2(new_n1114), .A3(KEYINPUT122), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1127), .A2(KEYINPUT57), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1120), .A2(new_n660), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1115), .A2(new_n695), .A3(new_n1118), .ZN(new_n1133));
  AOI211_X1 g0933(.A(G41), .B(new_n707), .C1(G77), .C2(new_n716), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT116), .Z(new_n1135));
  AOI22_X1  g0935(.A1(new_n382), .A2(new_n733), .B1(new_n738), .B2(G97), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT117), .Z(new_n1137));
  OAI221_X1 g0937(.A(new_n932), .B1(new_n756), .B2(new_n563), .C1(new_n216), .C2(new_n755), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n225), .B2(new_n753), .C1(new_n780), .C2(new_n782), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(G41), .B1(new_n707), .B2(G33), .ZN(new_n1143));
  INV_X1    g0943(.A(G132), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n750), .A2(new_n1144), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n717), .A2(new_n1064), .B1(new_n755), .B2(new_n1063), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT119), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n725), .A2(G125), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(new_n788), .C2(new_n734), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1145), .B(new_n1149), .C1(G150), .C2(new_n729), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT59), .ZN(new_n1151));
  AOI21_X1  g0951(.A(G33), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(G41), .B1(new_n722), .B2(G124), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(new_n984), .C2(new_n753), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1142), .B1(G50), .B2(new_n1143), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1156), .A2(new_n711), .B1(new_n220), .B2(new_n802), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n696), .B(new_n1157), .C1(new_n1107), .C2(new_n700), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1133), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1132), .A2(new_n1159), .ZN(G375));
  NAND2_X1  g0960(.A1(new_n868), .A2(new_n699), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n938), .B1(new_n212), .B2(new_n717), .C1(new_n779), .C2(new_n563), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n782), .A2(new_n718), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n734), .A2(new_n216), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n978), .B1(G283), .B2(new_n743), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1165), .B(new_n293), .C1(new_n527), .C2(new_n756), .ZN(new_n1166));
  NOR4_X1   g0966(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n733), .A2(G150), .B1(G50), .B2(new_n729), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n225), .B2(new_n753), .C1(new_n779), .C2(new_n1064), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n707), .B1(new_n788), .B2(new_n755), .C1(new_n782), .C2(new_n1063), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n717), .A2(new_n984), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n756), .A2(new_n1144), .ZN(new_n1172));
  NOR4_X1   g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n711), .B1(new_n1167), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1161), .A2(new_n696), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n268), .B2(new_n802), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1052), .A2(new_n1048), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1176), .B1(new_n1177), .B2(new_n695), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1052), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n914), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1178), .B1(new_n1180), .B2(new_n1053), .ZN(G381));
  NOR2_X1   g0981(.A1(G375), .A2(G378), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1183), .A2(G384), .A3(G381), .ZN(new_n1184));
  INV_X1    g0984(.A(G390), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n929), .A2(new_n962), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(G393), .A2(G396), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1184), .A2(new_n1187), .A3(new_n1188), .ZN(G407));
  OAI211_X1 g0989(.A(G407), .B(G213), .C1(G343), .C2(new_n1183), .ZN(G409));
  NAND2_X1  g0990(.A1(new_n641), .A2(G213), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1132), .A2(G378), .A3(new_n1159), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1127), .A2(new_n914), .A3(new_n1118), .A4(new_n1115), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1130), .A2(new_n695), .A3(new_n1129), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1158), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1058), .A2(new_n1078), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1056), .B2(new_n1054), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1192), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT60), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1179), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1179), .A2(new_n1201), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1202), .A2(new_n660), .A3(new_n1055), .A4(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1204), .A2(G384), .A3(new_n1178), .ZN(new_n1205));
  AOI21_X1  g1005(.A(G384), .B1(new_n1204), .B2(new_n1178), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1200), .A2(KEYINPUT62), .A3(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT126), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1193), .A2(KEYINPUT123), .A3(new_n1199), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT123), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT124), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n1191), .A4(new_n1207), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1193), .A2(new_n1199), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT123), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1193), .A2(KEYINPUT123), .A3(new_n1199), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1217), .A2(new_n1191), .A3(new_n1207), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(KEYINPUT124), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1214), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT62), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1209), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT61), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1207), .A2(G2897), .A3(new_n1192), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1207), .B1(G2897), .B2(new_n1192), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1224), .B1(new_n1227), .B2(new_n1200), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT125), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT127), .B1(new_n1223), .B2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(G393), .B(G396), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1185), .B1(new_n929), .B2(new_n962), .ZN(new_n1234));
  OR3_X1    g1034(.A1(new_n1187), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1187), .B2(new_n1234), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT127), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT62), .B1(new_n1214), .B2(new_n1220), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1229), .B(new_n1238), .C1(new_n1239), .C2(new_n1209), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1231), .A2(new_n1237), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT63), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1237), .B1(new_n1242), .B2(new_n1221), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1200), .A2(KEYINPUT63), .A3(new_n1207), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1212), .A2(new_n1191), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1226), .B2(new_n1225), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1224), .A3(new_n1244), .A4(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1241), .A2(new_n1247), .ZN(G405));
  NAND2_X1  g1048(.A1(G375), .A2(new_n1198), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1193), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(new_n1207), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1237), .B(new_n1251), .ZN(G402));
endmodule


