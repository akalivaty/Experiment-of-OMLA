//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n630, new_n632, new_n633,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT64), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OAI22_X1  g037(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n456), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n463), .B1(new_n461), .B2(new_n460), .ZN(new_n464));
  XOR2_X1   g039(.A(new_n464), .B(KEYINPUT66), .Z(G319));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT67), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT68), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n472), .A3(G2104), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n470), .A2(new_n471), .A3(new_n474), .A4(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n479), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n480));
  OAI22_X1  g055(.A1(new_n477), .A2(new_n478), .B1(new_n480), .B2(new_n471), .ZN(new_n481));
  INV_X1    g056(.A(G101), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT67), .B(G2104), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT69), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n467), .A2(new_n469), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n485), .A2(new_n486), .A3(new_n471), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n482), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n481), .A2(new_n488), .ZN(G160));
  INV_X1    g064(.A(new_n477), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT70), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G112), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n474), .A2(new_n476), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(G2105), .A3(new_n470), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n498), .B2(G124), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G162));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n470), .A2(new_n474), .A3(new_n476), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(G102), .A2(G2104), .ZN(new_n506));
  AOI21_X1  g081(.A(G2105), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n470), .A2(G126), .A3(new_n474), .A4(new_n476), .ZN(new_n508));
  NAND2_X1  g083(.A1(G114), .A2(G2104), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n471), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n503), .A2(G2105), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT4), .B1(new_n479), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g087(.A1(new_n507), .A2(new_n510), .A3(new_n512), .ZN(G164));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(G88), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(G50), .A3(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  OAI21_X1  g101(.A(G62), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n514), .B1(new_n523), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G62), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n517), .B2(new_n518), .ZN(new_n533));
  INV_X1    g108(.A(new_n528), .ZN(new_n534));
  OAI21_X1  g109(.A(G651), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n535), .A2(KEYINPUT71), .A3(new_n521), .A4(new_n522), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n531), .A2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  XOR2_X1   g114(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G63), .A2(G651), .ZN(new_n543));
  AND2_X1   g118(.A1(KEYINPUT6), .A2(G651), .ZN(new_n544));
  NOR2_X1   g119(.A1(KEYINPUT6), .A2(G651), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT73), .B(G89), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(new_n519), .ZN(new_n549));
  OR2_X1    g124(.A1(KEYINPUT6), .A2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(KEYINPUT6), .A2(G651), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n516), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G51), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n542), .A2(new_n549), .A3(new_n553), .ZN(G286));
  INV_X1    g129(.A(G286), .ZN(G168));
  AOI22_X1  g130(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n524), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n520), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G52), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n526), .A2(new_n525), .B1(new_n544), .B2(new_n545), .ZN(new_n560));
  INV_X1    g135(.A(G90), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n558), .A2(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n557), .A2(new_n562), .ZN(G171));
  AOI22_X1  g138(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n524), .ZN(new_n565));
  INV_X1    g140(.A(G43), .ZN(new_n566));
  INV_X1    g141(.A(G81), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n558), .A2(new_n566), .B1(new_n560), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  NOR2_X1   g149(.A1(new_n525), .A2(new_n526), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n546), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n576), .A2(KEYINPUT74), .A3(G91), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n578));
  INV_X1    g153(.A(G91), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n560), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G53), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT9), .B1(new_n558), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT9), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n552), .A2(new_n583), .A3(G53), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n577), .A2(new_n580), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G65), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n519), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n575), .A2(KEYINPUT75), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G78), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n585), .A2(new_n593), .ZN(G299));
  INV_X1    g169(.A(G171), .ZN(G301));
  NAND3_X1  g170(.A1(new_n519), .A2(new_n520), .A3(G87), .ZN(new_n596));
  INV_X1    g171(.A(G74), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n517), .A2(new_n597), .A3(new_n518), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n520), .A2(G49), .A3(G543), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(G288));
  AOI22_X1  g176(.A1(new_n576), .A2(G86), .B1(G48), .B2(new_n552), .ZN(new_n602));
  OAI21_X1  g177(.A(G61), .B1(new_n525), .B2(new_n526), .ZN(new_n603));
  NAND2_X1  g178(.A1(G73), .A2(G543), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n524), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(G305));
  NAND2_X1  g182(.A1(new_n552), .A2(G47), .ZN(new_n608));
  INV_X1    g183(.A(G85), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n560), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(new_n524), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n552), .A2(G54), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n576), .A2(KEYINPUT10), .A3(G92), .ZN(new_n617));
  AOI21_X1  g192(.A(KEYINPUT10), .B1(new_n576), .B2(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n519), .A2(new_n587), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n575), .A2(KEYINPUT75), .ZN(new_n621));
  OAI21_X1  g196(.A(G66), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(G79), .A2(G543), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n524), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n615), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n615), .B1(new_n625), .B2(G868), .ZN(G321));
  MUX2_X1   g202(.A(G299), .B(G286), .S(G868), .Z(G297));
  XNOR2_X1  g203(.A(G297), .B(KEYINPUT76), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n625), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n625), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g209(.A(KEYINPUT77), .B(KEYINPUT11), .ZN(new_n635));
  XNOR2_X1  g210(.A(G323), .B(new_n635), .ZN(G282));
  NAND2_X1  g211(.A1(new_n490), .A2(G135), .ZN(new_n637));
  INV_X1    g212(.A(G123), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n471), .A2(G111), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  OAI221_X1 g215(.A(new_n637), .B1(new_n497), .B2(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT79), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n484), .A2(new_n487), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(new_n479), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT12), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT78), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n646), .A2(new_n647), .A3(new_n653), .ZN(G156));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n660), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G14), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(G401));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT80), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT18), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n673), .B(KEYINPUT17), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n678), .B(new_n675), .C1(new_n672), .C2(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n679), .A2(new_n672), .A3(new_n674), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G2096), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT81), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT82), .ZN(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  AOI21_X1  g267(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n696), .A2(KEYINPUT20), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(KEYINPUT20), .ZN(new_n698));
  OAI221_X1 g273(.A(new_n695), .B1(new_n688), .B2(new_n694), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n703), .B1(new_n701), .B2(new_n702), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n686), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(new_n686), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n708), .A2(new_n709), .A3(new_n704), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  AND3_X1   g286(.A1(new_n707), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n711), .B1(new_n707), .B2(new_n710), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(G229));
  XOR2_X1   g289(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n715));
  AOI21_X1  g290(.A(G29), .B1(new_n715), .B2(G34), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G34), .B2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT93), .ZN(new_n718));
  INV_X1    g293(.A(G160), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G2084), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G5), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G171), .B2(new_n724), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT26), .Z(new_n728));
  INV_X1    g303(.A(G129), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n497), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G105), .B2(new_n648), .ZN(new_n731));
  INV_X1    g306(.A(G141), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n477), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT94), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(new_n720), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n720), .B2(G32), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n723), .B1(G1961), .B2(new_n726), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT97), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(new_n739), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT85), .B(G16), .Z(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(G19), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n569), .B2(new_n744), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT89), .B(G1341), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G29), .A2(G33), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT90), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n490), .A2(G139), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(new_n471), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n754));
  NAND3_X1  g329(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n751), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n750), .B1(new_n757), .B2(new_n720), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n748), .B1(new_n442), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n442), .B2(new_n758), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n724), .A2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G168), .B2(new_n724), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1966), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n721), .A2(new_n722), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n726), .A2(G1961), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G11), .ZN(new_n767));
  INV_X1    g342(.A(G28), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n768), .B2(KEYINPUT30), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(KEYINPUT30), .B2(new_n768), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n765), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n763), .A2(new_n764), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n643), .A2(G29), .A3(new_n644), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n742), .A2(new_n760), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n743), .A2(G20), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT99), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT23), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G16), .B2(G299), .ZN(new_n779));
  INV_X1    g354(.A(G1956), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n720), .A2(G26), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT28), .ZN(new_n783));
  INV_X1    g358(.A(G128), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n471), .A2(G116), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n786));
  OAI22_X1  g361(.A1(new_n497), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G140), .B2(new_n490), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n783), .B1(new_n788), .B2(new_n720), .ZN(new_n789));
  INV_X1    g364(.A(G2067), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(KEYINPUT96), .B2(new_n773), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n775), .A2(new_n781), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G4), .A2(G16), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n625), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT88), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1348), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n720), .A2(G35), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G162), .B2(new_n720), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT29), .Z(new_n800));
  INV_X1    g375(.A(G2090), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n741), .A2(new_n793), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n720), .A2(G27), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G164), .B2(new_n720), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G2078), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT98), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G6), .A2(G16), .ZN(new_n811));
  INV_X1    g386(.A(G48), .ZN(new_n812));
  INV_X1    g387(.A(G86), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n558), .A2(new_n812), .B1(new_n560), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(new_n605), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n811), .B1(new_n815), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT32), .ZN(new_n817));
  INV_X1    g392(.A(G1981), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n743), .A2(G22), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G166), .B2(new_n743), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G1971), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(G1971), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n724), .A2(G23), .ZN(new_n824));
  INV_X1    g399(.A(G288), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(new_n724), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT33), .B(G1976), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT86), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n826), .B(new_n828), .Z(new_n829));
  NAND4_X1  g404(.A1(new_n819), .A2(new_n822), .A3(new_n823), .A4(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT87), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT34), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n832), .A2(KEYINPUT34), .A3(new_n833), .ZN(new_n837));
  NOR2_X1   g412(.A1(G25), .A2(G29), .ZN(new_n838));
  OR2_X1    g413(.A1(G95), .A2(G2105), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n839), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n840));
  INV_X1    g415(.A(G131), .ZN(new_n841));
  INV_X1    g416(.A(G119), .ZN(new_n842));
  OAI221_X1 g417(.A(new_n840), .B1(new_n841), .B2(new_n477), .C1(new_n497), .C2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT84), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n838), .B1(new_n848), .B2(G29), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G1991), .Z(new_n850));
  XOR2_X1   g425(.A(new_n849), .B(new_n850), .Z(new_n851));
  NOR2_X1   g426(.A1(new_n744), .A2(G24), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n613), .B2(new_n744), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G1986), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n836), .A2(new_n837), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT36), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT36), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n836), .A2(new_n858), .A3(new_n837), .A4(new_n855), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n810), .B1(new_n857), .B2(new_n859), .ZN(G311));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n859), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n861), .A2(new_n809), .A3(new_n803), .ZN(G150));
  NAND2_X1  g437(.A1(new_n625), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n576), .A2(G93), .B1(G55), .B2(new_n552), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n524), .B2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n569), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n864), .B(new_n868), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n870), .A2(new_n871), .A3(G860), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(G860), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n874));
  XOR2_X1   g449(.A(new_n873), .B(new_n874), .Z(new_n875));
  OR2_X1    g450(.A1(new_n872), .A2(new_n875), .ZN(G145));
  NAND2_X1  g451(.A1(new_n490), .A2(G142), .ZN(new_n877));
  INV_X1    g452(.A(G130), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n471), .A2(KEYINPUT101), .A3(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT101), .B1(new_n471), .B2(G118), .ZN(new_n880));
  OR2_X1    g455(.A1(G106), .A2(G2105), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(G2104), .A3(new_n881), .ZN(new_n882));
  OAI221_X1 g457(.A(new_n877), .B1(new_n497), .B2(new_n878), .C1(new_n879), .C2(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n650), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n650), .A2(new_n883), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n847), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n847), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n505), .A2(new_n506), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n471), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n508), .A2(new_n509), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(G2105), .ZN(new_n892));
  INV_X1    g467(.A(new_n512), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n788), .B(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n757), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n731), .A2(new_n734), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n896), .B1(new_n731), .B2(new_n734), .ZN(new_n899));
  XNOR2_X1  g474(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n735), .A2(new_n757), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(new_n897), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n895), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n900), .B1(new_n898), .B2(new_n899), .ZN(new_n906));
  INV_X1    g481(.A(new_n895), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(new_n897), .A3(new_n902), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n888), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n905), .A2(new_n888), .A3(new_n909), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n645), .B(new_n719), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n911), .A2(KEYINPUT104), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n913), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(KEYINPUT104), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n915), .B1(new_n916), .B2(new_n910), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(G162), .ZN(new_n919));
  INV_X1    g494(.A(G37), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n917), .A3(new_n500), .ZN(new_n921));
  AND4_X1   g496(.A1(KEYINPUT40), .A2(new_n919), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G37), .B1(new_n918), .B2(G162), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT40), .B1(new_n923), .B2(new_n921), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n922), .A2(new_n924), .ZN(G395));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n611), .A2(new_n524), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n576), .A2(G85), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .A4(new_n608), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT106), .B1(new_n610), .B2(new_n612), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n930), .A2(new_n825), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n825), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(G305), .A2(new_n536), .A3(new_n530), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(G305), .B1(new_n536), .B2(new_n530), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n926), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  OAI221_X1 g514(.A(KEYINPUT107), .B1(new_n936), .B2(new_n937), .C1(new_n932), .C2(new_n933), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n930), .A2(new_n931), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(G288), .ZN(new_n943));
  INV_X1    g518(.A(new_n937), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n930), .A2(new_n825), .A3(new_n931), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n935), .A4(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n934), .A2(new_n938), .A3(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n941), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n941), .A2(new_n950), .A3(KEYINPUT109), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n625), .A2(G299), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n593), .B(new_n585), .C1(new_n619), .C2(new_n624), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n625), .A2(KEYINPUT105), .A3(G299), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(KEYINPUT41), .A3(new_n961), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT41), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n957), .A2(new_n964), .A3(new_n959), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n868), .B(new_n632), .ZN(new_n967));
  MUX2_X1   g542(.A(new_n962), .B(new_n966), .S(new_n967), .Z(new_n968));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n951), .A2(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n956), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n968), .B1(new_n956), .B2(new_n970), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  MUX2_X1   g548(.A(new_n867), .B(new_n973), .S(G868), .Z(G295));
  MUX2_X1   g549(.A(new_n867), .B(new_n973), .S(G868), .Z(G331));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  AND3_X1   g551(.A1(G286), .A2(KEYINPUT111), .A3(G171), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT111), .B1(G286), .B2(G171), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n868), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(G168), .B2(G301), .ZN(new_n982));
  NOR3_X1   g557(.A1(G286), .A2(G171), .A3(KEYINPUT110), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n979), .B(new_n980), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  OAI22_X1  g559(.A1(new_n982), .A2(new_n983), .B1(new_n977), .B2(new_n978), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n868), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT41), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n962), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n957), .A2(new_n959), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(KEYINPUT41), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n954), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT109), .B1(new_n941), .B2(new_n950), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n989), .B(new_n991), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n987), .A2(new_n966), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n984), .A2(new_n986), .A3(new_n962), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(new_n953), .A3(new_n954), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n994), .A2(new_n920), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n994), .A2(new_n998), .A3(KEYINPUT112), .A4(new_n920), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n976), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n998), .A2(new_n920), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n955), .A2(new_n996), .A3(new_n995), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT43), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT44), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n976), .A3(new_n994), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n976), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(G397));
  XOR2_X1   g588(.A(new_n847), .B(new_n850), .Z(new_n1014));
  XNOR2_X1  g589(.A(new_n788), .B(G2067), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n736), .A2(G1996), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n735), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1015), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(G290), .A2(G1986), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G290), .A2(G1986), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT45), .B1(new_n894), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G40), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n481), .A2(new_n1026), .A3(new_n488), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1023), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT124), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n894), .A2(new_n1027), .A3(new_n1024), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n1033));
  INV_X1    g608(.A(G1976), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G288), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g612(.A(KEYINPUT114), .B(KEYINPUT52), .C1(G288), .C2(new_n1034), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n825), .A2(G1976), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1032), .A2(new_n1039), .A3(G8), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n818), .ZN(new_n1042));
  OAI21_X1  g617(.A(G1981), .B1(new_n814), .B2(new_n605), .ZN(new_n1043));
  NOR2_X1   g618(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n818), .B1(new_n602), .B2(new_n606), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n814), .A2(G1981), .A3(new_n605), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1032), .A2(G8), .A3(new_n1046), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1041), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n512), .B1(new_n891), .B2(G2105), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1384), .B1(new_n1053), .B2(new_n890), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1054), .B2(new_n1027), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1036), .B1(new_n1055), .B2(new_n1040), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT117), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1032), .A2(G8), .A3(new_n1040), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT52), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1041), .A4(new_n1050), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1057), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n530), .A2(G8), .A3(new_n536), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT55), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT113), .B(G1971), .Z(new_n1065));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(G1384), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1027), .B1(G164), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1065), .B1(new_n1069), .B2(new_n1025), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n648), .A2(G101), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n496), .A2(G137), .A3(new_n471), .A4(new_n470), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n479), .A2(G125), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G113), .A2(G2104), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G2105), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1072), .A2(G40), .A3(new_n1073), .A4(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n894), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1071), .A2(new_n1080), .A3(new_n801), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1052), .B(new_n1064), .C1(new_n1070), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1070), .A2(new_n1081), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(G8), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1064), .ZN(new_n1086));
  AND4_X1   g661(.A1(new_n1031), .A2(new_n1062), .A3(new_n1083), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1064), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1084), .B2(G8), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(new_n1082), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1031), .B1(new_n1090), .B2(new_n1062), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT122), .B(KEYINPUT51), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1066), .B1(G164), .B2(G1384), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1078), .B1(new_n894), .B2(new_n1067), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1966), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1071), .A2(new_n1080), .A3(new_n722), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(G168), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1093), .B1(new_n1100), .B2(G8), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1079), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1027), .B1(G164), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n894), .B2(new_n1024), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1106), .A2(new_n722), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1052), .B1(new_n1107), .B2(G168), .ZN(new_n1108));
  OAI22_X1  g683(.A1(new_n1107), .A2(G168), .B1(KEYINPUT122), .B2(KEYINPUT51), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1101), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT125), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT119), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1113));
  INV_X1    g688(.A(G1961), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1071), .A2(new_n1080), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1096), .B2(G2078), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1094), .A2(new_n1095), .A3(KEYINPUT53), .A4(new_n443), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(G171), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1109), .A2(new_n1108), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1125), .B(KEYINPUT62), .C1(new_n1126), .C2(new_n1101), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1092), .A2(new_n1112), .A3(new_n1124), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1117), .A2(KEYINPUT123), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1113), .A2(new_n1130), .A3(new_n1116), .A4(new_n1114), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(G171), .B1(new_n1132), .B2(new_n1122), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1134), .B1(new_n1135), .B2(G301), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1110), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g712(.A(G171), .B(new_n1122), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1123), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1134), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(new_n1092), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n780), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G299), .B(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT56), .B(G2072), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1094), .A2(new_n1095), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1142), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n625), .ZN(new_n1148));
  INV_X1    g723(.A(G1348), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1113), .A2(new_n1149), .A3(new_n1116), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1054), .A2(new_n790), .A3(new_n1027), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1148), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1144), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1094), .A2(new_n1095), .A3(new_n1145), .ZN(new_n1154));
  AOI21_X1  g729(.A(G1956), .B1(new_n1071), .B2(new_n1080), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1147), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(KEYINPUT120), .B(new_n1147), .C1(new_n1152), .C2(new_n1157), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1156), .A2(new_n1147), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1094), .A2(new_n1095), .A3(new_n1017), .ZN(new_n1165));
  XOR2_X1   g740(.A(KEYINPUT58), .B(G1341), .Z(new_n1166));
  NAND2_X1  g741(.A1(new_n1032), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n569), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT59), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(new_n1171), .A3(new_n569), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1163), .A2(new_n1164), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1150), .A2(KEYINPUT60), .A3(new_n1151), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1176), .A2(new_n625), .A3(new_n1177), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1156), .A2(KEYINPUT61), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1147), .A2(KEYINPUT121), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1142), .A2(new_n1144), .A3(new_n1146), .A4(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1177), .A2(new_n625), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1173), .A2(new_n1178), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1162), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1128), .B1(new_n1141), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1050), .A2(new_n1034), .A3(new_n825), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1048), .B(KEYINPUT116), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1055), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1059), .A2(new_n1041), .A3(new_n1050), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1192), .B1(new_n1083), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(G168), .A2(G8), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1107), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1090), .A2(new_n1062), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT63), .ZN(new_n1199));
  AND2_X1   g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NOR4_X1   g775(.A1(new_n1193), .A2(new_n1107), .A3(new_n1199), .A4(new_n1196), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1201), .A2(new_n1090), .ZN(new_n1202));
  OAI211_X1 g777(.A(KEYINPUT118), .B(new_n1195), .C1(new_n1200), .C2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT118), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n1198), .A2(new_n1199), .B1(new_n1090), .B2(new_n1201), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1204), .B1(new_n1205), .B2(new_n1194), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1030), .B1(new_n1188), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1028), .B1(new_n1015), .B2(new_n736), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT46), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1029), .A2(new_n1017), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1212), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1213));
  XOR2_X1   g788(.A(new_n1213), .B(KEYINPUT47), .Z(new_n1214));
  NOR2_X1   g789(.A1(new_n1028), .A2(new_n1021), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT127), .ZN(new_n1216));
  XOR2_X1   g791(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1217));
  OAI22_X1  g792(.A1(new_n1020), .A2(new_n1028), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AND2_X1   g793(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n848), .A2(new_n850), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n1019), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1221), .B1(new_n790), .B2(new_n788), .ZN(new_n1222));
  OAI22_X1  g797(.A1(new_n1218), .A2(new_n1219), .B1(new_n1222), .B2(new_n1028), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n1214), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1208), .A2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g800(.A(new_n464), .B1(new_n668), .B2(new_n669), .ZN(new_n1227));
  NOR2_X1   g801(.A1(G227), .A2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g802(.A(new_n1228), .B1(new_n712), .B2(new_n713), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1230));
  NAND2_X1  g804(.A1(new_n1230), .A2(KEYINPUT43), .ZN(new_n1231));
  AOI21_X1  g805(.A(new_n1229), .B1(new_n1231), .B2(new_n1009), .ZN(new_n1232));
  NAND2_X1  g806(.A1(new_n923), .A2(new_n921), .ZN(new_n1233));
  AND2_X1   g807(.A1(new_n1232), .A2(new_n1233), .ZN(G308));
  NAND2_X1  g808(.A1(new_n1232), .A2(new_n1233), .ZN(G225));
endmodule


