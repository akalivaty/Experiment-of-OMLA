//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971;
  INV_X1    g000(.A(G127gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT74), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT74), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G127gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n205), .A3(G134gat), .ZN(new_n206));
  OR3_X1    g005(.A1(new_n202), .A2(KEYINPUT73), .A3(G134gat), .ZN(new_n207));
  INV_X1    g006(.A(G134gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G127gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT73), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212));
  INV_X1    g011(.A(G113gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G120gat), .ZN(new_n214));
  INV_X1    g013(.A(G120gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G113gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT75), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(new_n213), .B2(G120gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n215), .A2(KEYINPUT75), .A3(G113gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n219), .B(new_n220), .C1(G113gat), .C2(new_n215), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n202), .A2(G134gat), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n209), .A2(new_n222), .A3(new_n212), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n211), .A2(new_n217), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT27), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT27), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G183gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n227), .A2(new_n229), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT28), .ZN(new_n236));
  AND2_X1   g035(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT27), .B(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT69), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n235), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT70), .B1(new_n229), .B2(new_n231), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(KEYINPUT70), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n237), .A2(new_n238), .A3(new_n236), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n242), .A2(KEYINPUT71), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT71), .B1(new_n242), .B2(new_n247), .ZN(new_n249));
  NOR2_X1   g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT26), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT26), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(KEYINPUT72), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n256));
  AND3_X1   g055(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n253), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n248), .A2(new_n249), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G169gat), .ZN(new_n262));
  INV_X1    g061(.A(G176gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT23), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n257), .B2(new_n256), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(new_n250), .B2(KEYINPUT23), .ZN(new_n268));
  NAND3_X1  g067(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(G183gat), .B2(G190gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT24), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT64), .B1(new_n259), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n259), .A2(KEYINPUT64), .A3(new_n271), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n268), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n267), .A2(KEYINPUT66), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n266), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n227), .A2(new_n228), .A3(new_n232), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n271), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n269), .A2(KEYINPUT67), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n281), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n278), .A2(new_n279), .A3(new_n280), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n250), .A2(KEYINPUT23), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT25), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n277), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n224), .B1(new_n261), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G227gat), .ZN(new_n290));
  INV_X1    g089(.A(G233gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n277), .A2(new_n287), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n211), .A2(new_n217), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n221), .A2(new_n223), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n260), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT28), .B1(new_n233), .B2(new_n234), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT70), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(new_n243), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n241), .A2(new_n298), .B1(new_n300), .B2(new_n246), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n297), .B1(new_n301), .B2(KEYINPUT71), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n293), .B(new_n296), .C1(new_n302), .C2(new_n248), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n289), .A2(new_n292), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n289), .A2(KEYINPUT76), .A3(new_n303), .A4(new_n292), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT33), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n292), .B1(new_n289), .B2(new_n303), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT34), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G71gat), .B(G99gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT77), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(G15gat), .ZN(new_n316));
  INV_X1    g115(.A(G43gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n310), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n311), .B(KEYINPUT34), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT33), .B1(new_n306), .B2(new_n307), .ZN(new_n321));
  INV_X1    g120(.A(new_n318), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n308), .A2(KEYINPUT32), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(G8gat), .B(G36gat), .Z(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT80), .ZN(new_n328));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n328), .B(new_n329), .Z(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT78), .B(G197gat), .ZN(new_n331));
  INV_X1    g130(.A(G204gat), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n331), .A2(new_n332), .ZN(new_n334));
  INV_X1    g133(.A(G211gat), .ZN(new_n335));
  INV_X1    g134(.A(G218gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI22_X1  g136(.A1(new_n333), .A2(new_n334), .B1(KEYINPUT22), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G211gat), .B(G218gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n342));
  NAND2_X1  g141(.A1(G226gat), .A2(G233gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n293), .B1(new_n302), .B2(new_n248), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n242), .A2(new_n247), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT71), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n260), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n301), .A2(KEYINPUT71), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n288), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(new_n343), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n342), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n343), .B1(new_n352), .B2(KEYINPUT29), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT79), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n341), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n347), .A2(new_n353), .A3(new_n340), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n330), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n345), .A2(new_n344), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT79), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n342), .B1(new_n362), .B2(new_n343), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n340), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n358), .ZN(new_n365));
  INV_X1    g164(.A(new_n330), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n359), .A2(KEYINPUT30), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n364), .A2(new_n369), .A3(new_n365), .A4(new_n366), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n340), .B2(KEYINPUT29), .ZN(new_n374));
  INV_X1    g173(.A(G141gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G148gat), .ZN(new_n376));
  INV_X1    g175(.A(G148gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G141gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n376), .A2(new_n378), .B1(KEYINPUT2), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(KEYINPUT81), .A3(new_n379), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT81), .ZN(new_n384));
  INV_X1    g183(.A(new_n379), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(new_n381), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n380), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n382), .A2(new_n379), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n379), .A2(KEYINPUT2), .ZN(new_n389));
  XNOR2_X1  g188(.A(G141gat), .B(G148gat), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n388), .B(new_n384), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n372), .B1(new_n394), .B2(KEYINPUT84), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n373), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT82), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n398), .A3(new_n373), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n346), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n340), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n395), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G22gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n405), .A2(KEYINPUT85), .ZN(new_n406));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT31), .B(G50gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  MUX2_X1   g208(.A(new_n405), .B(new_n406), .S(new_n409), .Z(new_n410));
  XNOR2_X1  g209(.A(new_n404), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n325), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n319), .A2(new_n323), .A3(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n326), .A2(new_n371), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n224), .A2(new_n392), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT83), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n224), .B2(new_n392), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(KEYINPUT83), .A3(new_n416), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n296), .B1(new_n373), .B2(new_n392), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n420), .A2(new_n421), .B1(new_n400), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT5), .ZN(new_n425));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n296), .B(new_n392), .ZN(new_n428));
  INV_X1    g227(.A(new_n416), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n426), .B1(new_n429), .B2(new_n418), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n422), .B1(new_n397), .B2(new_n399), .ZN(new_n431));
  OAI221_X1 g230(.A(KEYINPUT5), .B1(new_n426), .B2(new_n428), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G1gat), .B(G29gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT0), .ZN(new_n434));
  XOR2_X1   g233(.A(G57gat), .B(G85gat), .Z(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n427), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n427), .B2(new_n432), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT6), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n440));
  AOI211_X1 g239(.A(new_n440), .B(new_n436), .C1(new_n427), .C2(new_n432), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n414), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n326), .A2(new_n444), .A3(new_n411), .A4(new_n413), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT35), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n446), .B(new_n445), .C1(new_n414), .C2(new_n442), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n442), .B1(new_n368), .B2(new_n370), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(new_n411), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT36), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n319), .A2(new_n323), .A3(new_n412), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n412), .B1(new_n319), .B2(new_n323), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n326), .A2(KEYINPUT36), .A3(new_n413), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT39), .ZN(new_n458));
  INV_X1    g257(.A(new_n426), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n420), .A2(new_n421), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n458), .B(new_n459), .C1(new_n460), .C2(new_n431), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n458), .B1(new_n428), .B2(new_n426), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(new_n424), .B2(new_n426), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n463), .A3(new_n436), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT40), .B1(new_n464), .B2(KEYINPUT86), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n461), .A2(new_n463), .A3(new_n466), .A4(new_n436), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n438), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT40), .A4(new_n436), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT87), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n368), .A2(new_n468), .A3(new_n370), .A4(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n364), .A2(new_n473), .A3(new_n365), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n474), .A2(new_n330), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT38), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n364), .A2(new_n365), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(KEYINPUT37), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n341), .B1(new_n361), .B2(new_n363), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n347), .A2(new_n353), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n473), .B1(new_n480), .B2(new_n340), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n474), .A2(new_n330), .A3(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n475), .A2(new_n478), .B1(new_n483), .B2(new_n476), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n442), .A2(new_n367), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n411), .B(new_n472), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n457), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n448), .B(new_n449), .C1(new_n451), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G229gat), .A2(G233gat), .ZN(new_n489));
  INV_X1    g288(.A(G1gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT16), .ZN(new_n491));
  INV_X1    g290(.A(G15gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G22gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n405), .A2(G15gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(G1gat), .B1(new_n493), .B2(new_n494), .ZN(new_n497));
  OAI21_X1  g296(.A(G8gat), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n497), .ZN(new_n499));
  INV_X1    g298(.A(G8gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n317), .A2(G50gat), .ZN(new_n503));
  INV_X1    g302(.A(G50gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G43gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n505), .A3(KEYINPUT15), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT90), .B(KEYINPUT15), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT91), .B1(new_n504), .B2(G43gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n504), .A2(G43gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n504), .A2(KEYINPUT91), .A3(G43gat), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G29gat), .ZN(new_n513));
  INV_X1    g312(.A(G36gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT89), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT89), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n517), .A3(KEYINPUT14), .ZN(new_n518));
  NAND2_X1  g317(.A1(G29gat), .A2(G36gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n516), .B(new_n520), .C1(G29gat), .C2(G36gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n506), .B1(new_n512), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n515), .A2(new_n517), .A3(KEYINPUT14), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n519), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n506), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n502), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n523), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n498), .A2(new_n501), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n530), .B1(new_n523), .B2(new_n528), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n489), .B(new_n529), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n317), .B2(G50gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(new_n503), .A3(new_n511), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT90), .B(KEYINPUT15), .Z(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n527), .B1(new_n526), .B2(new_n542), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n524), .A2(new_n506), .A3(new_n525), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n532), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n529), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n489), .B(KEYINPUT13), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT17), .B1(new_n543), .B2(new_n544), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n532), .A3(new_n531), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n489), .A4(new_n529), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n537), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G197gat), .ZN(new_n554));
  XOR2_X1   g353(.A(KEYINPUT11), .B(G169gat), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT12), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n537), .A2(new_n551), .A3(new_n557), .A4(new_n548), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n488), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G71gat), .B(G78gat), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(G57gat), .A2(G64gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(G57gat), .A2(G64gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n563), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n569), .A3(new_n563), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(new_n202), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n572), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n502), .B1(new_n578), .B2(KEYINPUT21), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n579), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n582));
  INV_X1    g381(.A(G155gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  AND3_X1   g385(.A1(new_n580), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n586), .B1(new_n580), .B2(new_n581), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT41), .ZN(new_n590));
  INV_X1    g389(.A(G232gat), .ZN(new_n591));
  NOR3_X1   g390(.A1(new_n590), .A2(new_n591), .A3(new_n291), .ZN(new_n592));
  INV_X1    g391(.A(new_n525), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n542), .A2(new_n518), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n544), .B1(new_n506), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G99gat), .B(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT8), .ZN(new_n599));
  OR2_X1    g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  OR2_X1    g399(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n601));
  AND2_X1   g400(.A1(G85gat), .A2(G92gat), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n599), .B(new_n600), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(G85gat), .A2(G92gat), .ZN(new_n607));
  NOR3_X1   g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n597), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(G85gat), .A2(G92gat), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n610), .B1(new_n607), .B2(new_n606), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n601), .A2(new_n604), .A3(new_n602), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n611), .A2(new_n612), .A3(new_n596), .A4(new_n599), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n592), .B1(new_n595), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n531), .A2(new_n614), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n616), .B1(new_n617), .B2(new_n534), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n616), .B(new_n621), .C1(new_n617), .C2(new_n534), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT94), .B(G134gat), .ZN(new_n623));
  INV_X1    g422(.A(G162gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n590), .B1(new_n591), .B2(new_n291), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  AND4_X1   g426(.A1(KEYINPUT96), .A2(new_n620), .A3(new_n622), .A4(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n630), .A2(new_n627), .B1(new_n620), .B2(new_n622), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n589), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n614), .A2(new_n571), .A3(new_n572), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n568), .A2(new_n569), .A3(new_n563), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n613), .B(new_n609), .C1(new_n637), .C2(new_n570), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n615), .A2(new_n578), .A3(KEYINPUT10), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n635), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(new_n638), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(new_n635), .ZN(new_n644));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT97), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n562), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n442), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT98), .B(G1gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1324gat));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660));
  INV_X1    g459(.A(new_n371), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n488), .A2(new_n661), .A3(new_n561), .A4(new_n654), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n500), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n660), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT100), .Z(new_n666));
  NOR3_X1   g465(.A1(new_n662), .A2(new_n660), .A3(new_n664), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n662), .A2(G8gat), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT101), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(KEYINPUT101), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n671), .ZN(G1325gat));
  NOR3_X1   g471(.A1(new_n655), .A2(new_n492), .A3(new_n457), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n453), .A2(new_n454), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n492), .B1(new_n655), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n678), .B(new_n492), .C1(new_n655), .C2(new_n675), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n673), .B1(new_n677), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n655), .A2(new_n411), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n371), .A2(new_n656), .ZN(new_n684));
  INV_X1    g483(.A(new_n411), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(KEYINPUT105), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n450), .B2(new_n411), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n457), .A2(new_n486), .A3(new_n686), .A4(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n448), .A3(new_n449), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n632), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n488), .A2(KEYINPUT44), .A3(new_n632), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n589), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n559), .A2(KEYINPUT104), .A3(new_n560), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT104), .B1(new_n559), .B2(new_n560), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n696), .A2(new_n700), .A3(new_n651), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G29gat), .B1(new_n702), .B2(new_n656), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n628), .A2(new_n631), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n696), .A2(new_n704), .A3(new_n651), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n562), .A2(new_n513), .A3(new_n442), .A4(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n703), .A2(new_n708), .ZN(G1328gat));
  OAI21_X1  g508(.A(G36gat), .B1(new_n702), .B2(new_n371), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  AOI21_X1  g510(.A(G36gat), .B1(new_n711), .B2(KEYINPUT46), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n562), .A2(new_n661), .A3(new_n705), .A4(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n711), .A2(KEYINPUT46), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n710), .A2(new_n715), .ZN(G1329gat));
  NAND2_X1  g515(.A1(new_n562), .A2(new_n705), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n317), .B1(new_n717), .B2(new_n675), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n457), .A2(new_n317), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n693), .A2(new_n694), .A3(new_n701), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT47), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n718), .A2(new_n723), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1330gat));
  OAI21_X1  g524(.A(new_n504), .B1(new_n717), .B2(new_n411), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n411), .A2(new_n504), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n693), .A2(new_n694), .A3(new_n701), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n726), .B2(new_n728), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(G1331gat));
  NOR4_X1   g531(.A1(new_n589), .A2(new_n699), .A3(new_n632), .A4(new_n652), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n690), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n442), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n661), .A2(new_n738), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n734), .A2(KEYINPUT108), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT108), .B1(new_n734), .B2(new_n739), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n742), .B(new_n743), .Z(G1333gat));
  OR3_X1    g543(.A1(new_n734), .A2(G71gat), .A3(new_n675), .ZN(new_n745));
  OAI21_X1  g544(.A(G71gat), .B1(new_n734), .B2(new_n457), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g547(.A1(new_n734), .A2(new_n411), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT109), .B(G78gat), .Z(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1335gat));
  NOR3_X1   g550(.A1(new_n696), .A2(new_n652), .A3(new_n699), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n693), .A2(new_n442), .A3(new_n694), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G85gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n696), .A2(new_n699), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n690), .A2(new_n632), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n690), .A2(KEYINPUT51), .A3(new_n632), .A4(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n656), .A2(G85gat), .A3(new_n652), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n754), .A2(KEYINPUT110), .A3(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1336gat));
  NAND4_X1  g566(.A1(new_n693), .A2(new_n661), .A3(new_n694), .A4(new_n752), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n371), .A2(G92gat), .A3(new_n652), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT52), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n769), .A2(new_n774), .A3(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1337gat));
  INV_X1    g575(.A(new_n457), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n695), .A2(new_n777), .A3(new_n752), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT111), .B(G99gat), .Z(new_n779));
  INV_X1    g578(.A(new_n760), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n674), .A2(new_n651), .A3(new_n779), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(G1338gat));
  NAND4_X1  g581(.A1(new_n693), .A2(new_n685), .A3(new_n694), .A4(new_n752), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G106gat), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n411), .A2(G106gat), .A3(new_n652), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n760), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n784), .B2(new_n786), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(G1339gat));
  NOR4_X1   g589(.A1(new_n589), .A2(new_n699), .A3(new_n632), .A4(new_n651), .ZN(new_n791));
  INV_X1    g590(.A(new_n547), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n545), .A2(new_n529), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT115), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n545), .A2(new_n795), .A3(new_n529), .A4(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n489), .B1(new_n550), .B2(new_n529), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n556), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n560), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n560), .A3(KEYINPUT116), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n632), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n640), .A2(new_n641), .A3(new_n635), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n640), .A2(new_n641), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n634), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n640), .A2(KEYINPUT113), .A3(new_n641), .A4(new_n635), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n807), .A2(new_n809), .A3(KEYINPUT54), .A4(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n648), .B1(new_n642), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT114), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n813), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n811), .A2(new_n819), .A3(KEYINPUT55), .A4(new_n813), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n815), .A2(new_n818), .A3(new_n650), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT117), .B1(new_n804), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n821), .ZN(new_n823));
  INV_X1    g622(.A(new_n803), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT116), .B1(new_n799), .B2(new_n560), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n824), .A2(new_n704), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n823), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n651), .A2(new_n560), .A3(new_n799), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n823), .B2(new_n699), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n822), .B(new_n828), .C1(new_n831), .C2(new_n632), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n791), .B1(new_n832), .B2(new_n589), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n833), .A2(new_n656), .A3(new_n414), .ZN(new_n834));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n699), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n833), .A2(new_n685), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n661), .A2(new_n656), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n836), .A2(new_n674), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n213), .B1(new_n559), .B2(new_n560), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(G1340gat));
  AOI21_X1  g639(.A(G120gat), .B1(new_n834), .B2(new_n651), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n652), .A2(new_n215), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n838), .B2(new_n842), .ZN(G1341gat));
  AND2_X1   g642(.A1(new_n203), .A2(new_n205), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n834), .A2(new_n844), .A3(new_n696), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n838), .A2(new_n696), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(new_n844), .ZN(G1342gat));
  AOI21_X1  g646(.A(new_n208), .B1(new_n838), .B2(new_n632), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n834), .A2(new_n208), .A3(new_n632), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(KEYINPUT56), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(KEYINPUT56), .B2(new_n849), .ZN(G1343gat));
  NAND2_X1  g650(.A1(new_n457), .A2(new_n837), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT118), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n823), .A2(new_n699), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n632), .B1(new_n854), .B2(new_n829), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n828), .A2(new_n822), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n589), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n791), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n411), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT119), .B1(new_n859), .B2(KEYINPUT57), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n861), .B(new_n862), .C1(new_n833), .C2(new_n411), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n411), .A2(new_n862), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n820), .A2(new_n650), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n867), .A2(new_n561), .A3(new_n818), .A4(new_n815), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT120), .B1(new_n868), .B2(new_n829), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n815), .A2(new_n650), .A3(new_n820), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n561), .A2(new_n818), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT120), .B(new_n829), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n704), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n856), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n696), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n791), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n829), .B1(new_n870), .B2(new_n871), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n632), .B1(new_n881), .B2(new_n872), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n589), .B1(new_n882), .B2(new_n856), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT121), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n866), .B1(new_n878), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n561), .B(new_n853), .C1(new_n864), .C2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n858), .B1(new_n883), .B2(KEYINPUT121), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n876), .A2(new_n877), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n865), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n860), .A3(new_n863), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n892), .A2(KEYINPUT123), .A3(new_n561), .A4(new_n853), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n888), .A2(G141gat), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n457), .A2(new_n685), .ZN(new_n895));
  NOR4_X1   g694(.A1(new_n833), .A2(new_n895), .A3(new_n656), .A4(new_n661), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n896), .A2(new_n375), .A3(new_n561), .ZN(new_n897));
  XNOR2_X1  g696(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n699), .B(new_n853), .C1(new_n864), .C2(new_n885), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n901), .A2(G141gat), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT58), .B1(new_n902), .B2(new_n897), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(G1344gat));
  NAND3_X1  g703(.A1(new_n896), .A2(new_n377), .A3(new_n651), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n853), .B1(new_n864), .B2(new_n885), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n652), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(KEYINPUT59), .A3(new_n377), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n804), .A2(new_n821), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n589), .B1(new_n882), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n561), .B2(new_n653), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT57), .B1(new_n911), .B2(new_n685), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n833), .A2(new_n866), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n853), .A2(new_n651), .ZN(new_n915));
  OAI21_X1  g714(.A(G148gat), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n905), .B1(new_n908), .B2(new_n918), .ZN(G1345gat));
  OAI21_X1  g718(.A(G155gat), .B1(new_n906), .B2(new_n589), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n896), .A2(new_n583), .A3(new_n696), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1346gat));
  NAND3_X1  g721(.A1(new_n896), .A2(new_n624), .A3(new_n632), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT125), .B1(new_n906), .B2(new_n704), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G162gat), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n906), .A2(KEYINPUT125), .A3(new_n704), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n833), .A2(new_n442), .ZN(new_n928));
  AND4_X1   g727(.A1(new_n661), .A2(new_n928), .A3(new_n411), .A4(new_n674), .ZN(new_n929));
  AOI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n699), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n371), .A2(new_n442), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NOR4_X1   g731(.A1(new_n833), .A2(new_n685), .A3(new_n675), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n262), .B1(new_n559), .B2(new_n560), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G1348gat));
  NAND3_X1  g734(.A1(new_n929), .A2(new_n263), .A3(new_n651), .ZN(new_n936));
  INV_X1    g735(.A(new_n933), .ZN(new_n937));
  OAI21_X1  g736(.A(G176gat), .B1(new_n937), .B2(new_n652), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1349gat));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n589), .A2(new_n243), .A3(new_n299), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n929), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G183gat), .B1(new_n937), .B2(new_n589), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n944), .A2(KEYINPUT60), .ZN(new_n945));
  AND4_X1   g744(.A1(new_n940), .A2(new_n942), .A3(new_n943), .A4(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n942), .A2(new_n943), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT60), .B1(new_n947), .B2(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n940), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(G1350gat));
  AOI21_X1  g749(.A(new_n226), .B1(new_n933), .B2(new_n632), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT61), .Z(new_n952));
  NAND3_X1  g751(.A1(new_n929), .A2(new_n239), .A3(new_n632), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1351gat));
  NOR4_X1   g753(.A1(new_n833), .A2(new_n895), .A3(new_n442), .A4(new_n371), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n699), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n914), .A2(new_n777), .A3(new_n932), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n561), .A2(G197gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(G1352gat));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n332), .A3(new_n651), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT62), .Z(new_n961));
  AND2_X1   g760(.A1(new_n957), .A2(new_n651), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n332), .ZN(G1353gat));
  NAND3_X1  g762(.A1(new_n955), .A2(new_n335), .A3(new_n696), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n777), .A2(new_n932), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n696), .B(new_n965), .C1(new_n912), .C2(new_n913), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n966), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT63), .B1(new_n966), .B2(G211gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(G1354gat));
  NAND3_X1  g768(.A1(new_n955), .A2(new_n336), .A3(new_n632), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n957), .A2(new_n632), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(new_n336), .ZN(G1355gat));
endmodule


