//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G237), .ZN(new_n192));
  INV_X1    g006(.A(G237), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(KEYINPUT68), .ZN(new_n194));
  OAI211_X1 g008(.A(G214), .B(new_n190), .C1(new_n192), .C2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(KEYINPUT68), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n191), .A2(G237), .ZN(new_n199));
  AOI21_X1  g013(.A(G953), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(G143), .B1(new_n200), .B2(G214), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n197), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT84), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT18), .A2(G131), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n195), .A2(new_n196), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n200), .A2(G143), .A3(G214), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n204), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT84), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(new_n209), .ZN(new_n212));
  XNOR2_X1  g026(.A(G125), .B(G140), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n213), .B(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(KEYINPUT16), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n219));
  INV_X1    g033(.A(G140), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G125), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n214), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n218), .A2(G146), .A3(new_n221), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(KEYINPUT17), .B(G131), .C1(new_n197), .C2(new_n201), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT86), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n206), .B2(new_n207), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT86), .B1(new_n231), .B2(KEYINPUT17), .ZN(new_n232));
  OAI211_X1 g046(.A(KEYINPUT87), .B(new_n226), .C1(new_n229), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n208), .A2(G131), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n206), .A2(new_n230), .A3(new_n207), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n227), .A2(new_n228), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n231), .A2(KEYINPUT86), .A3(KEYINPUT17), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n225), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(KEYINPUT87), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n189), .B(new_n217), .C1(new_n240), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n212), .A2(new_n215), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(new_n210), .B2(new_n205), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT19), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n213), .B(new_n248), .ZN(new_n249));
  MUX2_X1   g063(.A(new_n222), .B(new_n249), .S(new_n214), .Z(new_n250));
  AND2_X1   g064(.A1(new_n236), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT85), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n189), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT85), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n236), .A2(new_n250), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n217), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n252), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n245), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n259));
  NOR2_X1   g073(.A1(G475), .A2(G902), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT88), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT88), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n258), .A2(new_n263), .A3(new_n259), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n258), .A2(new_n260), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT20), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT89), .ZN(new_n268));
  INV_X1    g082(.A(G902), .ZN(new_n269));
  OR2_X1    g083(.A1(new_n243), .A2(KEYINPUT87), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n243), .A2(KEYINPUT87), .B1(new_n238), .B2(new_n237), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n247), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(new_n189), .ZN(new_n273));
  INV_X1    g087(.A(new_n245), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G475), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n267), .A2(new_n268), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n268), .B1(new_n267), .B2(new_n276), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G122), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G116), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT90), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G116), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G122), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT91), .ZN(new_n287));
  INV_X1    g101(.A(G107), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(KEYINPUT93), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n286), .A2(KEYINPUT91), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT91), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n291), .B1(new_n283), .B2(new_n285), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n288), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT93), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n283), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n285), .B(KEYINPUT14), .ZN(new_n297));
  OAI21_X1  g111(.A(G107), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n298), .A2(KEYINPUT94), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n196), .A2(G128), .ZN(new_n300));
  INV_X1    g114(.A(G128), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G143), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(G134), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n298), .B2(KEYINPUT94), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n289), .A2(new_n295), .A3(new_n299), .A4(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G134), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n196), .A2(KEYINPUT13), .A3(G128), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n309), .A2(KEYINPUT92), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(KEYINPUT92), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT13), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n300), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n310), .A2(new_n302), .A3(new_n311), .A4(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n308), .B1(new_n314), .B2(G134), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n287), .A2(new_n288), .ZN(new_n316));
  INV_X1    g130(.A(new_n293), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT9), .B(G234), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT74), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n320), .A2(G217), .A3(new_n190), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n306), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(new_n306), .B2(new_n318), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n269), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT15), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G478), .ZN(new_n326));
  INV_X1    g140(.A(G478), .ZN(new_n327));
  OAI221_X1 g141(.A(new_n269), .B1(KEYINPUT15), .B2(new_n327), .C1(new_n322), .C2(new_n323), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n279), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G214), .B1(G237), .B2(G902), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n214), .A2(G143), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n196), .A2(G146), .ZN(new_n335));
  AND2_X1   g149(.A1(KEYINPUT0), .A2(G128), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G143), .B(G146), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT0), .B(G128), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n334), .A2(new_n335), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n334), .A2(KEYINPUT1), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(G128), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n334), .B(new_n335), .C1(KEYINPUT1), .C2(new_n301), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n342), .B1(G125), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT7), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n348), .B1(KEYINPUT82), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n190), .A2(G224), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT7), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n348), .A2(KEYINPUT82), .A3(KEYINPUT7), .A4(new_n351), .ZN(new_n354));
  INV_X1    g168(.A(G119), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G116), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n284), .A2(G119), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT2), .B(G113), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT65), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT65), .B1(new_n356), .B2(new_n357), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT5), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G113), .B1(new_n356), .B2(KEYINPUT5), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G104), .B(G107), .ZN(new_n367));
  INV_X1    g181(.A(G101), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT78), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n288), .A2(G104), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n188), .A2(G107), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(G101), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n288), .A3(G104), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n375), .A2(new_n377), .A3(new_n368), .A4(new_n371), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n369), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n366), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G122), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT8), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT5), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n360), .B1(new_n365), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n380), .B(new_n382), .C1(new_n379), .C2(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n353), .A2(new_n354), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n375), .A2(new_n377), .A3(new_n371), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT76), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n368), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n375), .A2(new_n377), .A3(KEYINPUT76), .A4(new_n371), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT4), .A3(new_n378), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n361), .A2(new_n362), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n360), .B1(new_n393), .B2(new_n359), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n390), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n392), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n379), .A2(KEYINPUT79), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n369), .A2(new_n374), .A3(new_n400), .A4(new_n378), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n366), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n381), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(G902), .B1(new_n386), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n398), .A2(new_n402), .ZN(new_n405));
  INV_X1    g219(.A(new_n381), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n403), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n409), .A3(new_n406), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n348), .B(new_n351), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G210), .B1(G237), .B2(G902), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n404), .A2(new_n412), .A3(new_n414), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(KEYINPUT83), .A3(new_n415), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G952), .ZN(new_n422));
  AOI211_X1 g236(.A(G953), .B(new_n422), .C1(G234), .C2(G237), .ZN(new_n423));
  AOI211_X1 g237(.A(new_n269), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(G898), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR4_X1   g240(.A1(new_n331), .A2(new_n333), .A3(new_n421), .A4(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G472), .A2(G902), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT31), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT11), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n307), .B2(G137), .ZN(new_n431));
  INV_X1    g245(.A(G137), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT11), .A3(G134), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n307), .A2(G137), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G131), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n431), .A2(new_n433), .A3(new_n230), .A4(new_n434), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n341), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n307), .A2(G137), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n432), .A2(G134), .ZN(new_n441));
  OAI21_X1  g255(.A(G131), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n345), .A2(new_n437), .A3(new_n442), .A4(new_n346), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT67), .B1(new_n444), .B2(new_n395), .ZN(new_n445));
  INV_X1    g259(.A(new_n347), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n437), .A2(new_n442), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n446), .A2(new_n447), .B1(new_n438), .B2(new_n341), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT67), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n394), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT30), .B1(new_n444), .B2(KEYINPUT64), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT64), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT30), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n453), .B(new_n454), .C1(new_n439), .C2(new_n443), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n395), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT66), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n451), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n454), .B1(new_n448), .B2(new_n453), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n444), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n394), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(KEYINPUT66), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n200), .A2(G210), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n464), .B(KEYINPUT70), .Z(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT26), .B(G101), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n465), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n429), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n449), .B1(new_n448), .B2(new_n394), .ZN(new_n472));
  AND4_X1   g286(.A1(new_n449), .A2(new_n439), .A3(new_n394), .A4(new_n443), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n461), .B2(KEYINPUT66), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n456), .A2(new_n457), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n475), .A2(new_n429), .A3(new_n470), .A4(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT28), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT71), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n394), .B1(new_n448), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n444), .A2(KEYINPUT71), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n445), .A2(new_n450), .B1(new_n395), .B2(new_n444), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n482), .B1(new_n483), .B2(new_n478), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n469), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n477), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(KEYINPUT32), .B(new_n428), .C1(new_n471), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT72), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n428), .B1(new_n471), .B2(new_n486), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT32), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n475), .A2(new_n470), .A3(new_n476), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT31), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n485), .A3(new_n477), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n428), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n470), .B(new_n482), .C1(new_n483), .C2(new_n478), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n463), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n500), .B2(new_n469), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n269), .B1(new_n497), .B2(new_n498), .ZN(new_n502));
  OAI21_X1  g316(.A(G472), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n489), .A2(new_n492), .A3(new_n496), .A4(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G217), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(G234), .B2(new_n269), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT23), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n355), .B2(G128), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n301), .A2(KEYINPUT23), .A3(G119), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n509), .B(new_n510), .C1(G119), .C2(new_n301), .ZN(new_n511));
  XNOR2_X1  g325(.A(G119), .B(G128), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT24), .B(G110), .Z(new_n513));
  AOI22_X1  g327(.A1(new_n511), .A2(G110), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n225), .A2(new_n514), .ZN(new_n515));
  OAI22_X1  g329(.A1(new_n511), .A2(G110), .B1(new_n512), .B2(new_n513), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n213), .A2(new_n214), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n224), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT22), .B(G137), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(KEYINPUT73), .Z(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n515), .A2(new_n518), .A3(new_n522), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(KEYINPUT25), .A3(new_n269), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT25), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n526), .B2(G902), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n507), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n506), .A2(G902), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n504), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n320), .A2(new_n269), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G221), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT75), .ZN(new_n537));
  INV_X1    g351(.A(G469), .ZN(new_n538));
  XNOR2_X1  g352(.A(G110), .B(G140), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n190), .A2(G227), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n392), .A2(new_n397), .A3(new_n341), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT10), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n379), .B2(new_n347), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n399), .A2(KEYINPUT10), .A3(new_n401), .A4(new_n446), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n438), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT81), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(KEYINPUT81), .A3(new_n438), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n438), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n543), .A2(new_n553), .A3(new_n545), .A4(new_n546), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n542), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n542), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT80), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n379), .A2(new_n347), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n379), .A2(new_n347), .ZN(new_n559));
  OAI221_X1 g373(.A(new_n438), .B1(new_n557), .B2(KEYINPUT12), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n438), .B1(new_n558), .B2(new_n559), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT12), .B1(new_n438), .B2(new_n557), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n556), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n538), .B(new_n269), .C1(new_n555), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n560), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n542), .B1(new_n566), .B2(new_n554), .ZN(new_n567));
  INV_X1    g381(.A(new_n556), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n567), .B1(new_n552), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G469), .B1(new_n569), .B2(G902), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n537), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n534), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n427), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G101), .ZN(G3));
  OAI21_X1  g389(.A(KEYINPUT95), .B1(new_n322), .B2(new_n323), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(KEYINPUT95), .B(KEYINPUT33), .C1(new_n322), .C2(new_n323), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(G478), .A3(new_n269), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n324), .A2(new_n327), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n267), .A2(new_n276), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT89), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n267), .A2(new_n268), .A3(new_n276), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n583), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n426), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n333), .B1(new_n416), .B2(new_n418), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n495), .A2(new_n269), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n571), .A2(new_n592), .A3(new_n490), .A4(new_n533), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT34), .B(G104), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G6));
  NAND2_X1  g410(.A1(new_n266), .A2(new_n261), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n276), .ZN(new_n598));
  INV_X1    g412(.A(new_n589), .ZN(new_n599));
  NOR4_X1   g413(.A1(new_n598), .A2(new_n599), .A3(new_n330), .A4(new_n426), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n592), .A2(new_n490), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n572), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n602), .A3(new_n533), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G107), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  OR2_X1    g419(.A1(new_n523), .A2(KEYINPUT36), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n519), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n532), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n528), .A2(new_n530), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n507), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n607), .A2(G902), .A3(new_n506), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT96), .B1(new_n613), .B2(new_n531), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n602), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n427), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT37), .B(G110), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G12));
  AND4_X1   g433(.A1(new_n504), .A2(new_n571), .A3(new_n589), .A4(new_n615), .ZN(new_n620));
  INV_X1    g434(.A(G900), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n424), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n423), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n598), .A2(new_n330), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G128), .ZN(G30));
  XOR2_X1   g442(.A(new_n421), .B(KEYINPUT38), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n624), .B(KEYINPUT39), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n571), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n631), .A2(KEYINPUT40), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n585), .A2(new_n586), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n483), .B2(new_n469), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n463), .B2(new_n469), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n489), .A2(new_n492), .A3(new_n496), .A4(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n329), .A2(new_n332), .ZN(new_n639));
  AOI211_X1 g453(.A(new_n615), .B(new_n639), .C1(new_n631), .C2(KEYINPUT40), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n633), .A2(new_n634), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G143), .ZN(G45));
  NAND3_X1  g456(.A1(new_n620), .A2(new_n587), .A3(new_n624), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G146), .ZN(G48));
  INV_X1    g458(.A(new_n534), .ZN(new_n645));
  INV_X1    g459(.A(new_n551), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT81), .B1(new_n547), .B2(new_n438), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n554), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n564), .B1(new_n648), .B2(new_n541), .ZN(new_n649));
  OAI21_X1  g463(.A(G469), .B1(new_n649), .B2(G902), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n536), .A3(new_n565), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n590), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT41), .B(G113), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G15));
  NAND3_X1  g470(.A1(new_n645), .A2(new_n600), .A3(new_n652), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G116), .ZN(G18));
  NOR2_X1   g472(.A1(new_n634), .A2(new_n329), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n504), .A2(new_n615), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n589), .A2(new_n650), .A3(new_n536), .A4(new_n565), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n659), .A2(new_n588), .A3(new_n660), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G119), .ZN(G21));
  NOR2_X1   g478(.A1(new_n651), .A2(new_n426), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n428), .B(KEYINPUT97), .Z(new_n666));
  AOI22_X1  g480(.A1(new_n591), .A2(G472), .B1(new_n495), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n667), .A2(new_n533), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n589), .A2(new_n329), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n634), .A2(new_n665), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G122), .ZN(G24));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n581), .A2(new_n582), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n674), .B(new_n624), .C1(new_n277), .C2(new_n278), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n495), .A2(new_n666), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n592), .A2(new_n615), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n662), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n673), .B1(new_n675), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n677), .A2(new_n661), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n587), .A2(KEYINPUT98), .A3(new_n624), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G125), .ZN(G27));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n333), .B1(new_n419), .B2(new_n420), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT99), .ZN(new_n687));
  INV_X1    g501(.A(new_n536), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n565), .B2(new_n570), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n645), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n685), .B1(new_n690), .B2(new_n675), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT99), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n686), .A2(new_n692), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n693), .A2(new_n694), .A3(new_n689), .ZN(new_n695));
  INV_X1    g509(.A(new_n675), .ZN(new_n696));
  INV_X1    g510(.A(new_n533), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT32), .B1(new_n495), .B2(new_n428), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n698), .A2(KEYINPUT101), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n503), .B1(new_n698), .B2(KEYINPUT101), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n487), .B(KEYINPUT100), .Z(new_n702));
  AOI21_X1  g516(.A(new_n697), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n695), .A2(new_n696), .A3(new_n703), .A4(KEYINPUT42), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n691), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G131), .ZN(G33));
  INV_X1    g520(.A(new_n626), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n690), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n307), .ZN(G36));
  NOR2_X1   g523(.A1(new_n634), .A2(new_n583), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT43), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n601), .A2(new_n615), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n713), .A2(KEYINPUT44), .A3(new_n714), .A4(new_n715), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n687), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT104), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n569), .A2(KEYINPUT45), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n569), .A2(KEYINPUT45), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(G469), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(G469), .A2(G902), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT46), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n565), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n724), .A2(KEYINPUT46), .A3(new_n725), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n688), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n630), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT102), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n721), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT105), .B(G137), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G39));
  XNOR2_X1  g549(.A(new_n730), .B(KEYINPUT47), .ZN(new_n736));
  INV_X1    g550(.A(new_n687), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n737), .A2(new_n504), .A3(new_n533), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(new_n696), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT106), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G140), .ZN(G42));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n711), .A2(new_n423), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n737), .A2(new_n651), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n678), .A3(new_n744), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n638), .A2(new_n623), .A3(new_n697), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n279), .A2(new_n583), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n743), .A2(new_n668), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n629), .A2(new_n332), .A3(new_n651), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(KEYINPUT50), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n743), .A2(new_n668), .A3(new_n751), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n749), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(KEYINPUT114), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n650), .A2(new_n565), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT107), .ZN(new_n759));
  INV_X1    g573(.A(new_n537), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n750), .B(new_n687), .C1(new_n736), .C2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n756), .B2(KEYINPUT114), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n742), .B1(new_n757), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT115), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n756), .A2(KEYINPUT51), .A3(new_n762), .ZN(new_n766));
  INV_X1    g580(.A(new_n587), .ZN(new_n767));
  OAI211_X1 g581(.A(G952), .B(new_n190), .C1(new_n747), .C2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n750), .B2(new_n662), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n743), .A2(new_n703), .A3(new_n744), .ZN(new_n770));
  NAND2_X1  g584(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OR2_X1    g586(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n769), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n765), .A2(new_n766), .A3(new_n775), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n593), .A2(new_n333), .A3(new_n421), .A4(new_n426), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n634), .A2(new_n583), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n331), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n663), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n657), .B(new_n671), .C1(new_n590), .C2(new_n653), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n708), .B1(new_n691), .B2(new_n704), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n427), .B1(new_n573), .B2(new_n616), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n660), .A2(new_n571), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n329), .A2(new_n625), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n597), .A3(KEYINPUT109), .A4(new_n276), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n788));
  INV_X1    g602(.A(new_n786), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n788), .B1(new_n789), .B2(new_n598), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n687), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n687), .A2(new_n678), .A3(new_n689), .ZN(new_n792));
  OAI22_X1  g606(.A1(new_n785), .A2(new_n791), .B1(new_n792), .B2(new_n675), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n504), .A2(new_n571), .A3(new_n589), .A4(new_n615), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n675), .B2(new_n707), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n565), .A2(new_n570), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n613), .A2(new_n531), .A3(new_n625), .ZN(new_n800));
  AND4_X1   g614(.A1(KEYINPUT110), .A2(new_n799), .A3(new_n536), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT110), .B1(new_n689), .B2(new_n800), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n638), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n670), .B1(new_n277), .B2(new_n278), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n798), .A2(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n806), .A2(KEYINPUT111), .A3(new_n683), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT111), .B1(new_n806), .B2(new_n683), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n796), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT111), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n680), .A2(new_n682), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n689), .A2(new_n800), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n689), .A2(KEYINPUT110), .A3(new_n800), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n634), .A3(new_n638), .A4(new_n670), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n643), .A2(new_n627), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n810), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n806), .A2(new_n683), .A3(KEYINPUT111), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(KEYINPUT52), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n795), .A2(new_n809), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT52), .B1(new_n819), .B2(new_n820), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n796), .B1(new_n806), .B2(new_n683), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n827), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT112), .B1(new_n809), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n795), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n824), .B1(new_n831), .B2(new_n823), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT113), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n807), .A2(new_n808), .A3(new_n796), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n794), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT53), .B1(new_n837), .B2(new_n809), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n826), .B1(new_n825), .B2(new_n827), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n809), .A2(KEYINPUT112), .A3(new_n829), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n838), .B1(KEYINPUT53), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n833), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n841), .A2(KEYINPUT53), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n844), .B(KEYINPUT54), .C1(new_n845), .C2(new_n824), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n834), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  OAI22_X1  g661(.A1(new_n776), .A2(new_n847), .B1(G952), .B2(G953), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n533), .A2(new_n332), .A3(new_n760), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n629), .A2(new_n583), .A3(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n638), .B(new_n850), .C1(KEYINPUT49), .C2(new_n759), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n759), .A2(KEYINPUT49), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT108), .Z(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n279), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n848), .A2(new_n854), .ZN(G75));
  NOR2_X1   g669(.A1(new_n842), .A2(new_n269), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT56), .B1(new_n856), .B2(G210), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n408), .A2(new_n410), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(new_n411), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT55), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n857), .A2(new_n860), .B1(G952), .B2(new_n190), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n857), .B2(new_n860), .ZN(G51));
  NOR2_X1   g676(.A1(new_n190), .A2(G952), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n831), .A2(new_n823), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n864), .B(KEYINPUT54), .C1(new_n865), .C2(new_n838), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT117), .B1(new_n842), .B2(new_n833), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n843), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n725), .B(KEYINPUT57), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n869), .A2(new_n870), .B1(new_n555), .B2(new_n564), .ZN(new_n871));
  OR3_X1    g685(.A1(new_n842), .A2(new_n269), .A3(new_n724), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n863), .B1(new_n871), .B2(new_n872), .ZN(G54));
  NAND3_X1  g687(.A1(new_n856), .A2(KEYINPUT58), .A3(G475), .ZN(new_n874));
  INV_X1    g688(.A(new_n258), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n863), .B1(new_n874), .B2(new_n875), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G60));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n882));
  NAND2_X1  g696(.A1(G478), .A2(G902), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT59), .Z(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n578), .B2(new_n579), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n863), .B1(new_n868), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n884), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n580), .B1(new_n847), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI211_X1 g704(.A(KEYINPUT119), .B(new_n580), .C1(new_n847), .C2(new_n887), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n882), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n831), .A2(new_n823), .ZN(new_n893));
  INV_X1    g707(.A(new_n824), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n833), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n895), .A2(new_n844), .B1(new_n833), .B2(new_n842), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n884), .B1(new_n896), .B2(new_n834), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT119), .B1(new_n897), .B2(new_n580), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n888), .A2(new_n889), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(KEYINPUT120), .A3(new_n899), .A4(new_n886), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n892), .A2(new_n900), .ZN(G63));
  NAND2_X1  g715(.A1(G217), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT121), .Z(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT60), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n842), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n863), .B1(new_n905), .B2(new_n608), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n526), .B(KEYINPUT122), .Z(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT61), .Z(G66));
  INV_X1    g723(.A(new_n425), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n190), .B1(new_n910), .B2(G224), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n782), .A2(new_n784), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(new_n190), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n858), .B1(G898), .B2(new_n190), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n913), .B(new_n914), .Z(G69));
  NAND2_X1  g729(.A1(new_n459), .A2(new_n460), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n249), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n331), .A2(new_n778), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n737), .A2(new_n534), .A3(new_n631), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n740), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n811), .A2(new_n798), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n641), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n925), .B1(KEYINPUT62), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(KEYINPUT62), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT123), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n733), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n918), .B1(new_n933), .B2(new_n190), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n917), .B1(G900), .B2(G953), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n732), .A2(new_n634), .A3(new_n670), .A4(new_n703), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT125), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n938), .A2(new_n740), .A3(new_n783), .A4(new_n926), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n721), .B2(new_n732), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n940), .B2(new_n190), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT126), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n931), .B1(new_n721), .B2(new_n732), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n917), .B1(new_n944), .B2(G953), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n940), .A2(new_n190), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n943), .B(new_n945), .C1(new_n946), .C2(new_n936), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n942), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n948), .ZN(new_n950));
  OAI211_X1 g764(.A(KEYINPUT126), .B(new_n950), .C1(new_n934), .C2(new_n941), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(G72));
  NAND3_X1  g766(.A1(new_n944), .A2(new_n782), .A3(new_n784), .ZN(new_n953));
  NAND2_X1  g767(.A1(G472), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT63), .Z(new_n955));
  AOI211_X1 g769(.A(new_n469), .B(new_n463), .C1(new_n953), .C2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n940), .A2(new_n782), .A3(new_n784), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n470), .B(new_n500), .C1(new_n957), .C2(new_n955), .ZN(new_n958));
  INV_X1    g772(.A(new_n955), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n500), .A2(new_n469), .ZN(new_n960));
  AOI211_X1 g774(.A(new_n959), .B(new_n832), .C1(new_n493), .C2(new_n960), .ZN(new_n961));
  NOR4_X1   g775(.A1(new_n956), .A2(new_n958), .A3(new_n863), .A4(new_n961), .ZN(G57));
endmodule


