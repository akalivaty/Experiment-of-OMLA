//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT11), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n187), .B(new_n192), .C1(new_n188), .C2(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n196), .A3(new_n191), .A4(new_n193), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(KEYINPUT66), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n199), .A3(G131), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n198), .A2(KEYINPUT67), .A3(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT67), .B1(new_n198), .B2(new_n200), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT76), .B(G101), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n204), .A2(new_n206), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n206), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n205), .A2(G107), .ZN(new_n213));
  OAI211_X1 g027(.A(KEYINPUT77), .B(G101), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G143), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(new_n220), .A3(G143), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n218), .B(G146), .C1(new_n216), .C2(KEYINPUT1), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n212), .B2(new_n213), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n215), .A2(KEYINPUT10), .A3(new_n225), .A4(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n228), .A2(new_n225), .A3(new_n211), .A4(new_n214), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT10), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n210), .A2(new_n209), .A3(new_n206), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G101), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(KEYINPUT75), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(KEYINPUT75), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n233), .A2(G101), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n233), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n236), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  XOR2_X1   g055(.A(KEYINPUT0), .B(G128), .Z(new_n242));
  XNOR2_X1  g056(.A(G143), .B(G146), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT0), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n245), .B2(new_n216), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n229), .B(new_n232), .C1(new_n241), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n203), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n236), .A2(new_n238), .A3(new_n240), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n244), .A2(new_n246), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n250), .A2(new_n251), .B1(new_n231), .B2(new_n230), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n252), .B(new_n229), .C1(new_n201), .C2(new_n202), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G953), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT68), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G227), .ZN(new_n261));
  XNOR2_X1  g075(.A(G110), .B(G140), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT78), .B1(new_n254), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n228), .A2(new_n211), .A3(new_n214), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n230), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT12), .B1(new_n203), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(KEYINPUT12), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n198), .A2(new_n200), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n253), .B(new_n263), .C1(new_n270), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n268), .A2(new_n230), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n201), .A2(new_n276), .A3(new_n202), .ZN(new_n277));
  OAI22_X1  g091(.A1(new_n277), .A2(KEYINPUT12), .B1(new_n272), .B2(new_n271), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n278), .A2(KEYINPUT78), .A3(new_n253), .A4(new_n263), .ZN(new_n279));
  INV_X1    g093(.A(G469), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n275), .A2(new_n279), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n253), .B(new_n264), .C1(new_n270), .C2(new_n273), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n249), .A2(new_n253), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(new_n264), .ZN(new_n286));
  OAI21_X1  g100(.A(G469), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n280), .A2(new_n281), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n282), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  XOR2_X1   g104(.A(KEYINPUT9), .B(G234), .Z(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G221), .B1(new_n292), .B2(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G210), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G119), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G116), .ZN(new_n298));
  INV_X1    g112(.A(G116), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G119), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT2), .B(G113), .Z(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(new_n300), .A3(KEYINPUT5), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n304), .B(G113), .C1(KEYINPUT5), .C2(new_n298), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n215), .A2(new_n303), .A3(new_n228), .A4(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n301), .B(new_n302), .Z(new_n307));
  OAI21_X1  g121(.A(new_n306), .B1(new_n241), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G110), .B(G122), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n306), .B(new_n309), .C1(new_n241), .C2(new_n307), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(KEYINPUT6), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n247), .A2(G125), .ZN(new_n314));
  INV_X1    g128(.A(G125), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n267), .A2(KEYINPUT79), .A3(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n222), .A2(new_n315), .A3(new_n223), .A4(new_n224), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G224), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(G953), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT6), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n308), .A2(new_n325), .A3(new_n310), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n313), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n281), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n317), .A2(new_n318), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n317), .A2(new_n318), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n316), .A2(KEYINPUT81), .A3(new_n319), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n314), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n323), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT82), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n336), .A2(KEYINPUT7), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(KEYINPUT7), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n334), .A2(KEYINPUT83), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT83), .B1(new_n334), .B2(new_n339), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n312), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n305), .A2(new_n303), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n266), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n306), .A2(new_n344), .A3(KEYINPUT80), .ZN(new_n345));
  OR3_X1    g159(.A1(new_n266), .A2(new_n343), .A3(KEYINPUT80), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n309), .B(KEYINPUT8), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n314), .A2(KEYINPUT7), .A3(new_n320), .A4(new_n335), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n296), .B1(new_n328), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n348), .A2(new_n349), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n354), .B(new_n312), .C1(new_n341), .C2(new_n340), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n355), .A2(new_n281), .A3(new_n295), .A4(new_n327), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n356), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT84), .ZN(new_n359));
  OAI21_X1  g173(.A(G214), .B1(G237), .B2(G902), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n257), .A2(G952), .ZN(new_n362));
  INV_X1    g176(.A(G234), .ZN(new_n363));
  INV_X1    g177(.A(G237), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  XOR2_X1   g180(.A(KEYINPUT21), .B(G898), .Z(new_n367));
  OAI21_X1  g181(.A(G902), .B1(new_n363), .B2(new_n364), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n369), .B2(new_n259), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n294), .A2(new_n361), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT67), .ZN(new_n372));
  INV_X1    g186(.A(G137), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G134), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n192), .B1(new_n374), .B2(new_n187), .ZN(new_n375));
  AOI211_X1 g189(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n373), .C2(G134), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n196), .B1(new_n377), .B2(new_n191), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n197), .A2(KEYINPUT66), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n200), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n372), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n198), .A2(KEYINPUT67), .A3(new_n200), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n251), .A3(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n191), .A2(new_n374), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n197), .B(new_n225), .C1(new_n196), .C2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(KEYINPUT30), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n307), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n272), .B2(new_n247), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n384), .A2(new_n307), .A3(new_n386), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n257), .A2(KEYINPUT68), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n255), .A2(G953), .ZN(new_n395));
  AOI21_X1  g209(.A(G237), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G210), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(G101), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n392), .A2(new_n393), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT31), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n392), .A2(new_n393), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n393), .A2(KEYINPUT28), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT28), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n384), .A2(new_n406), .A3(new_n307), .A4(new_n386), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n405), .A2(new_n407), .B1(new_n388), .B2(new_n389), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n402), .B(new_n404), .C1(new_n400), .C2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(G472), .A2(G902), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT32), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n405), .A2(new_n407), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n389), .A2(new_n388), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n400), .ZN(new_n417));
  INV_X1    g231(.A(new_n400), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n392), .A2(new_n393), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT29), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n307), .B1(new_n384), .B2(new_n386), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n405), .B2(new_n407), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT29), .A3(new_n400), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n281), .ZN(new_n424));
  OAI21_X1  g238(.A(G472), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n409), .A2(KEYINPUT32), .A3(new_n410), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n413), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT22), .B(G137), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n216), .A2(KEYINPUT23), .A3(G119), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT70), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n297), .A2(G128), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n216), .A2(G119), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT23), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G110), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n433), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT24), .B(G110), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G140), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G125), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n315), .A2(G140), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT71), .A3(KEYINPUT16), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT71), .B1(new_n443), .B2(KEYINPUT16), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT16), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n450), .A3(G146), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(G146), .B1(new_n447), .B2(new_n450), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n438), .B(new_n441), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n439), .A2(new_n440), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(new_n437), .B2(G110), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n446), .A2(new_n220), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT72), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n454), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n454), .B2(new_n458), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n430), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n430), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n454), .A2(new_n458), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n463), .B1(new_n464), .B2(KEYINPUT72), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n281), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n469));
  INV_X1    g283(.A(new_n467), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n462), .A2(new_n281), .A3(new_n465), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G217), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(G234), .B2(new_n281), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(G902), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n462), .A2(new_n465), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT74), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G475), .ZN(new_n481));
  OAI211_X1 g295(.A(G214), .B(new_n364), .C1(new_n256), .C2(new_n258), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n218), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n396), .A2(G143), .A3(G214), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n196), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT17), .ZN(new_n488));
  INV_X1    g302(.A(new_n484), .ZN(new_n489));
  AOI21_X1  g303(.A(G143), .B1(new_n396), .B2(G214), .ZN(new_n490));
  OAI21_X1  g304(.A(G131), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n483), .A2(KEYINPUT85), .A3(new_n484), .A4(new_n196), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n487), .A2(new_n488), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n452), .A2(new_n453), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n483), .A2(new_n484), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT17), .A3(G131), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(G113), .B(G122), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n205), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n445), .B(G146), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(new_n196), .ZN(new_n502));
  OAI221_X1 g316(.A(new_n500), .B1(new_n495), .B2(new_n502), .C1(new_n491), .C2(new_n501), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT86), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n497), .A2(new_n506), .A3(new_n499), .A4(new_n503), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT88), .B1(new_n497), .B2(new_n503), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n497), .A2(KEYINPUT88), .A3(new_n503), .ZN(new_n510));
  INV_X1    g324(.A(new_n499), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n508), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n481), .B1(new_n513), .B2(new_n281), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n487), .A2(new_n491), .A3(new_n492), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n445), .B(KEYINPUT19), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n516), .B(new_n451), .C1(G146), .C2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n499), .B1(new_n518), .B2(new_n503), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n505), .B2(new_n507), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n519), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n508), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT87), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT87), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n525), .A2(new_n529), .A3(new_n527), .A4(new_n521), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n515), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(G128), .B(G143), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT13), .ZN(new_n534));
  OR3_X1    g348(.A1(new_n216), .A2(KEYINPUT13), .A3(G143), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(G134), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G122), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G116), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n299), .A2(G122), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G107), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n539), .A3(new_n208), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n533), .A2(new_n188), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n536), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n541), .A2(new_n542), .B1(new_n188), .B2(new_n533), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(KEYINPUT89), .A3(new_n536), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n539), .A2(KEYINPUT14), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n538), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT90), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n208), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT90), .B1(new_n539), .B2(KEYINPUT14), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n533), .B(new_n188), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n542), .A3(new_n557), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n292), .A2(new_n473), .A3(G953), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n550), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT91), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n550), .A2(new_n558), .A3(new_n559), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n559), .B1(new_n550), .B2(new_n558), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n562), .B1(new_n565), .B2(new_n561), .ZN(new_n566));
  INV_X1    g380(.A(G478), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT92), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n566), .A2(KEYINPUT93), .A3(new_n281), .A4(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n549), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT89), .B1(new_n548), .B2(new_n536), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n558), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n559), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(new_n561), .A3(new_n560), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n563), .A2(KEYINPUT91), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n281), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT93), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n572), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n580), .A2(KEYINPUT93), .A3(new_n581), .A4(new_n281), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n574), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n532), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n371), .A2(new_n427), .A3(new_n480), .A4(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(new_n589), .B(new_n204), .Z(G3));
  INV_X1    g404(.A(G472), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n409), .B2(new_n281), .ZN(new_n592));
  INV_X1    g406(.A(new_n410), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n416), .A2(new_n418), .B1(new_n401), .B2(KEYINPUT31), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n594), .B2(new_n404), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n592), .A2(new_n479), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n529), .B1(new_n508), .B2(new_n524), .ZN(new_n597));
  OAI22_X1  g411(.A1(new_n597), .A2(KEYINPUT20), .B1(new_n520), .B2(new_n522), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n514), .B1(new_n598), .B2(new_n530), .ZN(new_n599));
  INV_X1    g413(.A(new_n370), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n327), .A2(new_n281), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n295), .B1(new_n601), .B2(new_n355), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n360), .B(new_n600), .C1(new_n602), .C2(new_n358), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT94), .B(KEYINPUT33), .Z(new_n604));
  NAND3_X1  g418(.A1(new_n565), .A2(KEYINPUT95), .A3(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n579), .A2(KEYINPUT33), .A3(new_n560), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n566), .A2(new_n604), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n567), .A2(G902), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n609), .A2(new_n610), .B1(new_n567), .B2(new_n582), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n599), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n294), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n596), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT34), .B(G104), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NAND2_X1  g430(.A1(new_n596), .A2(new_n613), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n520), .B2(new_n522), .ZN(new_n619));
  INV_X1    g433(.A(new_n618), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n523), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n515), .A2(new_n619), .A3(new_n587), .A4(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n617), .A2(new_n603), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT35), .B(G107), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G9));
  NOR2_X1   g439(.A1(new_n463), .A2(KEYINPUT36), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(new_n464), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n472), .A2(new_n474), .B1(new_n476), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n371), .A2(new_n588), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(G902), .B1(new_n594), .B2(new_n404), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n411), .B1(new_n631), .B2(new_n591), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT37), .B(G110), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  INV_X1    g449(.A(G900), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n259), .A2(new_n636), .ZN(new_n637));
  OR3_X1    g451(.A1(new_n637), .A2(KEYINPUT97), .A3(new_n368), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT97), .B1(new_n637), .B2(new_n368), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n365), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n622), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n360), .B1(new_n602), .B2(new_n358), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n294), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n427), .A2(new_n642), .A3(new_n629), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  XNOR2_X1  g460(.A(new_n640), .B(KEYINPUT39), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n613), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(KEYINPUT40), .ZN(new_n649));
  INV_X1    g463(.A(new_n587), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n649), .A2(new_n599), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n357), .A2(new_n359), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT38), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n629), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n418), .B1(new_n392), .B2(new_n393), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n393), .A2(new_n418), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n281), .B1(new_n656), .B2(new_n421), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n413), .A2(new_n658), .A3(new_n426), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(KEYINPUT40), .B2(new_n648), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n651), .A2(new_n360), .A3(new_n654), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G143), .ZN(G45));
  NOR3_X1   g477(.A1(new_n599), .A2(new_n611), .A3(new_n641), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n427), .A2(new_n664), .A3(new_n629), .A4(new_n644), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  NAND3_X1  g480(.A1(new_n275), .A2(new_n279), .A3(new_n281), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G469), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(new_n293), .A3(new_n282), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n427), .A2(new_n612), .A3(new_n480), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT41), .B(G113), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G15));
  NOR2_X1   g487(.A1(new_n622), .A2(new_n643), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n669), .A2(new_n370), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n427), .A2(new_n674), .A3(new_n480), .A4(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT98), .B(G116), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G18));
  NOR3_X1   g492(.A1(new_n669), .A2(new_n643), .A3(new_n628), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n427), .A2(new_n679), .A3(new_n588), .A4(new_n600), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  INV_X1    g495(.A(new_n643), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n532), .A2(new_n682), .A3(new_n587), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n598), .A2(new_n530), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n650), .B1(new_n686), .B2(new_n515), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(KEYINPUT101), .A3(new_n682), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT100), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n631), .B2(new_n591), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n409), .A2(new_n281), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(KEYINPUT100), .A3(G472), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n402), .B1(new_n400), .B2(new_n422), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT99), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n402), .B(KEYINPUT99), .C1(new_n400), .C2(new_n422), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n404), .A3(new_n697), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n691), .A2(new_n693), .B1(new_n698), .B2(new_n410), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n689), .A2(new_n480), .A3(new_n675), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G122), .ZN(G24));
  AOI21_X1  g515(.A(new_n611), .B1(new_n686), .B2(new_n515), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT102), .B1(new_n702), .B2(new_n640), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n599), .A2(new_n704), .A3(new_n611), .A4(new_n641), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n699), .B(new_n679), .C1(new_n703), .C2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT103), .B(G125), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G27));
  INV_X1    g522(.A(new_n611), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n532), .A2(new_n709), .A3(new_n640), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n704), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n702), .A2(KEYINPUT102), .A3(new_n640), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n652), .A2(new_n360), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n294), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n716));
  AOI211_X1 g530(.A(new_n412), .B(new_n593), .C1(new_n594), .C2(new_n404), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT32), .B1(new_n409), .B2(new_n410), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n413), .A2(KEYINPUT104), .A3(new_n426), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n425), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n713), .A2(new_n480), .A3(new_n715), .A4(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n717), .A2(new_n718), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n479), .B1(new_n723), .B2(new_n425), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n724), .A2(new_n715), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT42), .B1(new_n711), .B2(new_n712), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n722), .A2(KEYINPUT42), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G131), .ZN(G33));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n724), .A2(new_n729), .A3(new_n642), .A4(new_n715), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n715), .A2(new_n427), .A3(new_n642), .A4(new_n480), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT105), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  NAND2_X1  g548(.A1(new_n599), .A2(new_n709), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT43), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n599), .A2(new_n737), .A3(new_n709), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n632), .A3(new_n629), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n714), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n739), .A2(KEYINPUT44), .A3(new_n632), .A4(new_n629), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT45), .B1(new_n284), .B2(new_n286), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n283), .B(new_n747), .C1(new_n264), .C2(new_n285), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(G469), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n746), .A2(KEYINPUT106), .A3(new_n748), .A4(G469), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n289), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT107), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n289), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n753), .A2(new_n759), .A3(KEYINPUT46), .A4(new_n289), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n755), .A2(new_n758), .A3(new_n282), .A4(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(new_n293), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n762), .A2(KEYINPUT108), .A3(new_n647), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT108), .B1(new_n762), .B2(new_n647), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n745), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G137), .ZN(G39));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n761), .A2(new_n767), .A3(new_n293), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n767), .B1(new_n761), .B2(new_n293), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR4_X1   g584(.A1(new_n427), .A2(new_n710), .A3(new_n480), .A4(new_n714), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT109), .Z(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  INV_X1    g588(.A(KEYINPUT120), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n722), .A2(KEYINPUT42), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n725), .A2(new_n726), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n733), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n671), .A2(new_n680), .A3(new_n676), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n587), .B(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(new_n599), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n371), .B(new_n596), .C1(new_n782), .C2(new_n702), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(new_n589), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n630), .A2(new_n632), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n779), .A2(new_n784), .A3(new_n700), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n699), .B1(new_n703), .B2(new_n705), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n781), .A2(new_n641), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n515), .A2(new_n619), .A3(new_n621), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n427), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n791), .A2(new_n629), .A3(new_n715), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n778), .A2(new_n786), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n627), .A2(new_n476), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n475), .A2(new_n795), .A3(new_n640), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n628), .A2(KEYINPUT113), .A3(new_n640), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n294), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT101), .B1(new_n687), .B2(new_n682), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n599), .A2(new_n643), .A3(new_n684), .A4(new_n650), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n659), .B(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n706), .A2(new_n803), .A3(new_n645), .A4(new_n665), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n645), .A2(new_n665), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n806), .A2(new_n807), .A3(new_n706), .A4(new_n803), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n794), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n805), .A2(new_n794), .A3(new_n808), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n793), .B(KEYINPUT53), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n812));
  XNOR2_X1  g626(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n675), .B1(new_n801), .B2(new_n802), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n699), .A2(new_n480), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n589), .B(new_n783), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n671), .A2(new_n680), .A3(new_n676), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n817), .A2(new_n633), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n791), .A2(new_n629), .A3(new_n715), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n727), .A3(new_n733), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n805), .A2(new_n808), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n814), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n811), .A2(new_n812), .A3(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n821), .A2(new_n822), .A3(new_n814), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n793), .B1(new_n810), .B2(new_n809), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n824), .B1(new_n828), .B2(new_n812), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n736), .A2(new_n366), .A3(new_n738), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n830), .A2(new_n669), .A3(new_n714), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n480), .A3(new_n721), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT48), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n816), .A2(new_n830), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n682), .A3(new_n670), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n480), .A2(new_n366), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n659), .A2(new_n836), .A3(new_n669), .A4(new_n714), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n702), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n833), .A2(new_n362), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n669), .A2(KEYINPUT117), .A3(new_n360), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT117), .B1(new_n669), .B2(new_n360), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n653), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n834), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(KEYINPUT119), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n816), .A2(new_n843), .A3(new_n830), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n849), .B1(new_n850), .B2(new_n846), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(KEYINPUT50), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n848), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n831), .A2(new_n629), .A3(new_n699), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n837), .A2(new_n599), .A3(new_n611), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(KEYINPUT116), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n668), .A2(new_n282), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n293), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n743), .B(new_n834), .C1(new_n770), .C2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n856), .A3(new_n853), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n853), .A2(new_n856), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n865), .A2(new_n862), .B1(new_n857), .B2(new_n858), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n840), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n775), .B1(new_n829), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n827), .A2(new_n826), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT54), .B1(new_n869), .B2(new_n825), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n859), .A2(new_n863), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n865), .A2(new_n858), .A3(new_n857), .A4(new_n862), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n839), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n870), .A2(new_n873), .A3(KEYINPUT120), .A4(new_n824), .ZN(new_n874));
  NOR2_X1   g688(.A1(G952), .A2(G953), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT121), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n868), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n735), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n480), .A3(new_n293), .A4(new_n360), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT110), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n879), .A2(new_n880), .B1(KEYINPUT49), .B2(new_n860), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n880), .B2(new_n879), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT111), .Z(new_n883));
  OR2_X1    g697(.A1(new_n860), .A2(KEYINPUT49), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n653), .A3(new_n660), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n877), .A2(new_n885), .ZN(G75));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n811), .A2(new_n823), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n887), .B1(new_n888), .B2(G902), .ZN(new_n889));
  AOI211_X1 g703(.A(KEYINPUT122), .B(new_n281), .C1(new_n811), .C2(new_n823), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n296), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n313), .A2(new_n326), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n324), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT55), .Z(new_n894));
  XNOR2_X1  g708(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n260), .A2(G952), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n888), .A2(G210), .A3(G902), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n894), .B1(new_n900), .B2(KEYINPUT56), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n897), .A2(new_n899), .A3(new_n901), .ZN(G51));
  NAND2_X1  g716(.A1(new_n289), .A2(KEYINPUT57), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n289), .A2(KEYINPUT57), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n811), .A2(new_n812), .A3(new_n823), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n812), .B1(new_n811), .B2(new_n823), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n903), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n275), .A3(new_n279), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n751), .B(new_n752), .C1(new_n889), .C2(new_n890), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n898), .B1(new_n908), .B2(new_n909), .ZN(G54));
  AND2_X1   g724(.A1(KEYINPUT58), .A2(G475), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n889), .B2(new_n890), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n520), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n525), .B(new_n911), .C1(new_n889), .C2(new_n890), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n913), .A2(new_n899), .A3(new_n914), .ZN(G60));
  INV_X1    g729(.A(new_n609), .ZN(new_n916));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT59), .Z(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n905), .B2(new_n906), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n920), .A2(KEYINPUT124), .A3(new_n899), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT124), .B1(new_n920), .B2(new_n899), .ZN(new_n922));
  INV_X1    g736(.A(new_n918), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n609), .B1(new_n829), .B2(new_n923), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(G63));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT60), .Z(new_n927));
  AND2_X1   g741(.A1(new_n888), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n898), .B1(new_n928), .B2(new_n627), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n462), .A2(new_n465), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n929), .B(KEYINPUT61), .C1(new_n931), .C2(new_n928), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n928), .A2(new_n931), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n888), .A2(new_n927), .ZN(new_n935));
  INV_X1    g749(.A(new_n627), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n899), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n933), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n932), .A2(new_n938), .ZN(G66));
  INV_X1    g753(.A(new_n367), .ZN(new_n940));
  OAI21_X1  g754(.A(G953), .B1(new_n940), .B2(new_n322), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n819), .B2(new_n259), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n892), .B1(G898), .B2(new_n260), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G69));
  AND3_X1   g758(.A1(new_n689), .A2(new_n480), .A3(new_n721), .ZN(new_n945));
  OAI22_X1  g759(.A1(new_n763), .A2(new_n764), .B1(new_n745), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n778), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n806), .A2(new_n706), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n946), .A2(new_n773), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n260), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n387), .A2(new_n391), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n517), .B(KEYINPUT125), .Z(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n637), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n948), .A2(new_n662), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n725), .B(new_n647), .C1(new_n702), .C2(new_n782), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n957), .A2(new_n765), .A3(new_n773), .A4(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n953), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n260), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT126), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(G227), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n259), .B1(new_n963), .B2(new_n636), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n962), .B(new_n964), .ZN(G72));
  XNOR2_X1  g779(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n966));
  NAND2_X1  g780(.A1(G472), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n959), .B2(new_n786), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n655), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n968), .B1(new_n949), .B2(new_n786), .ZN(new_n971));
  INV_X1    g785(.A(new_n419), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n898), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n828), .A2(new_n972), .A3(new_n655), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n968), .B2(new_n975), .ZN(G57));
endmodule


