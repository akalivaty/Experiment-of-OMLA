//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G146), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n191), .B1(KEYINPUT0), .B2(G128), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT0), .B(G128), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI22_X1  g011(.A1(KEYINPUT64), .A2(new_n196), .B1(new_n197), .B2(G137), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT11), .A4(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(KEYINPUT64), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n197), .A2(G137), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n198), .A2(new_n201), .A3(new_n202), .A4(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G131), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(G131), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n195), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n211), .A2(new_n188), .A3(new_n190), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n187), .B(G146), .C1(new_n210), .C2(KEYINPUT1), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n189), .A3(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n211), .A2(new_n188), .A3(new_n190), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n217), .A2(KEYINPUT66), .A3(new_n213), .A4(new_n214), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n200), .A2(G134), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(new_n203), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n204), .B2(G131), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n208), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n226), .A2(KEYINPUT73), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT2), .B(G113), .Z(new_n228));
  XNOR2_X1  g042(.A(G116), .B(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g046(.A1(new_n228), .A2(new_n229), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n232), .B(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n226), .B2(KEYINPUT73), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n227), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT28), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n239));
  INV_X1    g053(.A(G237), .ZN(new_n240));
  INV_X1    g054(.A(G953), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(G210), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n239), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G101), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT71), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n212), .A2(new_n215), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n224), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n234), .B1(new_n208), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT72), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n234), .B(new_n251), .C1(new_n208), .C2(new_n248), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n216), .A2(new_n218), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT67), .B1(new_n254), .B2(new_n224), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n225), .A2(new_n219), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n232), .B(new_n233), .Z(new_n260));
  XNOR2_X1  g074(.A(new_n204), .B(G131), .ZN(new_n261));
  INV_X1    g075(.A(new_n195), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n258), .A2(new_n259), .A3(new_n260), .A4(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n225), .A2(new_n219), .A3(new_n256), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n256), .B1(new_n225), .B2(new_n219), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n260), .B(new_n263), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT68), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n253), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n238), .B(new_n246), .C1(new_n269), .C2(new_n237), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n263), .B(new_n272), .C1(new_n247), .C2(new_n224), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n208), .B1(new_n255), .B2(new_n257), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n273), .B1(new_n274), .B2(new_n272), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n234), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n268), .A2(new_n264), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n245), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n270), .A2(new_n271), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT74), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n274), .A2(new_n260), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(new_n264), .B2(new_n268), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n238), .B1(new_n285), .B2(new_n237), .ZN(new_n286));
  OR3_X1    g100(.A1(new_n286), .A2(new_n271), .A3(new_n279), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n270), .A2(new_n288), .A3(new_n271), .A4(new_n280), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n282), .A2(new_n283), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G472), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n276), .A2(new_n277), .A3(new_n245), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT31), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT70), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n276), .A2(new_n277), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT31), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n245), .ZN(new_n299));
  INV_X1    g113(.A(new_n246), .ZN(new_n300));
  INV_X1    g114(.A(new_n253), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n237), .B1(new_n277), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT28), .B1(new_n227), .B2(new_n235), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n295), .A2(new_n296), .A3(new_n299), .A4(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT32), .B1(new_n305), .B2(new_n306), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT75), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n306), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT32), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n311), .A2(KEYINPUT75), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n291), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G104), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G107), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n317));
  INV_X1    g131(.A(G107), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(G104), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT81), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT82), .B(G107), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT83), .ZN(new_n322));
  NOR4_X1   g136(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT3), .A4(new_n315), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(KEYINPUT82), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G107), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n315), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT83), .B1(new_n327), .B2(new_n317), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n316), .B(new_n320), .C1(new_n323), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G101), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n325), .A2(G107), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n318), .A2(KEYINPUT82), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n317), .B(G104), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n322), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n327), .A2(KEYINPUT83), .A3(new_n317), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G101), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n336), .A2(new_n337), .A3(new_n316), .A4(new_n320), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n330), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n329), .A2(new_n340), .A3(G101), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n341), .A3(new_n262), .ZN(new_n342));
  INV_X1    g156(.A(new_n261), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n318), .A2(G104), .ZN(new_n344));
  INV_X1    g158(.A(new_n321), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(G104), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G101), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n217), .B(KEYINPUT84), .ZN(new_n348));
  INV_X1    g162(.A(new_n215), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n338), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n338), .A2(KEYINPUT10), .A3(new_n347), .A4(new_n219), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n342), .A2(new_n343), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G110), .B(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n241), .A2(G227), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n338), .A2(new_n347), .A3(new_n350), .ZN(new_n362));
  INV_X1    g176(.A(new_n247), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n338), .B2(new_n347), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n261), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT12), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n355), .A2(KEYINPUT85), .A3(new_n358), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n361), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n342), .A2(new_n353), .A3(new_n354), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n261), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n355), .ZN(new_n372));
  INV_X1    g186(.A(new_n358), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G469), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(G469), .A2(G902), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n365), .B(KEYINPUT12), .ZN(new_n379));
  INV_X1    g193(.A(new_n355), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n373), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n371), .A2(new_n355), .A3(new_n358), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(G469), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G221), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT9), .B(G234), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n385), .B1(new_n387), .B2(new_n283), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G125), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n392), .A2(KEYINPUT16), .A3(G140), .ZN(new_n393));
  XNOR2_X1  g207(.A(G125), .B(G140), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(KEYINPUT16), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n189), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n210), .A2(G119), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(KEYINPUT23), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n210), .A2(G119), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G110), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n400), .A2(new_n398), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT24), .B(G110), .Z(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n397), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G110), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n407), .A3(new_n400), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT76), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n408), .A2(new_n409), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n403), .A2(new_n404), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n395), .A2(G146), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n394), .A2(new_n189), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n406), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT77), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT77), .B(new_n406), .C1(new_n413), .C2(new_n416), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT22), .B(G137), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n241), .A2(G221), .A3(G234), .ZN(new_n422));
  XOR2_X1   g236(.A(new_n421), .B(new_n422), .Z(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n417), .A2(new_n418), .A3(new_n423), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G217), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(G234), .B2(new_n283), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n283), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT78), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT79), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT25), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n427), .B2(new_n283), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n427), .A2(new_n436), .A3(new_n283), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n429), .A3(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n435), .A2(KEYINPUT80), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT80), .B1(new_n435), .B2(new_n440), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G128), .B(G143), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT13), .ZN(new_n446));
  OR3_X1    g260(.A1(new_n210), .A2(KEYINPUT13), .A3(G143), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(G134), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n197), .ZN(new_n449));
  XNOR2_X1  g263(.A(G116), .B(G122), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n345), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(G116), .B(G122), .Z(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n321), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n448), .B(new_n449), .C1(new_n451), .C2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n445), .B(new_n197), .ZN(new_n455));
  INV_X1    g269(.A(new_n453), .ZN(new_n456));
  INV_X1    g270(.A(G116), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(KEYINPUT14), .A3(G122), .ZN(new_n458));
  OAI211_X1 g272(.A(G107), .B(new_n458), .C1(new_n452), .C2(KEYINPUT14), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n386), .A2(new_n428), .A3(G953), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n454), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n461), .B1(new_n454), .B2(new_n460), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G902), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT92), .ZN(new_n466));
  INV_X1    g280(.A(G478), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT91), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n466), .A2(new_n472), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT93), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G952), .ZN(new_n481));
  AOI211_X1 g295(.A(G953), .B(new_n481), .C1(G234), .C2(G237), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n283), .B(new_n241), .C1(G234), .C2(G237), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT21), .B(G898), .Z(new_n486));
  OAI21_X1  g300(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(G475), .A2(G902), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n489), .B(KEYINPUT90), .Z(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n240), .A2(new_n241), .A3(G214), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(G143), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT18), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n493), .B1(new_n494), .B2(new_n220), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n394), .B(new_n189), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n492), .B(new_n187), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G131), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n495), .B(new_n496), .C1(new_n494), .C2(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n394), .B(KEYINPUT19), .Z(new_n500));
  OAI21_X1  g314(.A(new_n414), .B1(new_n500), .B2(G146), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n493), .A2(new_n220), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G113), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n315), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n497), .A2(KEYINPUT17), .A3(G131), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n498), .A2(new_n502), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n396), .B(new_n509), .C1(new_n510), .C2(KEYINPUT17), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n506), .A3(new_n499), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(KEYINPUT89), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT89), .B1(new_n508), .B2(new_n512), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n491), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT20), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n490), .A2(KEYINPUT20), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n508), .B2(new_n512), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n511), .A2(new_n499), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n507), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n512), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n283), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n517), .A2(new_n521), .B1(G475), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n480), .A2(new_n488), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G214), .B1(G237), .B2(G902), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n339), .A2(new_n341), .A3(new_n234), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n457), .A2(KEYINPUT5), .A3(G119), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(new_n229), .B2(KEYINPUT5), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n533), .A2(G113), .B1(new_n229), .B2(new_n228), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n338), .A2(new_n347), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(G110), .B(G122), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n537), .B(KEYINPUT86), .Z(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n538), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n531), .A2(new_n540), .A3(new_n535), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(KEYINPUT6), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n195), .A2(G125), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(G125), .B2(new_n363), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n241), .A2(G224), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n545), .B(KEYINPUT87), .Z(new_n546));
  XNOR2_X1  g360(.A(new_n544), .B(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n536), .A2(new_n548), .A3(new_n538), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n542), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT7), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n543), .B2(KEYINPUT88), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n553), .B(new_n544), .Z(new_n554));
  NAND2_X1  g368(.A1(new_n338), .A2(new_n347), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(new_n534), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n538), .B(KEYINPUT8), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n541), .B(new_n554), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n550), .A2(new_n283), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G210), .B1(G237), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n550), .A2(new_n283), .A3(new_n560), .A4(new_n558), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n530), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n528), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n314), .A2(new_n391), .A3(new_n444), .A4(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G101), .ZN(G3));
  AND2_X1   g381(.A1(new_n305), .A2(new_n283), .ZN(new_n568));
  INV_X1    g382(.A(G472), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n311), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n443), .A2(new_n570), .A3(new_n390), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT94), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n562), .A2(new_n573), .A3(new_n563), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n559), .A2(KEYINPUT95), .A3(new_n561), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n574), .A2(new_n529), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT33), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n464), .A2(new_n578), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT33), .ZN(new_n580));
  OAI211_X1 g394(.A(G478), .B(new_n283), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n465), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n582), .A2(KEYINPUT96), .A3(new_n467), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT96), .B1(new_n582), .B2(new_n467), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n526), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n487), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n577), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT34), .B(G104), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  NAND2_X1  g406(.A1(new_n525), .A2(G475), .ZN(new_n593));
  INV_X1    g407(.A(new_n515), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n513), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n517), .B1(new_n596), .B2(new_n519), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n480), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n598), .A2(new_n487), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n577), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT35), .B(G107), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G9));
  INV_X1    g416(.A(new_n570), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n604));
  AOI211_X1 g418(.A(KEYINPUT25), .B(G902), .C1(new_n425), .C2(new_n426), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n437), .A2(new_n605), .A3(new_n430), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n424), .A2(KEYINPUT36), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n417), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n432), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n604), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n440), .A2(KEYINPUT97), .A3(new_n609), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n603), .A2(new_n565), .A3(new_n391), .A4(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT37), .B(G110), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G12));
  XNOR2_X1  g430(.A(KEYINPUT98), .B(G900), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n483), .B1(new_n485), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n598), .A2(new_n618), .ZN(new_n619));
  AND4_X1   g433(.A1(new_n529), .A2(new_n613), .A3(new_n575), .A4(new_n574), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n314), .A2(new_n391), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n311), .A2(new_n312), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n306), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(KEYINPUT75), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n311), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n309), .A3(KEYINPUT32), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n390), .B1(new_n629), .B2(new_n291), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n630), .A2(KEYINPUT99), .A3(new_n619), .A4(new_n620), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT100), .B(G128), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G30));
  XNOR2_X1  g448(.A(new_n618), .B(KEYINPUT39), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n391), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(KEYINPUT40), .Z(new_n637));
  NOR2_X1   g451(.A1(new_n285), .A2(new_n246), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n638), .A2(KEYINPUT101), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n292), .B1(new_n638), .B2(KEYINPUT101), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n283), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(G472), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n629), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n606), .A2(new_n610), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n480), .A2(new_n529), .A3(new_n527), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n562), .A2(new_n563), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT38), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n637), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G143), .ZN(G45));
  NAND2_X1  g466(.A1(new_n587), .A2(new_n618), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n314), .A2(new_n391), .A3(new_n620), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G146), .ZN(G48));
  NAND2_X1  g470(.A1(new_n369), .A2(new_n374), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n283), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(G469), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n375), .B2(new_n376), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n658), .A2(new_n660), .A3(G469), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n388), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n664), .A2(new_n576), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n665), .A2(new_n314), .A3(new_n444), .A4(new_n589), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT41), .B(G113), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G15));
  NAND4_X1  g482(.A1(new_n665), .A2(new_n314), .A3(new_n444), .A4(new_n599), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT103), .B(G116), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G18));
  NAND4_X1  g485(.A1(new_n665), .A2(new_n314), .A3(new_n528), .A4(new_n613), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G119), .ZN(G21));
  NAND2_X1  g487(.A1(new_n574), .A2(new_n575), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n674), .A2(new_n488), .A3(new_n647), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n569), .B1(new_n305), .B2(new_n283), .ZN(new_n676));
  INV_X1    g490(.A(new_n306), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n299), .A2(new_n293), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n286), .A2(new_n300), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n435), .A2(new_n440), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n676), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n675), .A2(new_n664), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G122), .ZN(G24));
  OR3_X1    g498(.A1(new_n676), .A2(new_n680), .A3(new_n645), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n653), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n665), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G125), .ZN(G27));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n625), .A2(KEYINPUT104), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n689), .B1(new_n625), .B2(KEYINPUT104), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n624), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n692), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n308), .A3(new_n690), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n695), .A3(new_n291), .ZN(new_n696));
  INV_X1    g510(.A(new_n681), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n649), .A2(new_n530), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n390), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n696), .A2(new_n697), .A3(new_n654), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT42), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n290), .A2(G472), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n626), .B2(new_n628), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n443), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n653), .A2(KEYINPUT42), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n700), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n220), .ZN(G33));
  NAND3_X1  g523(.A1(new_n705), .A2(new_n619), .A3(new_n700), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G134), .ZN(G36));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n358), .B1(new_n367), .B2(new_n355), .ZN(new_n713));
  INV_X1    g527(.A(new_n382), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n381), .A2(KEYINPUT45), .A3(new_n382), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(G469), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT46), .B1(new_n717), .B2(new_n378), .ZN(new_n718));
  INV_X1    g532(.A(new_n377), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n717), .A2(KEYINPUT46), .A3(new_n378), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n722), .A2(new_n389), .A3(new_n635), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT20), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n595), .B2(new_n491), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n585), .B(new_n593), .C1(new_n725), .C2(new_n520), .ZN(new_n726));
  OAI211_X1 g540(.A(KEYINPUT106), .B(new_n593), .C1(new_n725), .C2(new_n520), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n526), .B(new_n585), .C1(KEYINPUT106), .C2(KEYINPUT43), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n731), .B(new_n646), .C1(new_n627), .C2(new_n676), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n735), .B(new_n698), .C1(new_n732), .C2(new_n733), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n570), .A2(KEYINPUT44), .A3(new_n646), .A4(new_n731), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n735), .B1(new_n738), .B2(new_n698), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n723), .B(new_n734), .C1(new_n737), .C2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G137), .ZN(G39));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n742));
  INV_X1    g556(.A(new_n721), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n743), .A2(new_n718), .A3(new_n719), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n742), .B1(new_n744), .B2(new_n388), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n722), .A2(KEYINPUT47), .A3(new_n389), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n441), .A2(new_n442), .A3(new_n653), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n629), .A2(new_n748), .A3(new_n291), .A4(new_n698), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n704), .A2(KEYINPUT108), .A3(new_n698), .A4(new_n748), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n747), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G140), .ZN(G42));
  NOR2_X1   g568(.A1(new_n527), .A2(new_n476), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n587), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n571), .A2(new_n564), .A3(new_n487), .A4(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n566), .A3(new_n614), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n669), .A2(new_n672), .ZN(new_n760));
  INV_X1    g574(.A(new_n683), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n664), .A2(new_n576), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n704), .A2(new_n762), .A3(new_n443), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n761), .B1(new_n763), .B2(new_n589), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n760), .A2(new_n764), .A3(KEYINPUT109), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n666), .A2(new_n669), .A3(new_n672), .A4(new_n683), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n759), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  AND4_X1   g583(.A1(new_n593), .A2(new_n597), .A3(new_n476), .A4(new_n618), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n314), .A2(new_n613), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n700), .B1(new_n771), .B2(new_n686), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n702), .A2(new_n772), .A3(new_n707), .A4(new_n710), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n655), .A2(new_n687), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n623), .B2(new_n631), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n391), .A2(new_n575), .A3(new_n574), .A4(new_n618), .ZN(new_n777));
  INV_X1    g591(.A(new_n647), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n643), .A3(new_n645), .A4(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n655), .A2(new_n687), .ZN(new_n781));
  AND4_X1   g595(.A1(KEYINPUT52), .A2(new_n632), .A3(new_n781), .A4(new_n779), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n769), .B(new_n774), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n780), .B2(new_n782), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n576), .A2(new_n613), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n704), .A2(new_n390), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT99), .B1(new_n789), .B2(new_n619), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n621), .A2(new_n622), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n781), .B(new_n779), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n776), .A2(KEYINPUT52), .A3(new_n779), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n773), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT110), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n769), .B(new_n796), .C1(new_n797), .C2(KEYINPUT53), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n787), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n483), .B1(new_n729), .B2(new_n730), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n682), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n665), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n759), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n760), .A3(KEYINPUT53), .A4(new_n764), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n783), .A2(new_n784), .B1(new_n796), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n664), .A2(new_n698), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n801), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT116), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(new_n814), .A3(new_n801), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n696), .A2(new_n697), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n816), .A2(KEYINPUT48), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT48), .B1(new_n816), .B2(new_n817), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n685), .B1(new_n813), .B2(new_n815), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n644), .A2(new_n482), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n811), .A2(new_n444), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n527), .A2(new_n585), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n664), .A2(new_n530), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n803), .B1(new_n827), .B2(KEYINPUT113), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(KEYINPUT50), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n650), .B1(new_n827), .B2(KEYINPUT113), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n829), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n833), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n831), .B1(new_n835), .B2(new_n828), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n662), .A2(new_n663), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n388), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n745), .A2(new_n746), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n802), .A2(new_n699), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n826), .A2(KEYINPUT51), .A3(new_n837), .A4(new_n842), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n481), .B(G953), .C1(new_n824), .C2(new_n587), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n820), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n837), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n747), .A2(KEYINPUT112), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT112), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n745), .A2(new_n746), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n839), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n841), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT115), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n847), .A2(new_n826), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(KEYINPUT117), .A3(new_n855), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n845), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n800), .A2(new_n804), .A3(new_n810), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n481), .A2(new_n241), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n809), .B1(new_n787), .B2(new_n798), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT53), .B1(new_n796), .B2(new_n769), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n773), .B(new_n806), .C1(new_n794), .C2(new_n795), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n866), .A2(KEYINPUT54), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT118), .A3(new_n804), .A4(new_n860), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n863), .A2(new_n864), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n838), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n697), .B1(new_n872), .B2(KEYINPUT49), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(KEYINPUT49), .B2(new_n872), .ZN(new_n874));
  INV_X1    g688(.A(new_n650), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n726), .A2(new_n388), .A3(new_n530), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n874), .A2(new_n875), .A3(new_n644), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n871), .A2(new_n877), .ZN(G75));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n879));
  OAI211_X1 g693(.A(G210), .B(G902), .C1(new_n866), .C2(new_n867), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(KEYINPUT120), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(KEYINPUT119), .A3(new_n881), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n542), .A2(new_n549), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n547), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT55), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n879), .A2(new_n882), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n882), .A2(new_n879), .A3(new_n886), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n241), .A2(G952), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G51));
  NOR2_X1   g704(.A1(new_n808), .A2(new_n809), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n868), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n378), .B(KEYINPUT57), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n657), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n808), .A2(new_n283), .A3(new_n717), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(G54));
  NOR2_X1   g710(.A1(new_n808), .A2(new_n283), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n898), .A2(new_n596), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n596), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n889), .ZN(G60));
  NOR2_X1   g715(.A1(new_n579), .A2(new_n580), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT121), .Z(new_n903));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT59), .Z(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n869), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n889), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n892), .A2(new_n903), .A3(new_n905), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(G63));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n911));
  NAND2_X1  g725(.A1(G217), .A2(G902), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT60), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT122), .B1(new_n808), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n427), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n916));
  INV_X1    g730(.A(new_n913), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n916), .B(new_n917), .C1(new_n866), .C2(new_n867), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n907), .ZN(new_n920));
  INV_X1    g734(.A(new_n608), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n914), .B2(new_n918), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n911), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n922), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n924), .A2(KEYINPUT61), .A3(new_n907), .A4(new_n919), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(G66));
  AOI21_X1  g740(.A(new_n241), .B1(new_n486), .B2(G224), .ZN(new_n927));
  INV_X1    g741(.A(new_n769), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n241), .ZN(new_n929));
  INV_X1    g743(.A(G898), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n884), .B1(new_n930), .B2(G953), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n929), .B(new_n931), .ZN(G69));
  AOI21_X1  g746(.A(new_n241), .B1(G227), .B2(G900), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n753), .A2(new_n740), .A3(new_n710), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n708), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n632), .A2(new_n781), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT123), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n776), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n674), .A2(new_n647), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n696), .A2(new_n723), .A3(new_n697), .A4(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n935), .A2(new_n937), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n632), .A2(new_n938), .A3(new_n781), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n938), .B1(new_n632), .B2(new_n781), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n946), .A2(new_n947), .A3(new_n941), .A4(new_n935), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n943), .A2(new_n241), .A3(new_n948), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n275), .B(new_n500), .Z(new_n950));
  NAND2_X1  g764(.A1(G900), .A2(G953), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n933), .B1(new_n952), .B2(KEYINPUT125), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n705), .B(new_n698), .C1(KEYINPUT124), .C2(new_n756), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n636), .B(new_n954), .C1(KEYINPUT124), .C2(new_n756), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n937), .A2(new_n651), .A3(new_n939), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n937), .A2(new_n939), .A3(KEYINPUT62), .A4(new_n651), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n753), .A2(new_n740), .ZN(new_n961));
  AOI21_X1  g775(.A(G953), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n952), .B1(new_n962), .B2(new_n950), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n953), .B(new_n963), .Z(G72));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT63), .Z(new_n966));
  NAND2_X1  g780(.A1(new_n280), .A2(new_n292), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n799), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n960), .A2(new_n769), .A3(new_n961), .ZN(new_n969));
  AOI211_X1 g783(.A(new_n279), .B(new_n297), .C1(new_n969), .C2(new_n966), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n943), .A2(new_n769), .A3(new_n948), .ZN(new_n972));
  AOI211_X1 g786(.A(new_n245), .B(new_n278), .C1(new_n972), .C2(new_n966), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n973), .B2(new_n889), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n966), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(new_n279), .A3(new_n297), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(KEYINPUT127), .A3(new_n907), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n968), .B(new_n970), .C1(new_n974), .C2(new_n977), .ZN(G57));
endmodule


