

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U545 ( .A(n729), .ZN(n713) );
  OR2_X1 U546 ( .A1(n751), .A2(KEYINPUT33), .ZN(n755) );
  OR2_X1 U547 ( .A1(n753), .A2(n764), .ZN(n513) );
  XOR2_X1 U548 ( .A(n700), .B(KEYINPUT93), .Z(n514) );
  OR2_X1 U549 ( .A1(n697), .A2(n847), .ZN(n698) );
  NOR2_X1 U550 ( .A1(G299), .A2(n707), .ZN(n705) );
  NAND2_X1 U551 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U552 ( .A(n746), .B(KEYINPUT98), .ZN(n759) );
  AND2_X1 U553 ( .A1(n971), .A2(n513), .ZN(n754) );
  AND2_X1 U554 ( .A1(n688), .A2(G40), .ZN(n769) );
  NAND2_X1 U555 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U556 ( .A(n598), .B(n597), .ZN(n959) );
  XOR2_X1 U557 ( .A(KEYINPUT0), .B(G543), .Z(n635) );
  XNOR2_X1 U558 ( .A(n525), .B(KEYINPUT72), .ZN(G299) );
  NOR2_X1 U559 ( .A1(G651), .A2(n635), .ZN(n515) );
  XNOR2_X2 U560 ( .A(KEYINPUT64), .B(n515), .ZN(n650) );
  NAND2_X1 U561 ( .A1(n650), .A2(G53), .ZN(n524) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n646) );
  NAND2_X1 U563 ( .A1(G91), .A2(n646), .ZN(n517) );
  INV_X1 U564 ( .A(G651), .ZN(n518) );
  NOR2_X1 U565 ( .A1(n635), .A2(n518), .ZN(n644) );
  NAND2_X1 U566 ( .A1(G78), .A2(n644), .ZN(n516) );
  NAND2_X1 U567 ( .A1(n517), .A2(n516), .ZN(n522) );
  NOR2_X1 U568 ( .A1(G543), .A2(n518), .ZN(n519) );
  XOR2_X2 U569 ( .A(KEYINPUT1), .B(n519), .Z(n647) );
  NAND2_X1 U570 ( .A1(G65), .A2(n647), .ZN(n520) );
  XNOR2_X1 U571 ( .A(KEYINPUT71), .B(n520), .ZN(n521) );
  NOR2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U574 ( .A1(G62), .A2(n647), .ZN(n527) );
  NAND2_X1 U575 ( .A1(G50), .A2(n650), .ZN(n526) );
  NAND2_X1 U576 ( .A1(n527), .A2(n526), .ZN(n531) );
  NAND2_X1 U577 ( .A1(G88), .A2(n646), .ZN(n529) );
  NAND2_X1 U578 ( .A1(G75), .A2(n644), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U581 ( .A(n532), .B(KEYINPUT82), .ZN(G166) );
  INV_X1 U582 ( .A(G166), .ZN(G303) );
  NAND2_X1 U583 ( .A1(n647), .A2(G64), .ZN(n533) );
  XNOR2_X1 U584 ( .A(n533), .B(KEYINPUT68), .ZN(n535) );
  NAND2_X1 U585 ( .A1(G52), .A2(n650), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U587 ( .A(KEYINPUT69), .B(n536), .Z(n542) );
  NAND2_X1 U588 ( .A1(n646), .A2(G90), .ZN(n537) );
  XNOR2_X1 U589 ( .A(n537), .B(KEYINPUT70), .ZN(n539) );
  NAND2_X1 U590 ( .A1(G77), .A2(n644), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U592 ( .A(KEYINPUT9), .B(n540), .Z(n541) );
  NOR2_X1 U593 ( .A1(n542), .A2(n541), .ZN(G171) );
  XNOR2_X1 U594 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n544) );
  NOR2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n543) );
  XNOR2_X2 U596 ( .A(n544), .B(n543), .ZN(n878) );
  NAND2_X1 U597 ( .A1(G137), .A2(n878), .ZN(n546) );
  INV_X1 U598 ( .A(G2105), .ZN(n555) );
  NOR2_X2 U599 ( .A1(G2104), .A2(n555), .ZN(n882) );
  NAND2_X1 U600 ( .A1(G125), .A2(n882), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n553) );
  INV_X1 U602 ( .A(G2104), .ZN(n554) );
  NOR2_X4 U603 ( .A1(G2105), .A2(n554), .ZN(n877) );
  NAND2_X1 U604 ( .A1(G101), .A2(n877), .ZN(n547) );
  NAND2_X1 U605 ( .A1(KEYINPUT23), .A2(n547), .ZN(n551) );
  INV_X1 U606 ( .A(KEYINPUT23), .ZN(n549) );
  INV_X1 U607 ( .A(n547), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n558) );
  NOR2_X2 U611 ( .A1(n555), .A2(n554), .ZN(n881) );
  NAND2_X1 U612 ( .A1(G113), .A2(n881), .ZN(n556) );
  XNOR2_X1 U613 ( .A(n556), .B(KEYINPUT66), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U615 ( .A(n559), .B(KEYINPUT65), .ZN(n688) );
  BUF_X1 U616 ( .A(n688), .Z(G160) );
  XNOR2_X1 U617 ( .A(G2451), .B(G2427), .ZN(n569) );
  XOR2_X1 U618 ( .A(G2430), .B(G2443), .Z(n561) );
  XNOR2_X1 U619 ( .A(G2435), .B(G2438), .ZN(n560) );
  XNOR2_X1 U620 ( .A(n561), .B(n560), .ZN(n565) );
  XOR2_X1 U621 ( .A(G2454), .B(KEYINPUT105), .Z(n563) );
  XNOR2_X1 U622 ( .A(G1348), .B(G1341), .ZN(n562) );
  XNOR2_X1 U623 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U624 ( .A(n565), .B(n564), .Z(n567) );
  XNOR2_X1 U625 ( .A(G2446), .B(KEYINPUT106), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U627 ( .A(n569), .B(n568), .ZN(n570) );
  AND2_X1 U628 ( .A1(n570), .A2(G14), .ZN(G401) );
  AND2_X1 U629 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U630 ( .A1(G111), .A2(n881), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G135), .A2(n878), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n882), .A2(G123), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT18), .B(n573), .Z(n574) );
  NOR2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n877), .A2(G99), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n926) );
  XNOR2_X1 U638 ( .A(G2096), .B(n926), .ZN(n578) );
  OR2_X1 U639 ( .A1(G2100), .A2(n578), .ZN(G156) );
  INV_X1 U640 ( .A(G57), .ZN(G237) );
  INV_X1 U641 ( .A(G132), .ZN(G219) );
  NAND2_X1 U642 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n579), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U644 ( .A(G223), .ZN(n822) );
  NAND2_X1 U645 ( .A1(n822), .A2(G567), .ZN(n580) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(n580), .Z(G234) );
  NAND2_X1 U647 ( .A1(n646), .A2(G81), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT12), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G68), .A2(n644), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n585) );
  XOR2_X1 U651 ( .A(KEYINPUT74), .B(KEYINPUT13), .Z(n584) );
  XNOR2_X1 U652 ( .A(n585), .B(n584), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n647), .A2(G56), .ZN(n586) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(n586), .Z(n587) );
  NOR2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U656 ( .A1(G43), .A2(n650), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n953) );
  INV_X1 U658 ( .A(G860), .ZN(n614) );
  OR2_X1 U659 ( .A1(n953), .A2(n614), .ZN(G153) );
  INV_X1 U660 ( .A(G171), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U662 ( .A1(G92), .A2(n646), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G79), .A2(n644), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U665 ( .A1(G66), .A2(n647), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G54), .A2(n650), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n598) );
  XNOR2_X1 U669 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n597) );
  INV_X1 U670 ( .A(n959), .ZN(n847) );
  INV_X1 U671 ( .A(G868), .ZN(n664) );
  NAND2_X1 U672 ( .A1(n847), .A2(n664), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U674 ( .A1(G63), .A2(n647), .ZN(n602) );
  NAND2_X1 U675 ( .A1(G51), .A2(n650), .ZN(n601) );
  NAND2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U677 ( .A(KEYINPUT6), .B(n603), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n646), .A2(G89), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n604), .B(KEYINPUT4), .ZN(n606) );
  NAND2_X1 U680 ( .A1(G76), .A2(n644), .ZN(n605) );
  NAND2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U682 ( .A(n607), .B(KEYINPUT5), .Z(n608) );
  NOR2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U684 ( .A(KEYINPUT76), .B(n610), .Z(n611) );
  XNOR2_X1 U685 ( .A(KEYINPUT7), .B(n611), .ZN(G168) );
  XOR2_X1 U686 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U687 ( .A1(G868), .A2(G286), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G299), .A2(n664), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U690 ( .A1(n614), .A2(G559), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n615), .A2(n959), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U693 ( .A1(n847), .A2(n664), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n617), .B(KEYINPUT77), .ZN(n618) );
  NOR2_X1 U695 ( .A1(G559), .A2(n618), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n619), .B(KEYINPUT78), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n953), .A2(G868), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(G282) );
  NAND2_X1 U699 ( .A1(G559), .A2(n959), .ZN(n622) );
  XOR2_X1 U700 ( .A(n953), .B(n622), .Z(n661) );
  XNOR2_X1 U701 ( .A(KEYINPUT79), .B(n661), .ZN(n623) );
  NOR2_X1 U702 ( .A1(G860), .A2(n623), .ZN(n631) );
  NAND2_X1 U703 ( .A1(G93), .A2(n646), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G80), .A2(n644), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n650), .A2(G55), .ZN(n626) );
  XOR2_X1 U707 ( .A(KEYINPUT80), .B(n626), .Z(n627) );
  NOR2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n647), .A2(G67), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n663) );
  XOR2_X1 U711 ( .A(n631), .B(n663), .Z(G145) );
  NAND2_X1 U712 ( .A1(G651), .A2(G74), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G49), .A2(n650), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U715 ( .A1(n647), .A2(n634), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n635), .A2(G87), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(G288) );
  AND2_X1 U718 ( .A1(n647), .A2(G60), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G85), .A2(n646), .ZN(n639) );
  NAND2_X1 U720 ( .A1(G72), .A2(n644), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G47), .A2(n650), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(G290) );
  NAND2_X1 U725 ( .A1(G73), .A2(n644), .ZN(n645) );
  XNOR2_X1 U726 ( .A(n645), .B(KEYINPUT2), .ZN(n655) );
  NAND2_X1 U727 ( .A1(G86), .A2(n646), .ZN(n649) );
  NAND2_X1 U728 ( .A1(G61), .A2(n647), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U730 ( .A1(G48), .A2(n650), .ZN(n651) );
  XNOR2_X1 U731 ( .A(KEYINPUT81), .B(n651), .ZN(n652) );
  NOR2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(G305) );
  XNOR2_X1 U734 ( .A(G303), .B(G299), .ZN(n660) );
  XNOR2_X1 U735 ( .A(KEYINPUT19), .B(G288), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(n663), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n657), .B(G290), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n658), .B(G305), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n660), .B(n659), .ZN(n850) );
  XNOR2_X1 U740 ( .A(n661), .B(n850), .ZN(n662) );
  NAND2_X1 U741 ( .A1(n662), .A2(G868), .ZN(n666) );
  NAND2_X1 U742 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U743 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U748 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U750 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  NOR2_X1 U751 ( .A1(G219), .A2(G220), .ZN(n671) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U753 ( .A1(G218), .A2(n672), .ZN(n673) );
  XOR2_X1 U754 ( .A(KEYINPUT83), .B(n673), .Z(n674) );
  NAND2_X1 U755 ( .A1(G96), .A2(n674), .ZN(n827) );
  NAND2_X1 U756 ( .A1(G2106), .A2(n827), .ZN(n678) );
  NAND2_X1 U757 ( .A1(G69), .A2(G120), .ZN(n675) );
  NOR2_X1 U758 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U759 ( .A1(G108), .A2(n676), .ZN(n828) );
  NAND2_X1 U760 ( .A1(G567), .A2(n828), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U762 ( .A(KEYINPUT84), .B(n679), .Z(G319) );
  INV_X1 U763 ( .A(G319), .ZN(n898) );
  NAND2_X1 U764 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U765 ( .A1(n898), .A2(n680), .ZN(n824) );
  NAND2_X1 U766 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U767 ( .A1(n881), .A2(G114), .ZN(n683) );
  NAND2_X1 U768 ( .A1(G102), .A2(n877), .ZN(n681) );
  XOR2_X1 U769 ( .A(KEYINPUT85), .B(n681), .Z(n682) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n687) );
  NAND2_X1 U771 ( .A1(G138), .A2(n878), .ZN(n685) );
  NAND2_X1 U772 ( .A1(G126), .A2(n882), .ZN(n684) );
  NAND2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U774 ( .A1(n687), .A2(n686), .ZN(G164) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n771) );
  NAND2_X2 U776 ( .A1(n769), .A2(n771), .ZN(n729) );
  NAND2_X1 U777 ( .A1(G8), .A2(n729), .ZN(n764) );
  XNOR2_X1 U778 ( .A(G1996), .B(KEYINPUT92), .ZN(n906) );
  NAND2_X1 U779 ( .A1(n713), .A2(n906), .ZN(n689) );
  XNOR2_X1 U780 ( .A(n689), .B(KEYINPUT26), .ZN(n692) );
  AND2_X1 U781 ( .A1(n729), .A2(G1341), .ZN(n690) );
  NOR2_X1 U782 ( .A1(n690), .A2(n953), .ZN(n691) );
  AND2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n696) );
  NOR2_X1 U784 ( .A1(n713), .A2(G1348), .ZN(n694) );
  NOR2_X1 U785 ( .A1(G2067), .A2(n729), .ZN(n693) );
  NOR2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U787 ( .A1(n697), .A2(n847), .ZN(n695) );
  NAND2_X1 U788 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U789 ( .A1(n699), .A2(n698), .ZN(n700) );
  INV_X1 U790 ( .A(KEYINPUT27), .ZN(n702) );
  NAND2_X1 U791 ( .A1(n713), .A2(G2072), .ZN(n701) );
  XNOR2_X1 U792 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U793 ( .A1(G1956), .A2(n729), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n707) );
  XNOR2_X1 U795 ( .A(KEYINPUT94), .B(n705), .ZN(n706) );
  NOR2_X1 U796 ( .A1(n514), .A2(n706), .ZN(n710) );
  NAND2_X1 U797 ( .A1(G299), .A2(n707), .ZN(n708) );
  XOR2_X1 U798 ( .A(KEYINPUT28), .B(n708), .Z(n709) );
  NOR2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U800 ( .A(n711), .B(KEYINPUT29), .ZN(n717) );
  NOR2_X1 U801 ( .A1(n713), .A2(G1961), .ZN(n712) );
  XNOR2_X1 U802 ( .A(n712), .B(KEYINPUT91), .ZN(n715) );
  XNOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .ZN(n903) );
  NAND2_X1 U804 ( .A1(n713), .A2(n903), .ZN(n714) );
  NAND2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n721) );
  NAND2_X1 U806 ( .A1(G171), .A2(n721), .ZN(n716) );
  NAND2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n727) );
  NOR2_X1 U808 ( .A1(G1966), .A2(n764), .ZN(n741) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n729), .ZN(n738) );
  NOR2_X1 U810 ( .A1(n741), .A2(n738), .ZN(n718) );
  NAND2_X1 U811 ( .A1(G8), .A2(n718), .ZN(n719) );
  XNOR2_X1 U812 ( .A(KEYINPUT30), .B(n719), .ZN(n720) );
  NOR2_X1 U813 ( .A1(G168), .A2(n720), .ZN(n724) );
  NOR2_X1 U814 ( .A1(G171), .A2(n721), .ZN(n722) );
  XOR2_X1 U815 ( .A(KEYINPUT95), .B(n722), .Z(n723) );
  NOR2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U817 ( .A(KEYINPUT31), .B(n725), .Z(n726) );
  NAND2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n739) );
  NAND2_X1 U819 ( .A1(n739), .A2(G286), .ZN(n728) );
  XNOR2_X1 U820 ( .A(n728), .B(KEYINPUT96), .ZN(n734) );
  NOR2_X1 U821 ( .A1(G1971), .A2(n764), .ZN(n731) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n729), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U824 ( .A1(n732), .A2(G303), .ZN(n733) );
  NAND2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U826 ( .A1(n735), .A2(G8), .ZN(n737) );
  XOR2_X1 U827 ( .A(KEYINPUT97), .B(KEYINPUT32), .Z(n736) );
  XNOR2_X1 U828 ( .A(n737), .B(n736), .ZN(n745) );
  NAND2_X1 U829 ( .A1(G8), .A2(n738), .ZN(n743) );
  INV_X1 U830 ( .A(n739), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n752) );
  NOR2_X1 U834 ( .A1(G303), .A2(G1971), .ZN(n747) );
  NOR2_X1 U835 ( .A1(n752), .A2(n747), .ZN(n956) );
  NAND2_X1 U836 ( .A1(n759), .A2(n956), .ZN(n749) );
  NAND2_X1 U837 ( .A1(G288), .A2(G1976), .ZN(n748) );
  XOR2_X1 U838 ( .A(KEYINPUT99), .B(n748), .Z(n962) );
  NAND2_X1 U839 ( .A1(n749), .A2(n962), .ZN(n750) );
  NOR2_X1 U840 ( .A1(n764), .A2(n750), .ZN(n751) );
  XOR2_X1 U841 ( .A(G1981), .B(G305), .Z(n971) );
  NAND2_X1 U842 ( .A1(n752), .A2(KEYINPUT33), .ZN(n753) );
  XNOR2_X1 U843 ( .A(n756), .B(KEYINPUT100), .ZN(n768) );
  NOR2_X1 U844 ( .A1(G303), .A2(G2090), .ZN(n757) );
  XOR2_X1 U845 ( .A(KEYINPUT101), .B(n757), .Z(n758) );
  NAND2_X1 U846 ( .A1(G8), .A2(n758), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n761) );
  AND2_X1 U848 ( .A1(n761), .A2(n764), .ZN(n766) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U850 ( .A(n762), .B(KEYINPUT24), .Z(n763) );
  NOR2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n804) );
  INV_X1 U854 ( .A(n769), .ZN(n770) );
  NOR2_X1 U855 ( .A1(n771), .A2(n770), .ZN(n817) );
  NAND2_X1 U856 ( .A1(n877), .A2(G104), .ZN(n772) );
  XNOR2_X1 U857 ( .A(n772), .B(KEYINPUT86), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G140), .A2(n878), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n775), .ZN(n781) );
  NAND2_X1 U861 ( .A1(n882), .A2(G128), .ZN(n776) );
  XOR2_X1 U862 ( .A(KEYINPUT87), .B(n776), .Z(n778) );
  NAND2_X1 U863 ( .A1(n881), .A2(G116), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U865 ( .A(KEYINPUT35), .B(n779), .Z(n780) );
  NOR2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(n782), .ZN(n864) );
  XNOR2_X1 U868 ( .A(KEYINPUT37), .B(G2067), .ZN(n815) );
  NOR2_X1 U869 ( .A1(n864), .A2(n815), .ZN(n942) );
  NAND2_X1 U870 ( .A1(n817), .A2(n942), .ZN(n812) );
  XOR2_X1 U871 ( .A(G1986), .B(G290), .Z(n963) );
  NAND2_X1 U872 ( .A1(G107), .A2(n881), .ZN(n784) );
  NAND2_X1 U873 ( .A1(G131), .A2(n878), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G95), .A2(n877), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G119), .A2(n882), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n787) );
  OR2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n892) );
  NAND2_X1 U879 ( .A1(G1991), .A2(n892), .ZN(n799) );
  NAND2_X1 U880 ( .A1(G105), .A2(n877), .ZN(n789) );
  XNOR2_X1 U881 ( .A(n789), .B(KEYINPUT38), .ZN(n796) );
  NAND2_X1 U882 ( .A1(G117), .A2(n881), .ZN(n791) );
  NAND2_X1 U883 ( .A1(G141), .A2(n878), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n882), .A2(G129), .ZN(n792) );
  XOR2_X1 U886 ( .A(KEYINPUT88), .B(n792), .Z(n793) );
  NOR2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U889 ( .A(KEYINPUT89), .B(n797), .Z(n865) );
  NAND2_X1 U890 ( .A1(G1996), .A2(n865), .ZN(n798) );
  NAND2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U892 ( .A(KEYINPUT90), .B(n800), .Z(n947) );
  NAND2_X1 U893 ( .A1(n963), .A2(n947), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n801), .A2(n817), .ZN(n802) );
  AND2_X1 U895 ( .A1(n812), .A2(n802), .ZN(n803) );
  NAND2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n820) );
  INV_X1 U897 ( .A(n947), .ZN(n807) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U899 ( .A1(G1991), .A2(n892), .ZN(n929) );
  NOR2_X1 U900 ( .A1(n805), .A2(n929), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n809) );
  NOR2_X1 U902 ( .A1(n865), .A2(G1996), .ZN(n808) );
  XNOR2_X1 U903 ( .A(n808), .B(KEYINPUT102), .ZN(n933) );
  NOR2_X1 U904 ( .A1(n809), .A2(n933), .ZN(n810) );
  XOR2_X1 U905 ( .A(KEYINPUT103), .B(n810), .Z(n811) );
  XNOR2_X1 U906 ( .A(KEYINPUT39), .B(n811), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U908 ( .A(n814), .B(KEYINPUT104), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n864), .A2(n815), .ZN(n930) );
  NAND2_X1 U910 ( .A1(n816), .A2(n930), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U913 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U916 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U919 ( .A(KEYINPUT107), .B(n826), .Z(G188) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U926 ( .A(G1991), .B(KEYINPUT41), .ZN(n838) );
  XOR2_X1 U927 ( .A(G1971), .B(G1956), .Z(n830) );
  XNOR2_X1 U928 ( .A(G1996), .B(G1986), .ZN(n829) );
  XNOR2_X1 U929 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U930 ( .A(G1976), .B(G1981), .Z(n832) );
  XNOR2_X1 U931 ( .A(G1966), .B(G1961), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U933 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U934 ( .A(G2474), .B(KEYINPUT108), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(G229) );
  XOR2_X1 U937 ( .A(G2100), .B(G2096), .Z(n840) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2072), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2090), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(G227) );
  XNOR2_X1 U946 ( .A(KEYINPUT112), .B(n847), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n848), .B(n953), .ZN(n849) );
  XNOR2_X1 U948 ( .A(KEYINPUT111), .B(n849), .ZN(n852) );
  XNOR2_X1 U949 ( .A(G286), .B(n850), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n853), .B(G171), .ZN(n854) );
  NOR2_X1 U952 ( .A1(G37), .A2(n854), .ZN(G397) );
  NAND2_X1 U953 ( .A1(G124), .A2(n882), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U955 ( .A1(n881), .A2(G112), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G100), .A2(n877), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G136), .A2(n878), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U960 ( .A1(n861), .A2(n860), .ZN(G162) );
  XNOR2_X1 U961 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n926), .B(KEYINPUT110), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n891) );
  XNOR2_X1 U964 ( .A(G160), .B(n864), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n876) );
  NAND2_X1 U966 ( .A1(G118), .A2(n881), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G130), .A2(n882), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U969 ( .A1(G106), .A2(n877), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G142), .A2(n878), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U972 ( .A(KEYINPUT45), .B(n871), .ZN(n872) );
  XNOR2_X1 U973 ( .A(KEYINPUT109), .B(n872), .ZN(n873) );
  NOR2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U975 ( .A(n876), .B(n875), .Z(n889) );
  NAND2_X1 U976 ( .A1(G103), .A2(n877), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G139), .A2(n878), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U979 ( .A1(G115), .A2(n881), .ZN(n884) );
  NAND2_X1 U980 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n936) );
  XNOR2_X1 U984 ( .A(G164), .B(n936), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n894) );
  XNOR2_X1 U987 ( .A(n892), .B(G162), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U989 ( .A1(G37), .A2(n895), .ZN(G395) );
  NOR2_X1 U990 ( .A1(G229), .A2(G227), .ZN(n896) );
  XNOR2_X1 U991 ( .A(KEYINPUT49), .B(n896), .ZN(n897) );
  NOR2_X1 U992 ( .A1(G401), .A2(n897), .ZN(n900) );
  NOR2_X1 U993 ( .A1(G397), .A2(n898), .ZN(n899) );
  NAND2_X1 U994 ( .A1(n900), .A2(n899), .ZN(n901) );
  NOR2_X1 U995 ( .A1(n901), .A2(G395), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n902), .B(KEYINPUT113), .ZN(G225) );
  INV_X1 U997 ( .A(G225), .ZN(G308) );
  INV_X1 U998 ( .A(G108), .ZN(G238) );
  XOR2_X1 U999 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1009) );
  XNOR2_X1 U1000 ( .A(G2090), .B(G35), .ZN(n918) );
  XOR2_X1 U1001 ( .A(G2067), .B(G26), .Z(n905) );
  XNOR2_X1 U1002 ( .A(n903), .B(G27), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(G32), .B(n906), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n911) );
  XOR2_X1 U1006 ( .A(G2072), .B(G33), .Z(n909) );
  XNOR2_X1 U1007 ( .A(KEYINPUT116), .B(n909), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(KEYINPUT117), .B(n912), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n913), .A2(G28), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(G25), .B(G1991), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(KEYINPUT53), .B(n916), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n919), .B(KEYINPUT118), .ZN(n922) );
  XOR2_X1 U1016 ( .A(G2084), .B(G34), .Z(n920) );
  XNOR2_X1 U1017 ( .A(KEYINPUT54), .B(n920), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(KEYINPUT119), .B(n923), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G29), .A2(n924), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(n925), .B(KEYINPUT55), .ZN(n952) );
  XNOR2_X1 U1022 ( .A(G160), .B(G2084), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n931) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n946) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1028 ( .A(KEYINPUT114), .B(n934), .Z(n935) );
  XNOR2_X1 U1029 ( .A(KEYINPUT51), .B(n935), .ZN(n944) );
  XNOR2_X1 U1030 ( .A(G2072), .B(n936), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(G164), .B(G2078), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1033 ( .A(n939), .B(KEYINPUT50), .Z(n940) );
  XNOR2_X1 U1034 ( .A(KEYINPUT115), .B(n940), .ZN(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n948) );
  NAND2_X1 U1038 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1039 ( .A(KEYINPUT52), .B(n949), .ZN(n950) );
  NAND2_X1 U1040 ( .A1(G29), .A2(n950), .ZN(n951) );
  NAND2_X1 U1041 ( .A1(n952), .A2(n951), .ZN(n1006) );
  XNOR2_X1 U1042 ( .A(G16), .B(KEYINPUT56), .ZN(n978) );
  XNOR2_X1 U1043 ( .A(G1341), .B(KEYINPUT122), .ZN(n954) );
  XNOR2_X1 U1044 ( .A(n954), .B(n953), .ZN(n958) );
  NAND2_X1 U1045 ( .A1(G303), .A2(G1971), .ZN(n955) );
  NAND2_X1 U1046 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1047 ( .A1(n958), .A2(n957), .ZN(n967) );
  XOR2_X1 U1048 ( .A(G299), .B(G1956), .Z(n961) );
  XNOR2_X1 U1049 ( .A(G1348), .B(n959), .ZN(n960) );
  NAND2_X1 U1050 ( .A1(n961), .A2(n960), .ZN(n965) );
  NAND2_X1 U1051 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1052 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1053 ( .A1(n967), .A2(n966), .ZN(n970) );
  XOR2_X1 U1054 ( .A(G1961), .B(G301), .Z(n968) );
  XNOR2_X1 U1055 ( .A(KEYINPUT121), .B(n968), .ZN(n969) );
  NOR2_X1 U1056 ( .A1(n970), .A2(n969), .ZN(n976) );
  XNOR2_X1 U1057 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n974) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G168), .ZN(n972) );
  NAND2_X1 U1059 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1060 ( .A(n974), .B(n973), .ZN(n975) );
  NAND2_X1 U1061 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1062 ( .A1(n978), .A2(n977), .ZN(n1003) );
  XOR2_X1 U1063 ( .A(G1956), .B(G20), .Z(n983) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n980) );
  XNOR2_X1 U1065 ( .A(G6), .B(G1981), .ZN(n979) );
  NOR2_X1 U1066 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1067 ( .A(KEYINPUT124), .B(n981), .ZN(n982) );
  NAND2_X1 U1068 ( .A1(n983), .A2(n982), .ZN(n986) );
  XOR2_X1 U1069 ( .A(KEYINPUT59), .B(G1348), .Z(n984) );
  XNOR2_X1 U1070 ( .A(G4), .B(n984), .ZN(n985) );
  NOR2_X1 U1071 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1072 ( .A(KEYINPUT60), .B(n987), .ZN(n991) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G21), .ZN(n989) );
  XNOR2_X1 U1074 ( .A(G1961), .B(G5), .ZN(n988) );
  NOR2_X1 U1075 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1076 ( .A1(n991), .A2(n990), .ZN(n998) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n993) );
  XNOR2_X1 U1078 ( .A(G23), .B(G1976), .ZN(n992) );
  NOR2_X1 U1079 ( .A1(n993), .A2(n992), .ZN(n995) );
  XOR2_X1 U1080 ( .A(G1986), .B(G24), .Z(n994) );
  NAND2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(KEYINPUT58), .B(n996), .ZN(n997) );
  NOR2_X1 U1083 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(n999), .B(KEYINPUT61), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(G16), .B(KEYINPUT123), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1088 ( .A(KEYINPUT125), .B(n1004), .Z(n1005) );
  NOR2_X1 U1089 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1090 ( .A1(n1007), .A2(G11), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(n1009), .B(n1008), .ZN(G311) );
  XNOR2_X1 U1092 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

