//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961;
  NAND2_X1  g000(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT26), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n205), .B(new_n206), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  AND2_X1   g011(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT28), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g016(.A(KEYINPUT28), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n218));
  AOI211_X1 g017(.A(KEYINPUT66), .B(new_n211), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n218), .ZN(new_n221));
  INV_X1    g020(.A(new_n211), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(KEYINPUT23), .B2(new_n209), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n203), .A2(KEYINPUT65), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G169gat), .ZN(new_n228));
  AOI21_X1  g027(.A(G176gat), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n225), .B1(new_n229), .B2(KEYINPUT23), .ZN(new_n230));
  OR2_X1    g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(KEYINPUT24), .A3(new_n206), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n206), .A2(KEYINPUT24), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT25), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n203), .A2(new_n204), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n210), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(new_n224), .B2(KEYINPUT23), .ZN(new_n240));
  AND4_X1   g039(.A1(new_n232), .A2(new_n238), .A3(new_n233), .A4(new_n240), .ZN(new_n241));
  OAI22_X1  g040(.A1(new_n219), .A2(new_n223), .B1(new_n235), .B2(new_n241), .ZN(new_n242));
  OR2_X1    g041(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G113gat), .ZN(new_n246));
  INV_X1    g045(.A(G113gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G120gat), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT1), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G127gat), .B(G134gat), .ZN(new_n250));
  XOR2_X1   g049(.A(G127gat), .B(G134gat), .Z(new_n251));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n251), .B(new_n252), .C1(KEYINPUT1), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G113gat), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT1), .B1(new_n248), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT67), .B1(new_n257), .B2(new_n250), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n249), .A2(new_n250), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n258), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n247), .B1(new_n243), .B2(new_n244), .ZN(new_n264));
  INV_X1    g063(.A(new_n248), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n263), .B(new_n250), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n260), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n242), .A2(new_n261), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n226), .A2(new_n228), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT23), .A3(new_n204), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n271), .A2(new_n232), .A3(new_n233), .A4(new_n238), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n239), .ZN(new_n273));
  INV_X1    g072(.A(new_n241), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n275), .B(new_n267), .C1(new_n223), .C2(new_n219), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT34), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n278), .B(KEYINPUT64), .Z(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n269), .A2(new_n282), .A3(new_n276), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT32), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT34), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n277), .A2(new_n285), .A3(new_n281), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n283), .A2(KEYINPUT32), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n285), .B1(new_n277), .B2(new_n278), .ZN(new_n289));
  AOI211_X1 g088(.A(KEYINPUT34), .B(new_n282), .C1(new_n269), .C2(new_n276), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G15gat), .B(G43gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(G71gat), .ZN(new_n295));
  INV_X1    g094(.A(G99gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n287), .A2(new_n291), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n287), .B2(new_n291), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n202), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n291), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n298), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n291), .A3(new_n299), .ZN(new_n305));
  XOR2_X1   g104(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT72), .B(G211gat), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT22), .B1(new_n311), .B2(G218gat), .ZN(new_n312));
  XOR2_X1   g111(.A(G197gat), .B(G204gat), .Z(new_n313));
  NOR3_X1   g112(.A1(new_n312), .A2(KEYINPUT73), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n315));
  INV_X1    g114(.A(G211gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G211gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n319), .A3(G218gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT22), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n313), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n315), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n310), .B1(new_n314), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT73), .B1(new_n312), .B2(new_n313), .ZN(new_n326));
  INV_X1    g125(.A(new_n310), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n322), .A2(new_n323), .A3(new_n315), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n221), .A2(new_n222), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n275), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT74), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n242), .A2(KEYINPUT75), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n275), .B(new_n338), .C1(new_n223), .C2(new_n219), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT29), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n331), .B(new_n336), .C1(new_n340), .C2(new_n335), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n339), .A3(new_n335), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343));
  INV_X1    g142(.A(new_n335), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n333), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n330), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347));
  INV_X1    g146(.A(G64gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G92gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n341), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT30), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n341), .B2(new_n346), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n346), .ZN(new_n357));
  INV_X1    g156(.A(new_n351), .ZN(new_n358));
  AND4_X1   g157(.A1(KEYINPUT76), .A2(new_n357), .A3(KEYINPUT30), .A4(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT76), .B1(new_n354), .B2(KEYINPUT30), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n356), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n262), .A2(new_n266), .ZN(new_n363));
  XNOR2_X1  g162(.A(G141gat), .B(G148gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT78), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT2), .ZN(new_n369));
  NAND2_X1  g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n370), .B(KEYINPUT77), .Z(new_n373));
  INV_X1    g172(.A(G155gat), .ZN(new_n374));
  INV_X1    g173(.A(G162gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n372), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  OR2_X1    g176(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(G162gat), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n364), .B1(new_n380), .B2(KEYINPUT2), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n370), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n362), .B1(new_n363), .B2(new_n384), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n365), .A2(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n386), .A2(new_n373), .B1(new_n381), .B2(new_n382), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n259), .A2(KEYINPUT80), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT4), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n363), .A2(new_n384), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT4), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(new_n377), .B2(new_n383), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n387), .A2(new_n394), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(new_n363), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n391), .A2(new_n393), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n363), .A2(new_n384), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n388), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n389), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(KEYINPUT5), .A3(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n377), .A2(new_n383), .A3(new_n394), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n405), .A2(new_n395), .A3(new_n259), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n406), .A2(new_n407), .B1(new_n363), .B2(new_n384), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n385), .B2(new_n388), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n402), .A2(KEYINPUT5), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT0), .B(G57gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G85gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  NAND3_X1  g215(.A1(new_n404), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n412), .ZN(new_n420));
  INV_X1    g219(.A(new_n416), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n419), .B(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n361), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G78gat), .B(G106gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G22gat), .B(G50gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT29), .B1(new_n325), .B2(new_n329), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n384), .B1(new_n429), .B2(KEYINPUT3), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT82), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n329), .B(new_n325), .C1(new_n405), .C2(KEYINPUT29), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n433), .B(new_n384), .C1(new_n429), .C2(KEYINPUT3), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(G228gat), .A2(G233gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n439), .B(new_n430), .C1(new_n438), .C2(new_n432), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT31), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n437), .B2(new_n440), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n428), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n437), .A2(new_n440), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT31), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(new_n442), .A3(new_n427), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n309), .B1(new_n424), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT83), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n361), .A2(KEYINPUT84), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n356), .B(new_n453), .C1(new_n359), .C2(new_n360), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT40), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n392), .B1(new_n398), .B2(KEYINPUT4), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n402), .B1(new_n456), .B2(new_n409), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n401), .A2(new_n402), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n457), .A2(KEYINPUT39), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n416), .B1(new_n457), .B2(KEYINPUT39), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n422), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n459), .A2(new_n460), .A3(new_n455), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n452), .A2(new_n454), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n358), .B1(new_n357), .B2(KEYINPUT38), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT37), .B1(new_n341), .B2(new_n346), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n330), .B1(new_n342), .B2(new_n345), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n336), .B1(new_n340), .B2(new_n335), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(new_n330), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n467), .B1(KEYINPUT37), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT38), .B1(new_n471), .B2(new_n351), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT38), .B1(new_n357), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(new_n467), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n423), .B(new_n466), .C1(new_n472), .C2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(new_n449), .A3(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n448), .B(new_n445), .C1(new_n361), .C2(new_n423), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n309), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n451), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n300), .A2(new_n301), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n443), .A2(new_n444), .A3(new_n428), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n427), .B1(new_n447), .B2(new_n442), .ZN(new_n484));
  OAI211_X1 g283(.A(KEYINPUT35), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n416), .B1(new_n404), .B2(new_n412), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n419), .B(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n487), .B(new_n356), .C1(new_n360), .C2(new_n359), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n452), .A2(new_n454), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n304), .A2(new_n305), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n445), .B2(new_n448), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n487), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n481), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(G1gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT91), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n497), .ZN(new_n501));
  INV_X1    g300(.A(G1gat), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(KEYINPUT16), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(G8gat), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(KEYINPUT92), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n505), .B(new_n506), .C1(new_n503), .C2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT21), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n348), .A2(G57gat), .ZN(new_n515));
  INV_X1    g314(.A(G57gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(G64gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G71gat), .B(G78gat), .Z(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT94), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n517), .B1(new_n521), .B2(new_n515), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n521), .B2(new_n515), .ZN(new_n523));
  INV_X1    g322(.A(new_n519), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n514), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n527), .B(KEYINPUT95), .Z(new_n528));
  AND2_X1   g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n529), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n511), .ZN(new_n533));
  XOR2_X1   g332(.A(G127gat), .B(G155gat), .Z(new_n534));
  XOR2_X1   g333(.A(new_n533), .B(new_n534), .Z(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n537));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n535), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n530), .A2(new_n531), .A3(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n536), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n539), .B1(new_n536), .B2(new_n541), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G134gat), .B(G162gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT86), .ZN(new_n548));
  NOR3_X1   g347(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n549), .A2(KEYINPUT90), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(KEYINPUT90), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553));
  INV_X1    g352(.A(G43gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(KEYINPUT88), .A3(G50gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(G50gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT88), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n554), .A2(G50gat), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n553), .B(new_n555), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n556), .ZN(new_n563));
  OR3_X1    g362(.A1(new_n563), .A2(new_n553), .A3(new_n559), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n552), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G29gat), .ZN(new_n566));
  INV_X1    g365(.A(G36gat), .ZN(new_n567));
  OAI221_X1 g366(.A(new_n565), .B1(new_n561), .B2(new_n560), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n549), .A2(KEYINPUT87), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n548), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n549), .A2(KEYINPUT87), .ZN(new_n571));
  OAI22_X1  g370(.A1(new_n570), .A2(new_n571), .B1(new_n566), .B2(new_n567), .ZN(new_n572));
  INV_X1    g371(.A(new_n564), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G85gat), .A2(G92gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT7), .ZN(new_n577));
  INV_X1    g376(.A(G106gat), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT8), .B1(new_n296), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT97), .B(G85gat), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n577), .B(new_n579), .C1(G92gat), .C2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G99gat), .B(G106gat), .Z(new_n582));
  XOR2_X1   g381(.A(new_n581), .B(new_n582), .Z(new_n583));
  NAND2_X1  g382(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT96), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT41), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n584), .A2(KEYINPUT98), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n590));
  INV_X1    g389(.A(new_n583), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n568), .B2(new_n574), .ZN(new_n592));
  INV_X1    g391(.A(new_n588), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n587), .A2(KEYINPUT41), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n568), .A2(new_n598), .A3(new_n574), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n568), .B2(new_n574), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n591), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n595), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n597), .B1(new_n595), .B2(new_n601), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n604), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT98), .B1(new_n584), .B2(new_n588), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n592), .A2(new_n590), .A3(new_n593), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n601), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n596), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n607), .B1(new_n611), .B2(new_n602), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n546), .B1(new_n606), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n604), .B1(new_n603), .B2(new_n605), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n611), .A2(new_n607), .A3(new_n602), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n545), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n544), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n510), .B1(new_n599), .B2(new_n600), .ZN(new_n619));
  INV_X1    g418(.A(new_n510), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n575), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n510), .A2(new_n568), .A3(new_n574), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n622), .B(KEYINPUT13), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n619), .A2(KEYINPUT18), .A3(new_n621), .A4(new_n622), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT11), .B(G169gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G197gat), .ZN(new_n633));
  XOR2_X1   g432(.A(G113gat), .B(G141gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT85), .Z(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n625), .A2(new_n639), .A3(new_n629), .A4(new_n630), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(G230gat), .ZN(new_n642));
  INV_X1    g441(.A(G233gat), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n526), .A2(KEYINPUT99), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n526), .A2(KEYINPUT99), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n583), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n591), .B1(new_n526), .B2(KEYINPUT99), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n583), .A2(KEYINPUT10), .A3(new_n520), .A4(new_n525), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n644), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n648), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n652), .B1(new_n644), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT100), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n255), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n652), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n653), .A2(new_n644), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n661), .A3(new_n658), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n641), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n496), .A2(new_n618), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n487), .B(KEYINPUT101), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G1gat), .ZN(G1324gat));
  INV_X1    g468(.A(new_n490), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n672));
  OR2_X1    g471(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n676), .B(new_n677), .C1(new_n506), .C2(new_n671), .ZN(G1325gat));
  AOI21_X1  g477(.A(G15gat), .B1(new_n665), .B2(new_n482), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n302), .A2(new_n308), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(G15gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT102), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n679), .B1(new_n665), .B2(new_n682), .ZN(G1326gat));
  INV_X1    g482(.A(new_n449), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n685), .B(new_n687), .ZN(G1327gat));
  NAND2_X1  g487(.A1(new_n496), .A2(new_n617), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n544), .A2(new_n664), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n566), .A3(new_n667), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT45), .ZN(new_n695));
  OR3_X1    g494(.A1(new_n424), .A2(KEYINPUT105), .A3(new_n449), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n680), .B1(new_n478), .B2(KEYINPUT105), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n477), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n495), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n617), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n606), .A2(new_n612), .A3(new_n546), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n545), .B1(new_n614), .B2(new_n615), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n698), .B2(new_n495), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(KEYINPUT107), .A3(new_n700), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n703), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n691), .B(KEYINPUT104), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n666), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n713), .ZN(G1328gat));
  NOR3_X1   g513(.A1(new_n692), .A2(G36gat), .A3(new_n490), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT46), .ZN(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n712), .B2(new_n490), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1329gat));
  OAI21_X1  g517(.A(G43gat), .B1(new_n712), .B2(new_n309), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n693), .A2(new_n554), .A3(new_n482), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(G1330gat));
  XNOR2_X1  g523(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n684), .A3(new_n711), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G50gat), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n692), .A2(G50gat), .A3(new_n449), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n725), .B1(new_n730), .B2(KEYINPUT108), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n728), .B1(new_n726), .B2(G50gat), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733));
  INV_X1    g532(.A(new_n725), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n731), .A2(new_n735), .ZN(G1331gat));
  AND3_X1   g535(.A1(new_n699), .A2(new_n618), .A3(new_n641), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n663), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n666), .B(KEYINPUT110), .Z(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n516), .ZN(G1332gat));
  OAI22_X1  g540(.A1(new_n738), .A2(new_n490), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  INV_X1    g541(.A(new_n738), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n670), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT49), .B(G64gat), .Z(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT111), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n738), .B2(new_n309), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n738), .A2(G71gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(new_n491), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g550(.A1(new_n743), .A2(new_n684), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  INV_X1    g552(.A(new_n544), .ZN(new_n754));
  INV_X1    g553(.A(new_n641), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n699), .A2(KEYINPUT51), .A3(new_n617), .A4(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n708), .A2(KEYINPUT112), .A3(KEYINPUT51), .A4(new_n756), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n708), .A2(new_n756), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n759), .A2(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n663), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n580), .B1(new_n765), .B2(new_n667), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n710), .A2(new_n663), .A3(new_n756), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n666), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n580), .B2(new_n768), .ZN(G1336gat));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  NOR4_X1   g569(.A1(new_n763), .A2(G92gat), .A3(new_n764), .A4(new_n490), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(KEYINPUT114), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n490), .A2(G92gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n765), .A2(KEYINPUT114), .A3(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n710), .A2(new_n663), .A3(new_n670), .A4(new_n756), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G92gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n708), .A2(KEYINPUT113), .A3(new_n756), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n761), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n759), .A2(new_n760), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n764), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n783), .A2(new_n773), .B1(new_n775), .B2(G92gat), .ZN(new_n784));
  OAI22_X1  g583(.A1(new_n772), .A2(new_n777), .B1(new_n784), .B2(new_n770), .ZN(G1337gat));
  NAND3_X1  g584(.A1(new_n765), .A2(new_n296), .A3(new_n482), .ZN(new_n786));
  OAI21_X1  g585(.A(G99gat), .B1(new_n767), .B2(new_n309), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1338gat));
  OAI21_X1  g587(.A(G106gat), .B1(new_n767), .B2(new_n449), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n764), .A2(new_n449), .A3(G106gat), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n789), .B(new_n790), .C1(new_n763), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n781), .A2(new_n782), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n791), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n789), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n793), .B1(new_n796), .B2(new_n790), .ZN(G1339gat));
  NAND3_X1  g596(.A1(new_n650), .A2(new_n644), .A3(new_n651), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n660), .A2(KEYINPUT54), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n658), .B1(new_n652), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(KEYINPUT55), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT55), .B1(new_n799), .B2(new_n801), .ZN(new_n804));
  INV_X1    g603(.A(new_n662), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n631), .ZN(new_n807));
  INV_X1    g606(.A(new_n622), .ZN(new_n808));
  INV_X1    g607(.A(new_n600), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n568), .A2(new_n598), .A3(new_n574), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n620), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n621), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n808), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n621), .A2(new_n626), .A3(new_n628), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT116), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT115), .B(new_n808), .C1(new_n811), .C2(new_n812), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n807), .A2(new_n639), .B1(new_n819), .B2(new_n635), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n806), .B(new_n820), .C1(new_n705), .C2(new_n706), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT117), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n635), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n663), .A3(new_n640), .ZN(new_n824));
  INV_X1    g623(.A(new_n804), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n662), .A3(new_n802), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n826), .B2(new_n641), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n707), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n617), .A2(new_n829), .A3(new_n806), .A4(new_n820), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n822), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n544), .ZN(new_n832));
  NOR4_X1   g631(.A1(new_n544), .A2(new_n617), .A3(new_n755), .A4(new_n663), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(new_n449), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n833), .B1(new_n831), .B2(new_n544), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT118), .B1(new_n838), .B2(new_n684), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n670), .A2(new_n666), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n482), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n641), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n838), .A2(new_n670), .A3(new_n739), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n492), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n247), .A3(new_n755), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n843), .A2(new_n847), .ZN(G1340gat));
  OAI21_X1  g647(.A(G120gat), .B1(new_n842), .B2(new_n764), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n663), .A2(new_n245), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT119), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n849), .B1(new_n845), .B2(new_n851), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n846), .B2(new_n754), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n842), .A2(new_n544), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(G127gat), .ZN(G1342gat));
  NOR3_X1   g654(.A1(new_n845), .A2(G134gat), .A3(new_n707), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT56), .ZN(new_n857));
  OAI21_X1  g656(.A(G134gat), .B1(new_n842), .B2(new_n707), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1343gat));
  AOI21_X1  g658(.A(new_n641), .B1(new_n806), .B2(KEYINPUT121), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n826), .A2(new_n861), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n860), .A2(new_n862), .B1(new_n663), .B2(new_n820), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n822), .B(new_n830), .C1(new_n863), .C2(new_n617), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n833), .B1(new_n864), .B2(new_n544), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT57), .B1(new_n865), .B2(new_n449), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n835), .A2(new_n867), .A3(new_n684), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n841), .A2(new_n309), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT120), .Z(new_n870));
  NAND4_X1  g669(.A1(new_n866), .A2(new_n868), .A3(new_n755), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G141gat), .ZN(new_n872));
  INV_X1    g671(.A(G141gat), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n680), .A2(new_n449), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n844), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n755), .ZN(new_n876));
  XNOR2_X1  g675(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n872), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n872), .B2(new_n876), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n844), .A2(new_n874), .ZN(new_n881));
  OR3_X1    g680(.A1(new_n881), .A2(G148gat), .A3(new_n764), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n825), .A2(KEYINPUT121), .A3(new_n662), .A4(new_n802), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n862), .A2(new_n755), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n617), .B1(new_n885), .B2(new_n824), .ZN(new_n886));
  INV_X1    g685(.A(new_n821), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n544), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n888), .A2(new_n889), .A3(new_n834), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n888), .B2(new_n834), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n867), .B(new_n684), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT57), .B1(new_n838), .B2(new_n449), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n892), .A2(new_n663), .A3(new_n870), .A4(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n883), .B1(new_n894), .B2(G148gat), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n866), .A2(new_n868), .A3(new_n663), .A4(new_n870), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n896), .A2(new_n883), .A3(G148gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n882), .B1(new_n895), .B2(new_n897), .ZN(G1345gat));
  AND3_X1   g697(.A1(new_n866), .A2(new_n868), .A3(new_n870), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n899), .A2(new_n378), .A3(new_n379), .A4(new_n754), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n378), .A2(new_n379), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n901), .B1(new_n881), .B2(new_n544), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n900), .A2(new_n902), .ZN(G1346gat));
  NAND3_X1  g702(.A1(new_n899), .A2(G162gat), .A3(new_n617), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n375), .B1(new_n881), .B2(new_n707), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1347gat));
  AND2_X1   g705(.A1(new_n739), .A2(new_n670), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n840), .A2(new_n482), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G169gat), .B1(new_n908), .B2(new_n641), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n838), .A2(new_n667), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n490), .A2(new_n491), .A3(new_n684), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n755), .A3(new_n270), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n913), .ZN(G1348gat));
  AOI21_X1  g713(.A(G176gat), .B1(new_n912), .B2(new_n663), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n908), .A2(new_n764), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(G176gat), .ZN(G1349gat));
  NAND2_X1  g716(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n840), .A2(new_n754), .A3(new_n482), .A4(new_n907), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G183gat), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n213), .A2(new_n214), .ZN(new_n922));
  AND4_X1   g721(.A1(new_n754), .A2(new_n910), .A3(new_n922), .A4(new_n911), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n919), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  AOI211_X1 g724(.A(new_n918), .B(new_n923), .C1(new_n920), .C2(G183gat), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n908), .B2(new_n707), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(KEYINPUT61), .B(G190gat), .C1(new_n908), .C2(new_n707), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n910), .A2(new_n212), .A3(new_n617), .A4(new_n911), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT125), .Z(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(G1351gat));
  INV_X1    g733(.A(new_n874), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT126), .B1(new_n935), .B2(new_n490), .ZN(new_n936));
  OR3_X1    g735(.A1(new_n935), .A2(KEYINPUT126), .A3(new_n490), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n910), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(G197gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n755), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n892), .A2(new_n893), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n907), .A2(new_n309), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n941), .A2(new_n755), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n943), .B2(new_n939), .ZN(G1352gat));
  NAND3_X1  g743(.A1(new_n941), .A2(new_n663), .A3(new_n942), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G204gat), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n764), .A2(G204gat), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n910), .A2(new_n936), .A3(new_n937), .A4(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n948), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n949));
  XNOR2_X1  g748(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n946), .A2(new_n951), .ZN(G1353gat));
  INV_X1    g751(.A(new_n311), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n938), .A2(new_n754), .A3(new_n953), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n892), .A2(new_n754), .A3(new_n893), .A4(new_n942), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1354gat));
  INV_X1    g757(.A(G218gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n938), .A2(new_n959), .A3(new_n617), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n941), .A2(new_n617), .A3(new_n942), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(new_n959), .ZN(G1355gat));
endmodule


