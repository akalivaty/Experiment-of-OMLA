//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT22), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(G137), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT80), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n194));
  OR2_X1    g008(.A1(KEYINPUT77), .A2(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT77), .A2(G125), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(G140), .A3(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(G125), .A2(G140), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n194), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT77), .B(G125), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n201), .A2(KEYINPUT16), .A3(G140), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n193), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT77), .A2(G125), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT77), .A2(G125), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n194), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n198), .B1(new_n206), .B2(G140), .ZN(new_n209));
  OAI211_X1 g023(.A(G146), .B(new_n208), .C1(new_n209), .C2(new_n194), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n203), .A2(new_n210), .A3(KEYINPUT78), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n200), .A2(new_n202), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT78), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G146), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT76), .ZN(new_n217));
  INV_X1    g031(.A(G119), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G128), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT76), .A3(G119), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n219), .A2(new_n221), .B1(new_n218), .B2(G128), .ZN(new_n222));
  XOR2_X1   g036(.A(KEYINPUT24), .B(G110), .Z(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(G119), .B2(new_n220), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n218), .A2(KEYINPUT23), .A3(G128), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n226), .A2(new_n227), .B1(G119), .B2(new_n220), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G110), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n215), .A2(new_n216), .A3(new_n224), .A4(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n211), .A2(new_n224), .A3(new_n229), .A4(new_n214), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT79), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G125), .B(G140), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n193), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n228), .A2(G110), .B1(new_n222), .B2(new_n223), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n210), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n192), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  AOI211_X1 g053(.A(KEYINPUT80), .B(new_n237), .C1(new_n230), .C2(new_n232), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n191), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G902), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n233), .A2(new_n238), .A3(new_n190), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n247));
  INV_X1    g061(.A(new_n245), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n241), .A2(new_n242), .A3(new_n243), .A4(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(G217), .A2(G902), .ZN(new_n251));
  INV_X1    g065(.A(G217), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(G234), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT75), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n241), .A2(new_n243), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n254), .A2(G902), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G475), .A2(G902), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT92), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n211), .A2(new_n214), .ZN(new_n263));
  INV_X1    g077(.A(G237), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n187), .A3(G214), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT17), .A3(G131), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT90), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n269), .B(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT17), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT90), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n263), .A2(new_n277), .A3(new_n270), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n272), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G113), .B(G122), .ZN(new_n280));
  INV_X1    g094(.A(G104), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT87), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n269), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT18), .B1(new_n269), .B2(new_n283), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(new_n273), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n209), .A2(G146), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n235), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n269), .A2(new_n283), .A3(KEYINPUT18), .A4(G131), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n279), .A2(new_n282), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n274), .B(KEYINPUT88), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n209), .A2(KEYINPUT19), .ZN(new_n293));
  OR2_X1    g107(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n294));
  NAND2_X1  g108(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n234), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n210), .B1(new_n297), .B2(G146), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n290), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n282), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n291), .A2(new_n301), .A3(KEYINPUT91), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT91), .B1(new_n291), .B2(new_n301), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n262), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT20), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n291), .A2(new_n301), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT20), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(new_n262), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(G234), .A2(G237), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n310), .A2(G952), .A3(new_n187), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(G902), .A3(G953), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n312), .B(KEYINPUT97), .Z(new_n313));
  XOR2_X1   g127(.A(KEYINPUT21), .B(G898), .Z(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT3), .B1(new_n281), .B2(G107), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n319));
  INV_X1    g133(.A(G107), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(G104), .ZN(new_n321));
  INV_X1    g135(.A(G101), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n281), .A2(G107), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n318), .A2(new_n321), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT4), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n318), .A2(new_n321), .A3(new_n323), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G101), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n325), .B(new_n327), .ZN(new_n328));
  OR2_X1    g142(.A1(KEYINPUT0), .A2(G128), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT0), .A2(G128), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n266), .A2(G146), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n193), .A2(G143), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n329), .B(new_n330), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n193), .A2(G143), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n266), .A2(G146), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT0), .A4(G128), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n328), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n323), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n281), .A2(G107), .ZN(new_n340));
  OAI21_X1  g154(.A(G101), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n324), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G143), .B(G146), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G128), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n332), .A2(KEYINPUT1), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n344), .B2(G128), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n343), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT65), .ZN(new_n353));
  AOI21_X1  g167(.A(G128), .B1(new_n334), .B2(new_n335), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n335), .A2(new_n345), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n348), .B(KEYINPUT65), .C1(new_n344), .C2(G128), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n346), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT10), .A3(new_n343), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n338), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT11), .ZN(new_n361));
  INV_X1    g175(.A(G134), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(G137), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(G137), .ZN(new_n364));
  INV_X1    g178(.A(G137), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT11), .A3(G134), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G131), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n363), .A2(new_n366), .A3(new_n273), .A4(new_n364), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(KEYINPUT64), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT64), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n367), .A2(new_n371), .A3(G131), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n360), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n338), .A2(new_n373), .A3(new_n352), .A4(new_n359), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G140), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n187), .A2(G227), .ZN(new_n378));
  XOR2_X1   g192(.A(new_n377), .B(new_n378), .Z(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n376), .ZN(new_n381));
  OR3_X1    g195(.A1(new_n358), .A2(new_n343), .A3(KEYINPUT82), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT82), .B1(new_n358), .B2(new_n343), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n350), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n374), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT12), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(KEYINPUT12), .A3(new_n374), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n381), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n380), .B(G469), .C1(new_n389), .C2(new_n379), .ZN(new_n390));
  INV_X1    g204(.A(G469), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n376), .A2(new_n379), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n387), .B2(new_n388), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n379), .B1(new_n375), .B2(new_n376), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n391), .B(new_n242), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(G469), .A2(G902), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n390), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT9), .B(G234), .Z(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G221), .B1(new_n399), .B2(G902), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G116), .B(G122), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(new_n320), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT93), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n220), .A2(G143), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n266), .A2(G128), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n362), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT94), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n406), .A2(KEYINPUT13), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(new_n407), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n406), .A2(KEYINPUT13), .ZN(new_n413));
  INV_X1    g227(.A(new_n407), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n414), .B(KEYINPUT94), .C1(KEYINPUT13), .C2(new_n406), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G134), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n405), .A2(new_n409), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT95), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n405), .A2(KEYINPUT95), .A3(new_n409), .A4(new_n417), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n408), .B(new_n362), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n403), .A2(new_n320), .ZN(new_n424));
  INV_X1    g238(.A(G116), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(KEYINPUT14), .A3(G122), .ZN(new_n426));
  INV_X1    g240(.A(new_n403), .ZN(new_n427));
  OAI211_X1 g241(.A(G107), .B(new_n426), .C1(new_n427), .C2(KEYINPUT14), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n423), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n399), .A2(new_n252), .A3(G953), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n422), .A2(new_n430), .A3(new_n432), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G478), .ZN(new_n437));
  NOR2_X1   g251(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n242), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n432), .B1(new_n422), .B2(new_n430), .ZN(new_n444));
  AOI211_X1 g258(.A(new_n429), .B(new_n433), .C1(new_n420), .C2(new_n421), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n242), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n441), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G475), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n279), .A2(new_n290), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n300), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n291), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n449), .B1(new_n452), .B2(new_n242), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n309), .A2(new_n317), .A3(new_n402), .A4(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n456));
  MUX2_X1   g270(.A(new_n337), .B(new_n358), .S(new_n201), .Z(new_n457));
  NAND2_X1  g271(.A1(new_n187), .A2(G224), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n458), .B(KEYINPUT84), .Z(new_n459));
  NOR2_X1   g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g274(.A(KEYINPUT2), .B(G113), .Z(new_n461));
  XNOR2_X1  g275(.A(G116), .B(G119), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n218), .A2(G116), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n467), .B(G113), .C1(KEYINPUT5), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n342), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n466), .A2(new_n343), .A3(new_n469), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(G110), .B(G122), .Z(new_n474));
  XOR2_X1   g288(.A(KEYINPUT85), .B(KEYINPUT8), .Z(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n460), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n328), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n461), .A2(new_n462), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n464), .B2(new_n465), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n472), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OR2_X1    g295(.A1(new_n481), .A2(new_n474), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n457), .A2(KEYINPUT7), .A3(new_n459), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n457), .A2(KEYINPUT7), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n477), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(KEYINPUT83), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n481), .A2(new_n474), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n481), .B2(new_n474), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n481), .A2(new_n474), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n457), .B(new_n459), .Z(new_n492));
  OAI211_X1 g306(.A(new_n242), .B(new_n485), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n489), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n481), .A2(new_n474), .A3(new_n487), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n482), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n492), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n501), .A2(new_n242), .A3(new_n494), .A4(new_n485), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G214), .B1(G237), .B2(G902), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n456), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  AOI211_X1 g320(.A(KEYINPUT86), .B(new_n506), .C1(new_n496), .C2(new_n502), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n455), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT31), .ZN(new_n510));
  INV_X1    g324(.A(new_n364), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n362), .A2(G137), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n513), .A2(new_n369), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n358), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT68), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n370), .A2(new_n337), .A3(new_n372), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n358), .A2(new_n518), .A3(new_n514), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n516), .A2(KEYINPUT30), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n518), .B1(new_n358), .B2(new_n514), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n370), .A2(new_n372), .A3(new_n337), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n525), .A2(KEYINPUT69), .A3(KEYINPUT30), .A4(new_n519), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT66), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n515), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n358), .A2(KEYINPUT66), .A3(new_n514), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n517), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n480), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT26), .B(G101), .Z(new_n535));
  NAND3_X1  g349(.A1(new_n264), .A2(new_n187), .A3(G210), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n525), .A2(new_n480), .A3(new_n519), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n534), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n540), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n527), .B2(new_n533), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(KEYINPUT71), .A3(new_n539), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n510), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n534), .A2(new_n510), .A3(new_n539), .A4(new_n540), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT72), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT72), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n545), .A2(new_n550), .A3(new_n510), .A4(new_n539), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT28), .ZN(new_n553));
  INV_X1    g367(.A(new_n480), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n531), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n555), .B2(new_n540), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT73), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n480), .A2(new_n515), .A3(new_n517), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n553), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n539), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n547), .A2(new_n552), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G472), .A2(G902), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT74), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  AND4_X1   g379(.A1(KEYINPUT71), .A2(new_n534), .A3(new_n539), .A4(new_n540), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT71), .B1(new_n545), .B2(new_n539), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT31), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n556), .A2(KEYINPUT73), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n556), .A2(KEYINPUT73), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n560), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n539), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n568), .A2(new_n573), .A3(new_n549), .A4(new_n551), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT74), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n563), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT32), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n563), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT32), .ZN(new_n579));
  INV_X1    g393(.A(G472), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT29), .ZN(new_n581));
  INV_X1    g395(.A(new_n545), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n572), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n581), .B(new_n583), .C1(new_n571), .C2(new_n572), .ZN(new_n584));
  INV_X1    g398(.A(new_n560), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n554), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n540), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n585), .B1(new_n588), .B2(KEYINPUT28), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n572), .A2(new_n581), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  OAI22_X1  g406(.A1(new_n578), .A2(new_n579), .B1(new_n580), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n260), .B(new_n509), .C1(new_n577), .C2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  AOI21_X1  g409(.A(new_n580), .B1(new_n574), .B2(new_n242), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n565), .B2(new_n576), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n434), .A2(new_n598), .A3(new_n435), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT33), .B1(new_n444), .B2(new_n445), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(G478), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n436), .A2(new_n437), .A3(new_n242), .ZN(new_n602));
  NAND2_X1  g416(.A1(G478), .A2(G902), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n308), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n304), .B2(KEYINPUT20), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n606), .B2(new_n453), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n506), .B1(new_n496), .B2(new_n502), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n607), .A2(new_n609), .A3(new_n316), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n255), .A2(new_n258), .A3(new_n402), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n597), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT34), .B(G104), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  INV_X1    g428(.A(new_n453), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n448), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n316), .B(KEYINPUT99), .Z(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n608), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT91), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n306), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n291), .A2(new_n301), .A3(KEYINPUT91), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n307), .B1(new_n624), .B2(new_n262), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n307), .B(new_n262), .C1(new_n302), .C2(new_n303), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n620), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n305), .A2(KEYINPUT98), .A3(new_n626), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n616), .B(new_n619), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n597), .A3(new_n611), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NOR2_X1   g447(.A1(new_n239), .A2(new_n240), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT36), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n635), .A3(new_n190), .ZN(new_n636));
  OAI22_X1  g450(.A1(new_n239), .A2(new_n240), .B1(KEYINPUT36), .B2(new_n191), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n636), .A2(new_n637), .A3(new_n257), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n255), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n255), .A2(KEYINPUT100), .A3(new_n639), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n597), .A2(new_n642), .A3(new_n509), .A4(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n644), .B(KEYINPUT37), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G110), .ZN(G12));
  AOI21_X1  g460(.A(KEYINPUT100), .B1(new_n255), .B2(new_n639), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n641), .B(new_n638), .C1(new_n250), .C2(new_n254), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n647), .A2(new_n648), .A3(new_n401), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n574), .A2(new_n575), .A3(new_n563), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n575), .B1(new_n574), .B2(new_n563), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n579), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n580), .B1(new_n584), .B2(new_n591), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n562), .A2(new_n564), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n653), .B1(new_n654), .B2(KEYINPUT32), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n313), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n311), .ZN(new_n659));
  AOI211_X1 g473(.A(new_n659), .B(new_n616), .C1(new_n628), .C2(new_n629), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n649), .A2(new_n656), .A3(new_n608), .A4(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT101), .B(G128), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G30));
  XNOR2_X1  g477(.A(new_n659), .B(KEYINPUT39), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n402), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT40), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n503), .B(KEYINPUT38), .Z(new_n668));
  NOR3_X1   g482(.A1(new_n667), .A2(new_n506), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n566), .A2(new_n567), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n588), .A2(new_n572), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT102), .Z(new_n672));
  OAI21_X1  g486(.A(new_n242), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n652), .B(new_n674), .C1(new_n579), .C2(new_n578), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n647), .A2(new_n648), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n309), .A2(new_n615), .B1(new_n443), .B2(new_n447), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n669), .A2(new_n675), .A3(new_n677), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  INV_X1    g494(.A(new_n659), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n604), .B(new_n681), .C1(new_n606), .C2(new_n453), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n649), .A2(new_n656), .A3(new_n608), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  OR2_X1    g499(.A1(new_n393), .A2(new_n394), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n242), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G469), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n400), .A3(new_n395), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT103), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n656), .A2(new_n260), .A3(new_n610), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND4_X1  g507(.A1(new_n656), .A2(new_n260), .A3(new_n630), .A4(new_n690), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  NOR4_X1   g509(.A1(new_n606), .A2(new_n316), .A3(new_n453), .A4(new_n448), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n577), .B2(new_n593), .ZN(new_n697));
  INV_X1    g511(.A(new_n689), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n642), .A2(new_n608), .A3(new_n643), .A4(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT104), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  OAI21_X1  g516(.A(G472), .B1(new_n562), .B2(G902), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n589), .A2(KEYINPUT105), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n589), .A2(KEYINPUT105), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n572), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n568), .A2(new_n549), .A3(new_n551), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n563), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n259), .ZN(new_n710));
  INV_X1    g524(.A(new_n619), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n678), .A4(new_n690), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  NOR2_X1   g527(.A1(new_n709), .A2(new_n682), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n676), .A2(new_n714), .A3(new_n608), .A4(new_n698), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  AOI21_X1  g530(.A(new_n259), .B1(new_n652), .B2(new_n655), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n401), .B(KEYINPUT106), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n503), .A2(new_n506), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n717), .A2(new_n683), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT107), .B1(new_n578), .B2(new_n579), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n725));
  AOI211_X1 g539(.A(new_n725), .B(KEYINPUT32), .C1(new_n574), .C2(new_n563), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n259), .B1(new_n727), .B2(new_n655), .ZN(new_n728));
  INV_X1    g542(.A(new_n720), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n659), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n718), .A2(new_n607), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n728), .A2(KEYINPUT42), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n723), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  AND4_X1   g548(.A1(new_n717), .A2(new_n660), .A3(new_n719), .A4(new_n720), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n362), .ZN(G36));
  INV_X1    g550(.A(new_n379), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n387), .A2(new_n388), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n737), .B1(new_n738), .B2(new_n381), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n380), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(KEYINPUT45), .A3(new_n380), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(G469), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n396), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n744), .A2(KEYINPUT46), .A3(new_n396), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n395), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n400), .A3(new_n665), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n615), .B(new_n604), .C1(new_n625), .C2(new_n605), .ZN(new_n751));
  NAND2_X1  g565(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n752));
  OR2_X1    g566(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n606), .A2(new_n453), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT43), .A3(new_n604), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n751), .A2(KEYINPUT109), .A3(new_n752), .A4(new_n753), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n597), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n676), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n729), .B(new_n750), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n760), .A2(KEYINPUT44), .A3(new_n761), .A4(new_n676), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n765), .A2(new_n766), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G137), .ZN(G39));
  NAND2_X1  g585(.A1(new_n749), .A2(new_n400), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT47), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n652), .A2(new_n655), .A3(new_n259), .A4(new_n720), .ZN(new_n774));
  OR3_X1    g588(.A1(new_n773), .A2(new_n682), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  NOR2_X1   g590(.A1(new_n675), .A2(new_n259), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n729), .A2(new_n689), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n777), .A2(new_n311), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n604), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n757), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT114), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n760), .A2(new_n311), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n778), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n677), .A3(new_n709), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n783), .A2(new_n710), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n688), .A2(new_n395), .ZN(new_n787));
  INV_X1    g601(.A(new_n400), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n729), .B1(new_n773), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n785), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n786), .A2(new_n698), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n668), .A2(new_n506), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(KEYINPUT50), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n792), .A2(new_n796), .A3(new_n793), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n782), .B(new_n791), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT51), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n508), .A2(new_n617), .ZN(new_n800));
  INV_X1    g614(.A(new_n607), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n597), .A2(new_n611), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n594), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n594), .A2(new_n802), .A3(KEYINPUT111), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n401), .B1(new_n628), .B2(new_n629), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n656), .A2(new_n454), .A3(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n709), .A2(new_n607), .A3(new_n718), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n676), .B(new_n730), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n691), .A2(new_n694), .A3(new_n712), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n616), .A2(new_n606), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n597), .A2(new_n611), .A3(new_n800), .A4(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n644), .B(new_n814), .C1(new_n697), .C2(new_n699), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n807), .A2(new_n811), .A3(new_n812), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n735), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n733), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n661), .A2(new_n715), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n678), .A2(new_n608), .A3(new_n402), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n640), .A2(new_n659), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n675), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(KEYINPUT52), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n661), .A2(KEYINPUT112), .A3(new_n715), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n823), .A2(new_n684), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n661), .A2(new_n826), .A3(new_n684), .A4(new_n715), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT53), .B1(new_n820), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n830), .B(KEYINPUT52), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n735), .B1(new_n723), .B2(new_n732), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n691), .A2(new_n694), .A3(new_n712), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n815), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n836), .A2(new_n811), .A3(new_n838), .A4(new_n807), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n835), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT54), .B1(new_n834), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n820), .A2(new_n833), .A3(KEYINPUT53), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n835), .B2(new_n839), .ZN(new_n844));
  XNOR2_X1  g658(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n799), .A2(new_n842), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(G952), .B(new_n187), .C1(new_n792), .C2(new_n609), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n801), .B2(new_n779), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n783), .A2(new_n728), .A3(new_n778), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT48), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT115), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n848), .A2(new_n854), .B1(G952), .B2(G953), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n787), .B(KEYINPUT49), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n504), .A2(new_n856), .A3(new_n604), .A4(new_n668), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n777), .A2(new_n400), .A3(new_n757), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n858), .ZN(G75));
  NAND2_X1  g673(.A1(new_n491), .A2(new_n492), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n860), .A2(new_n501), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT55), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n242), .B1(new_n843), .B2(new_n844), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT116), .B1(new_n864), .B2(G210), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT56), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n820), .A2(new_n833), .A3(KEYINPUT53), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n830), .B(new_n831), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT53), .B1(new_n820), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(G210), .B(G902), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n868), .A2(new_n872), .A3(new_n863), .A4(new_n866), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n862), .B1(new_n867), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n187), .A2(G952), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n872), .A2(new_n868), .A3(new_n866), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT55), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n865), .A2(new_n863), .A3(new_n866), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n879), .A3(new_n861), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n874), .A2(new_n876), .A3(new_n880), .ZN(G51));
  NAND2_X1  g695(.A1(new_n843), .A2(new_n844), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n845), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n847), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n882), .A2(KEYINPUT118), .A3(new_n845), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n396), .B(KEYINPUT117), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n686), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n744), .B(KEYINPUT119), .Z(new_n892));
  NAND2_X1  g706(.A1(new_n864), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n875), .B1(new_n891), .B2(new_n893), .ZN(G54));
  AND2_X1   g708(.A1(new_n864), .A2(KEYINPUT58), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n895), .A2(G475), .A3(new_n624), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n624), .B1(new_n895), .B2(G475), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n875), .ZN(G60));
  NAND2_X1  g712(.A1(new_n599), .A2(new_n600), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n603), .B(KEYINPUT59), .ZN(new_n900));
  AND4_X1   g714(.A1(new_n899), .A2(new_n885), .A3(new_n886), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n842), .A2(new_n847), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n899), .B1(new_n902), .B2(new_n900), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n901), .A2(new_n903), .A3(new_n875), .ZN(G63));
  AND2_X1   g718(.A1(new_n636), .A2(new_n637), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n251), .B(KEYINPUT60), .Z(new_n906));
  NAND3_X1  g720(.A1(new_n882), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n882), .A2(new_n906), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n256), .B(KEYINPUT122), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n882), .A2(KEYINPUT121), .A3(new_n905), .A4(new_n906), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n909), .A2(new_n912), .A3(new_n876), .A4(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n914), .A2(KEYINPUT120), .A3(KEYINPUT61), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT61), .B1(new_n914), .B2(KEYINPUT120), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(G66));
  AND2_X1   g731(.A1(new_n838), .A2(new_n807), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(G953), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n187), .B1(new_n314), .B2(G224), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT123), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n491), .B1(G898), .B2(new_n187), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n922), .B(new_n923), .Z(G69));
  AOI22_X1  g738(.A1(new_n522), .A2(new_n526), .B1(new_n532), .B2(new_n531), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(new_n297), .Z(new_n926));
  NAND2_X1  g740(.A1(G900), .A2(G953), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n762), .A2(new_n763), .ZN(new_n929));
  INV_X1    g743(.A(new_n750), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n720), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n769), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n767), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n823), .A2(new_n684), .A3(new_n828), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n928), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n930), .A2(new_n728), .A3(new_n608), .A4(new_n678), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n936), .A2(KEYINPUT125), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n735), .B1(new_n936), .B2(KEYINPUT125), .ZN(new_n938));
  AND4_X1   g752(.A1(new_n733), .A2(new_n775), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n823), .A2(new_n684), .A3(new_n828), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n770), .A3(KEYINPUT124), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n935), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n926), .B(new_n927), .C1(new_n942), .C2(G953), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n823), .A2(new_n679), .A3(new_n684), .A4(new_n828), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n770), .A2(new_n775), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n801), .A2(new_n813), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n948), .A2(new_n666), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n717), .A2(new_n949), .A3(new_n720), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n946), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n951), .A2(new_n187), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n943), .B1(new_n952), .B2(new_n926), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G72));
  NAND4_X1  g769(.A1(new_n946), .A2(new_n918), .A3(new_n947), .A4(new_n950), .ZN(new_n956));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n539), .A3(new_n582), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n583), .B1(new_n566), .B2(new_n567), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n958), .B(new_n961), .C1(new_n834), .C2(new_n841), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n935), .A2(new_n941), .A3(new_n918), .A4(new_n939), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n958), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(KEYINPUT126), .A3(new_n958), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n967), .A2(new_n572), .A3(new_n545), .A4(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n963), .A2(new_n969), .A3(KEYINPUT127), .A4(new_n876), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n971));
  INV_X1    g785(.A(new_n969), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n960), .A2(new_n876), .A3(new_n962), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n974), .ZN(G57));
endmodule


