//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(G58), .A2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n225), .A2(G50), .A3(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n206), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n211), .A2(new_n222), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XOR2_X1   g0044(.A(G58), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT67), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  NAND2_X1  g0052(.A1(new_n207), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n229), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT72), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n206), .A2(G33), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n258), .A2(new_n213), .B1(new_n206), .B2(G68), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n254), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT11), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n261), .ZN(new_n263));
  INV_X1    g0063(.A(G13), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n264), .A2(new_n206), .A3(G1), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OR3_X1    g0066(.A1(new_n266), .A2(KEYINPUT12), .A3(G68), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT12), .B1(new_n266), .B2(G68), .ZN(new_n268));
  INV_X1    g0068(.A(new_n229), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n207), .B2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n266), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G68), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n205), .B2(G20), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n267), .A2(new_n268), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n262), .A2(new_n263), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G238), .ZN(new_n284));
  OR2_X1    g0084(.A1(new_n277), .A2(new_n282), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT71), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n283), .B(KEYINPUT71), .C1(new_n284), .C2(new_n285), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G97), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G226), .ZN(new_n295));
  INV_X1    g0095(.A(G232), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(G1698), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n291), .B1(new_n294), .B2(new_n295), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n298), .A2(KEYINPUT70), .A3(new_n277), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT70), .B1(new_n298), .B2(new_n277), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n290), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT13), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT13), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n303), .B(new_n290), .C1(new_n299), .C2(new_n300), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT14), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(new_n306), .A3(G169), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n302), .A2(G179), .A3(new_n304), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n306), .B1(new_n305), .B2(G169), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n276), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n276), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n305), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n302), .B2(new_n304), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n311), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n255), .A2(G150), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n258), .ZN(new_n322));
  INV_X1    g0122(.A(G50), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n206), .B1(new_n223), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n254), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n205), .A2(G20), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G50), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n325), .B1(G50), .B2(new_n266), .C1(new_n271), .C2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT9), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n283), .B1(new_n295), .B2(new_n285), .ZN(new_n330));
  INV_X1    g0130(.A(G33), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT3), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G33), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(new_n293), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(G223), .B1(G77), .B2(new_n335), .ZN(new_n337));
  INV_X1    g0137(.A(G222), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(new_n294), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n330), .B1(new_n339), .B2(new_n277), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G190), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT69), .B(G200), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n329), .B(new_n341), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT10), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n328), .B1(new_n340), .B2(G169), .ZN(new_n345));
  INV_X1    g0145(.A(G179), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n345), .A2(KEYINPUT68), .B1(new_n346), .B2(new_n340), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(KEYINPUT68), .B2(new_n345), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n321), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n326), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n271), .A2(new_n351), .B1(new_n266), .B2(new_n350), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT7), .B1(new_n335), .B2(new_n206), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  AOI211_X1 g0154(.A(new_n354), .B(G20), .C1(new_n332), .C2(new_n334), .ZN(new_n355));
  OAI21_X1  g0155(.A(G68), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT73), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n354), .B1(new_n292), .B2(G20), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n333), .A2(G33), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n331), .A2(KEYINPUT3), .ZN(new_n361));
  OAI211_X1 g0161(.A(KEYINPUT7), .B(new_n206), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(KEYINPUT73), .A3(G68), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(G58), .A2(G68), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n366), .B2(new_n223), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n255), .A2(G159), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n270), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n359), .A2(KEYINPUT74), .A3(new_n362), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT74), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n374), .B(new_n354), .C1(new_n292), .C2(G20), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(G68), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n369), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n370), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n352), .B1(new_n372), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT76), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n332), .A2(new_n334), .A3(G223), .A4(new_n293), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G87), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n332), .A2(new_n334), .A3(G226), .A4(G1698), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT75), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n292), .A2(KEYINPUT75), .A3(G226), .A4(G1698), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n277), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n381), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n387), .A2(new_n388), .ZN(new_n392));
  OAI211_X1 g0192(.A(KEYINPUT76), .B(new_n277), .C1(new_n392), .C2(new_n384), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n283), .B1(new_n296), .B2(new_n285), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(G179), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n391), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G169), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n389), .A2(new_n390), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(new_n394), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT18), .B1(new_n380), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n394), .A2(G190), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n391), .A2(new_n393), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n315), .B1(new_n398), .B2(new_n394), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT73), .B1(new_n363), .B2(G68), .ZN(new_n406));
  AOI211_X1 g0206(.A(new_n357), .B(new_n273), .C1(new_n359), .C2(new_n362), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n371), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n379), .A2(new_n254), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n352), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n409), .A2(new_n410), .ZN(new_n414));
  INV_X1    g0214(.A(new_n400), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n380), .A2(KEYINPUT17), .A3(new_n405), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n401), .A2(new_n413), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n326), .A2(G77), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n271), .A2(new_n420), .B1(G77), .B2(new_n266), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n350), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT15), .B(G87), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n258), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n421), .B1(new_n254), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n285), .ZN(new_n426));
  AOI22_X1  g0226(.A1(G244), .A2(new_n426), .B1(new_n279), .B2(new_n282), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n297), .A2(new_n284), .B1(new_n215), .B2(new_n292), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n294), .A2(new_n296), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n277), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n425), .B1(new_n431), .B2(new_n397), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n427), .A2(new_n346), .A3(new_n430), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n342), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n436), .B(new_n425), .C1(new_n313), .C2(new_n431), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NOR4_X1   g0238(.A1(new_n319), .A2(new_n349), .A3(new_n419), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G116), .ZN(new_n440));
  OAI221_X1 g0240(.A(new_n440), .B1(new_n294), .B2(new_n284), .C1(new_n214), .C2(new_n297), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n277), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n390), .B(G250), .C1(G1), .C2(new_n281), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n281), .A2(G1), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n279), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n342), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n441), .B2(new_n277), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n313), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n292), .A2(new_n206), .A3(G68), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT19), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n206), .B1(new_n291), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(G87), .B2(new_n203), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n258), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n453), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n254), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n423), .A2(new_n265), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n205), .A2(G33), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n270), .A2(new_n266), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G87), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n452), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT81), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n442), .A2(new_n346), .A3(new_n447), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n460), .B(new_n461), .C1(new_n423), .C2(new_n464), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n472), .C1(G169), .C2(new_n450), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n292), .A2(new_n206), .A3(G87), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT22), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT23), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(new_n215), .A3(G20), .ZN(new_n479));
  INV_X1    g0279(.A(G116), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n477), .B(new_n479), .C1(new_n480), .C2(new_n258), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT84), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g0284(.A(KEYINPUT83), .B(KEYINPUT24), .Z(new_n485));
  AND2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n484), .A2(new_n485), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n254), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n265), .A2(KEYINPUT25), .A3(new_n215), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT25), .B1(new_n265), .B2(new_n215), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n464), .A2(new_n215), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT5), .B(G41), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n444), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n496), .A2(new_n390), .A3(G264), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT85), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n496), .A2(new_n278), .A3(new_n277), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n292), .A2(G257), .A3(G1698), .ZN(new_n500));
  INV_X1    g0300(.A(G294), .ZN(new_n501));
  INV_X1    g0301(.A(G250), .ZN(new_n502));
  OAI221_X1 g0302(.A(new_n500), .B1(new_n331), .B2(new_n501), .C1(new_n294), .C2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n499), .B1(new_n503), .B2(new_n277), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n397), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n498), .A2(new_n346), .A3(new_n504), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n494), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n473), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n467), .B1(new_n449), .B2(new_n451), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT81), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n505), .A2(G200), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n498), .A2(G190), .A3(new_n504), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n488), .A2(new_n512), .A3(new_n493), .A4(new_n513), .ZN(new_n514));
  AND4_X1   g0314(.A1(new_n474), .A2(new_n508), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n465), .A2(G116), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n265), .A2(new_n480), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n253), .A2(new_n229), .B1(G20), .B2(new_n480), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n519), .B(new_n206), .C1(G33), .C2(new_n457), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n518), .A2(KEYINPUT20), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT20), .B1(new_n518), .B2(new_n520), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n516), .B(new_n517), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n292), .A2(G257), .A3(new_n293), .ZN(new_n524));
  INV_X1    g0324(.A(G303), .ZN(new_n525));
  OAI221_X1 g0325(.A(new_n524), .B1(new_n525), .B2(new_n292), .C1(new_n297), .C2(new_n216), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n277), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n277), .B1(new_n444), .B2(new_n495), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n499), .B1(G270), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n523), .B1(new_n530), .B2(G200), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n313), .B2(new_n530), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n523), .A2(new_n530), .A3(G169), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT21), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n530), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(G179), .A3(new_n523), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n523), .A2(new_n530), .A3(KEYINPUT21), .A4(G169), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n532), .A2(new_n535), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT82), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n537), .A2(new_n538), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n542), .A2(KEYINPUT82), .A3(new_n535), .A4(new_n532), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT80), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n464), .A2(G97), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT77), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n266), .A2(new_n457), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n373), .A2(G107), .A3(new_n375), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n215), .A2(KEYINPUT6), .A3(G97), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n457), .A2(new_n215), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(new_n202), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n555), .B2(KEYINPUT6), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n270), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  OR3_X1    g0358(.A1(new_n551), .A2(KEYINPUT79), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT79), .B1(new_n551), .B2(new_n558), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n294), .B2(new_n214), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n336), .A2(G250), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n292), .A2(KEYINPUT4), .A3(G244), .A4(new_n293), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n519), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n277), .ZN(new_n566));
  INV_X1    g0366(.A(new_n499), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n528), .A2(G257), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G179), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(G169), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n559), .A2(new_n560), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n313), .B1(new_n315), .B2(KEYINPUT78), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n551), .A2(new_n558), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n569), .A2(KEYINPUT78), .A3(G200), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n545), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n559), .A2(new_n560), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n571), .A2(new_n572), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(KEYINPUT80), .A3(new_n578), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n515), .A2(new_n544), .A3(new_n580), .A4(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n439), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g0387(.A(new_n587), .B(KEYINPUT86), .Z(G372));
  OAI211_X1 g0388(.A(new_n433), .B(new_n432), .C1(new_n314), .C2(new_n316), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n311), .A2(KEYINPUT88), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT88), .B1(new_n311), .B2(new_n589), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n413), .A2(new_n418), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n401), .A2(new_n417), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n344), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n573), .A2(new_n579), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n508), .A2(new_n535), .A3(new_n542), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT87), .B1(new_n462), .B2(new_n466), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n462), .A2(KEYINPUT87), .A3(new_n466), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n452), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n514), .A2(new_n473), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n474), .A2(new_n511), .A3(new_n573), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT26), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n599), .A2(new_n598), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n509), .B1(new_n605), .B2(new_n452), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT26), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n576), .B1(new_n571), .B2(new_n572), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n602), .A2(new_n604), .A3(new_n473), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n439), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n595), .A2(new_n348), .A3(new_n611), .ZN(G369));
  NAND3_X1  g0412(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n613), .A2(KEYINPUT27), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(KEYINPUT27), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(G213), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G343), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n523), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n544), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n542), .A2(new_n535), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(new_n619), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(KEYINPUT89), .A3(G330), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT89), .ZN(new_n626));
  INV_X1    g0426(.A(G330), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n494), .A2(new_n506), .A3(new_n507), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n494), .A2(new_n618), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n514), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n508), .A2(new_n618), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n621), .A2(new_n618), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n633), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(G399));
  NAND2_X1  g0438(.A1(new_n209), .A2(new_n280), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G1), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n227), .B2(new_n639), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n642), .B(KEYINPUT28), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n603), .A2(new_n607), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT91), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n606), .A2(KEYINPUT26), .A3(new_n608), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT91), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n603), .A2(new_n647), .A3(new_n607), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n602), .A2(new_n473), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n618), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(KEYINPUT29), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n610), .A2(new_n652), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT29), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n580), .A2(new_n584), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n658), .A2(new_n544), .A3(new_n515), .A4(new_n652), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT31), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n498), .A2(new_n450), .A3(new_n504), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n566), .A2(new_n568), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT90), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n530), .B2(new_n346), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n536), .A2(KEYINPUT90), .A3(G179), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT30), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n663), .A2(KEYINPUT30), .A3(new_n665), .A4(new_n666), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n536), .A2(G179), .A3(new_n450), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n505), .A3(new_n569), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n660), .B1(new_n673), .B2(new_n618), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n673), .A2(new_n660), .A3(new_n618), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n627), .B1(new_n659), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n657), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n643), .B1(new_n681), .B2(G1), .ZN(G364));
  INV_X1    g0482(.A(new_n629), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n264), .A2(G20), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT92), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G45), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G1), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n639), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n683), .B(new_n689), .C1(G330), .C2(new_n624), .ZN(new_n690));
  INV_X1    g0490(.A(new_n689), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n209), .A2(new_n292), .ZN(new_n692));
  INV_X1    g0492(.A(G355), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n692), .A2(new_n693), .B1(G116), .B2(new_n209), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n247), .A2(G45), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n209), .A2(new_n335), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n228), .B2(new_n281), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n694), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(G13), .A2(G33), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G20), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n229), .B1(G20), .B2(new_n397), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n691), .B1(new_n698), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n702), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n206), .A2(new_n346), .ZN(new_n707));
  NOR2_X1   g0507(.A1(G190), .A2(G200), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n292), .B1(new_n709), .B2(new_n213), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(G200), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G190), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n206), .A2(G179), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n708), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G159), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n713), .A2(new_n273), .B1(new_n717), .B2(KEYINPUT32), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n707), .A2(G190), .A3(new_n315), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n710), .B(new_n718), .C1(G58), .C2(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n313), .A2(G179), .A3(G200), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n206), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n457), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n711), .A2(new_n313), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n323), .ZN(new_n727));
  AOI211_X1 g0527(.A(new_n724), .B(new_n727), .C1(KEYINPUT32), .C2(new_n717), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n435), .A2(new_n714), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G190), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G107), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n729), .A2(new_n313), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G87), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n721), .A2(new_n728), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT33), .B(G317), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n712), .A2(new_n735), .B1(new_n720), .B2(G322), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT93), .ZN(new_n737));
  INV_X1    g0537(.A(G311), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n335), .B1(new_n709), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(G329), .B2(new_n716), .ZN(new_n740));
  INV_X1    g0540(.A(new_n723), .ZN(new_n741));
  AOI22_X1  g0541(.A1(G294), .A2(new_n741), .B1(new_n725), .B2(G326), .ZN(new_n742));
  AOI22_X1  g0542(.A1(G283), .A2(new_n730), .B1(new_n732), .B2(G303), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n737), .A2(new_n740), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n706), .B1(new_n734), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n705), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n701), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n746), .B1(new_n624), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n690), .A2(new_n748), .ZN(G396));
  NOR2_X1   g0549(.A1(new_n434), .A2(new_n618), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n437), .B1(new_n425), .B2(new_n652), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n750), .B1(new_n434), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n610), .A2(new_n652), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n654), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n752), .B(KEYINPUT96), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n691), .B1(new_n756), .B2(new_n679), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(new_n679), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n706), .A2(new_n700), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n691), .B1(G77), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT94), .Z(new_n761));
  INV_X1    g0561(.A(new_n709), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n720), .A2(G143), .B1(new_n762), .B2(G159), .ZN(new_n763));
  INV_X1    g0563(.A(G150), .ZN(new_n764));
  INV_X1    g0564(.A(G137), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n763), .B1(new_n713), .B2(new_n764), .C1(new_n765), .C2(new_n726), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT34), .Z(new_n767));
  NAND2_X1  g0567(.A1(new_n730), .A2(G68), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n732), .A2(G50), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n741), .A2(G58), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n335), .B1(new_n716), .B2(G132), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n768), .A2(new_n769), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n335), .B1(new_n715), .B2(new_n738), .C1(new_n719), .C2(new_n501), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n724), .B(new_n773), .C1(G303), .C2(new_n725), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n730), .A2(G87), .ZN(new_n775));
  INV_X1    g0575(.A(new_n732), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n774), .B(new_n775), .C1(new_n215), .C2(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n712), .A2(G283), .B1(new_n762), .B2(G116), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT95), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n767), .A2(new_n772), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n761), .B1(new_n780), .B2(new_n702), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n752), .B2(new_n700), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n758), .A2(new_n782), .ZN(G384));
  OR2_X1    g0583(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n784), .A2(G116), .A3(new_n230), .A4(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT36), .Z(new_n787));
  OR3_X1    g0587(.A1(new_n227), .A2(new_n213), .A3(new_n366), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n323), .A2(G68), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n205), .B(G13), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n594), .A2(new_n616), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n750), .B(KEYINPUT97), .Z(new_n793));
  NAND2_X1  g0593(.A1(new_n753), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n276), .A2(new_n618), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n311), .A2(new_n318), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n305), .A2(G169), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(KEYINPUT14), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(new_n308), .A3(new_n307), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n276), .B(new_n618), .C1(new_n799), .C2(new_n317), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT98), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n377), .B1(new_n406), .B2(new_n407), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n370), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n803), .B(new_n352), .C1(new_n372), .C2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n369), .B1(new_n358), .B2(new_n364), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n254), .B(new_n408), .C1(new_n807), .C2(KEYINPUT16), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT98), .B1(new_n808), .B2(new_n410), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n806), .A2(new_n809), .A3(new_n616), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n419), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT37), .ZN(new_n812));
  AOI21_X1  g0612(.A(KEYINPUT16), .B1(new_n365), .B2(new_n377), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n408), .A2(new_n254), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n410), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n803), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n400), .A2(new_n616), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n808), .A2(KEYINPUT98), .A3(new_n410), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n812), .B1(new_n819), .B2(new_n411), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n414), .A2(new_n415), .ZN(new_n821));
  INV_X1    g0621(.A(new_n616), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n414), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n821), .A2(new_n823), .A3(new_n812), .A4(new_n411), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n811), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n811), .B(KEYINPUT38), .C1(new_n820), .C2(new_n825), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n828), .A2(KEYINPUT99), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT99), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n826), .A2(new_n831), .A3(new_n827), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n792), .B1(new_n802), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT100), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n799), .A2(new_n276), .A3(new_n652), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n829), .A2(KEYINPUT99), .ZN(new_n838));
  INV_X1    g0638(.A(new_n411), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n806), .A2(new_n809), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(new_n840), .B2(new_n817), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n824), .B1(new_n841), .B2(new_n812), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT38), .B1(new_n842), .B2(new_n811), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n832), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT39), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT101), .ZN(new_n847));
  INV_X1    g0647(.A(new_n419), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n821), .A2(new_n823), .A3(new_n411), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n848), .A2(new_n823), .B1(new_n850), .B2(new_n825), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n827), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT39), .B1(new_n852), .B2(new_n829), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n846), .A2(new_n847), .A3(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n830), .B2(new_n832), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT101), .B1(new_n858), .B2(new_n853), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n837), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n835), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n653), .A2(new_n439), .A3(new_n656), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n348), .A3(new_n595), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n862), .B(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n676), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n585), .A2(new_n618), .B1(new_n866), .B2(new_n674), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(new_n801), .A3(new_n752), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT102), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n844), .A2(new_n845), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT102), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(KEYINPUT40), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n869), .B(new_n870), .C1(new_n868), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n852), .A2(new_n829), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT40), .B1(new_n875), .B2(new_n868), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n439), .A2(new_n867), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n627), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n878), .B2(new_n877), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n865), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n205), .B2(new_n685), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n865), .A2(new_n880), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n791), .B1(new_n882), .B2(new_n883), .ZN(G367));
  XOR2_X1   g0684(.A(new_n634), .B(new_n636), .Z(new_n885));
  NAND2_X1  g0685(.A1(new_n683), .A2(KEYINPUT103), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT103), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n629), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n885), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n886), .A2(new_n885), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT44), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n596), .B1(new_n576), .B2(new_n652), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n608), .A2(new_n618), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n893), .B1(new_n637), .B2(new_n896), .ZN(new_n897));
  OR3_X1    g0697(.A1(new_n637), .A2(new_n893), .A3(new_n896), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT45), .B1(new_n637), .B2(new_n896), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n637), .A2(KEYINPUT45), .A3(new_n896), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n897), .A2(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(new_n635), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n681), .B1(new_n892), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n639), .B(KEYINPUT41), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n687), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT104), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n605), .A2(new_n652), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n606), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n473), .B2(new_n910), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n896), .A2(new_n634), .A3(new_n636), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT42), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n896), .A2(new_n630), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n618), .B1(new_n916), .B2(new_n583), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n913), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n918), .B(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n896), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n635), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n908), .A2(new_n909), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n923), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT104), .B1(new_n907), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n241), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n703), .B1(new_n209), .B2(new_n423), .C1(new_n928), .C2(new_n696), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n691), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT105), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n335), .B1(new_n719), .B2(new_n525), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n713), .A2(new_n501), .B1(new_n726), .B2(new_n738), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n932), .B(new_n933), .C1(G317), .C2(new_n716), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n732), .A2(KEYINPUT46), .A3(G116), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n730), .A2(G97), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT46), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n776), .B2(new_n480), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G283), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n723), .A2(new_n215), .B1(new_n709), .B2(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT106), .Z(new_n942));
  NOR2_X1   g0742(.A1(new_n719), .A2(new_n764), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n723), .A2(new_n273), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(G143), .C2(new_n725), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n292), .B1(new_n715), .B2(new_n765), .C1(new_n323), .C2(new_n709), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(G159), .B2(new_n712), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n732), .A2(G58), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n730), .A2(G77), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n947), .A2(new_n949), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n939), .A2(new_n942), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT47), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n702), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n953), .A2(new_n954), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n931), .B1(new_n956), .B2(new_n957), .C1(new_n912), .C2(new_n747), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n927), .A2(new_n958), .ZN(G387));
  NAND2_X1  g0759(.A1(new_n892), .A2(new_n680), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n886), .A2(new_n885), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(new_n889), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n681), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n639), .B(KEYINPUT111), .Z(new_n964));
  NAND3_X1  g0764(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n692), .A2(new_n640), .B1(G107), .B2(new_n209), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n238), .A2(G45), .ZN(new_n967));
  INV_X1    g0767(.A(new_n640), .ZN(new_n968));
  AOI211_X1 g0768(.A(G45), .B(new_n968), .C1(G68), .C2(G77), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n321), .A2(G50), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT50), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n696), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n966), .B1(new_n967), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n691), .B1(new_n973), .B2(new_n704), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT108), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n723), .A2(new_n423), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n323), .B2(new_n719), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT109), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n292), .B1(new_n715), .B2(new_n764), .C1(new_n273), .C2(new_n709), .ZN(new_n980));
  INV_X1    g0780(.A(G159), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n981), .A2(new_n726), .B1(new_n713), .B2(new_n321), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n732), .A2(G77), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n936), .A2(new_n983), .ZN(new_n984));
  NOR4_X1   g0784(.A1(new_n979), .A2(new_n980), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n732), .A2(G294), .B1(G283), .B2(new_n741), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n720), .A2(G317), .B1(new_n762), .B2(G303), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n725), .A2(G322), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n738), .C2(new_n713), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT48), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT110), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n990), .B2(new_n989), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT49), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n292), .B1(new_n716), .B2(G326), .ZN(new_n995));
  INV_X1    g0795(.A(new_n730), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n995), .B1(new_n996), .B2(new_n480), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n993), .B2(KEYINPUT49), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n985), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n975), .B1(new_n999), .B2(new_n706), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n634), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n701), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n962), .B2(new_n687), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n965), .A2(new_n1003), .ZN(G393));
  OR2_X1    g0804(.A1(new_n903), .A2(new_n688), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n703), .B1(new_n457), .B2(new_n209), .C1(new_n250), .C2(new_n696), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n335), .B1(new_n709), .B2(new_n501), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n713), .A2(new_n525), .B1(new_n480), .B2(new_n723), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(G322), .C2(new_n716), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G317), .A2(new_n725), .B1(new_n720), .B2(G311), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT52), .Z(new_n1011));
  NAND2_X1  g0811(.A1(new_n732), .A2(G283), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n731), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n292), .B1(new_n709), .B2(new_n321), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n723), .A2(new_n213), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(G50), .C2(new_n712), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n732), .A2(G68), .B1(G143), .B2(new_n716), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n775), .C1(KEYINPUT112), .C2(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n726), .A2(new_n764), .B1(new_n981), .B2(new_n719), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT51), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(KEYINPUT112), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1013), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT113), .Z(new_n1024));
  OAI211_X1 g0824(.A(new_n691), .B(new_n1006), .C1(new_n1024), .C2(new_n706), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT114), .Z(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n747), .B2(new_n896), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n963), .A2(new_n903), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n964), .B1(new_n963), .B2(new_n903), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1005), .B(new_n1027), .C1(new_n1029), .C2(new_n1030), .ZN(G390));
  NAND2_X1  g0831(.A1(new_n802), .A2(new_n836), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n855), .A2(new_n859), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n618), .B1(new_n649), .B2(new_n650), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n751), .A2(new_n434), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n750), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n801), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n836), .B(new_n874), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n867), .A2(new_n801), .A3(G330), .A4(new_n752), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(KEYINPUT115), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT115), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n678), .A2(new_n1041), .A3(new_n752), .A4(new_n801), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1033), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1039), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n855), .A2(new_n859), .A3(new_n699), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n691), .B1(new_n350), .B2(new_n759), .ZN(new_n1048));
  INV_X1    g0848(.A(G128), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n713), .A2(new_n765), .B1(new_n726), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G159), .B2(new_n741), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n730), .A2(G50), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(KEYINPUT54), .B(G143), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n335), .B1(new_n762), .B2(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n720), .A2(G132), .B1(new_n716), .B2(G125), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1051), .A2(new_n1052), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n732), .A2(G150), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT53), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1015), .B1(G283), .B2(new_n725), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n215), .B2(new_n713), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n719), .A2(new_n480), .B1(new_n715), .B2(new_n501), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n292), .B(new_n1062), .C1(G97), .C2(new_n762), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1063), .A2(new_n733), .A3(new_n768), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n1057), .A2(new_n1059), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1048), .B1(new_n1065), .B2(new_n702), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1046), .A2(new_n687), .B1(new_n1047), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n867), .A2(G330), .A3(new_n755), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n1037), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1040), .A2(new_n1042), .A3(new_n1036), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n801), .B1(new_n678), .B2(new_n752), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1039), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n794), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n678), .A2(new_n439), .ZN(new_n1075));
  AND4_X1   g0875(.A1(new_n348), .A2(new_n863), .A3(new_n595), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1044), .A2(new_n1045), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n964), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT117), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT116), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1045), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1033), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1082), .B1(new_n1085), .B2(new_n1077), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1082), .B(new_n1077), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1080), .B(new_n1081), .C1(new_n1086), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1077), .ZN(new_n1091));
  OAI21_X1  g0891(.A(KEYINPUT116), .B1(new_n1046), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n1087), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1081), .B1(new_n1093), .B2(new_n1080), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1067), .B1(new_n1090), .B2(new_n1094), .ZN(G378));
  XNOR2_X1  g0895(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n328), .A2(new_n822), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n349), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n349), .A2(new_n1098), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1101), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n1099), .A3(new_n1096), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n877), .A2(G330), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1105), .B1(new_n877), .B2(G330), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n862), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n877), .A2(G330), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1105), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1112), .A2(new_n861), .A3(new_n835), .A4(new_n1106), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1111), .A2(new_n699), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n691), .B1(G50), .B2(new_n759), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n331), .A2(new_n280), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT118), .ZN(new_n1118));
  AOI211_X1 g0918(.A(G50), .B(new_n1118), .C1(new_n280), .C2(new_n335), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n726), .A2(new_n480), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n944), .B(new_n1120), .C1(G97), .C2(new_n712), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n730), .A2(G58), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n280), .B(new_n335), .C1(new_n719), .C2(new_n215), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n709), .A2(new_n423), .B1(new_n715), .B2(new_n940), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1121), .A2(new_n983), .A3(new_n1122), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT58), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1119), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n719), .A2(new_n1049), .B1(new_n709), .B2(new_n765), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G132), .B2(new_n712), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G150), .A2(new_n741), .B1(new_n725), .B2(G125), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(new_n776), .C2(new_n1053), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(KEYINPUT59), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(KEYINPUT59), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n730), .A2(G159), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n716), .A2(G124), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .A4(new_n1118), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1128), .B1(new_n1127), .B2(new_n1126), .C1(new_n1133), .C2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1116), .B1(new_n1138), .B2(new_n702), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1114), .A2(new_n687), .B1(new_n1115), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT57), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT119), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1076), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1078), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1083), .A2(new_n1091), .A3(new_n1084), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT119), .B1(new_n1146), .B2(new_n1076), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1142), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n964), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1143), .B1(new_n1078), .B2(new_n1144), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1146), .A2(KEYINPUT119), .A3(new_n1076), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT57), .B1(new_n1152), .B2(new_n1114), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1140), .B1(new_n1149), .B2(new_n1153), .ZN(G375));
  OR2_X1    g0954(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n906), .A3(new_n1077), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT120), .Z(new_n1157));
  NAND2_X1  g0957(.A1(new_n1037), .A2(new_n699), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n691), .B1(G68), .B2(new_n759), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n977), .B1(new_n713), .B2(new_n480), .C1(new_n501), .C2(new_n726), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n732), .A2(G97), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n292), .B1(new_n720), .B2(G283), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G107), .A2(new_n762), .B1(new_n716), .B2(G303), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n951), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n732), .A2(G159), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n335), .B1(new_n762), .B2(G150), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n720), .A2(G137), .B1(new_n716), .B2(G128), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1122), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G132), .A2(new_n725), .B1(new_n712), .B2(new_n1054), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n323), .B2(new_n723), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n1160), .A2(new_n1164), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1159), .B1(new_n1171), .B2(new_n702), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1074), .A2(new_n687), .B1(new_n1158), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1157), .A2(new_n1173), .ZN(G381));
  INV_X1    g0974(.A(G396), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n965), .A2(new_n1003), .A3(new_n1175), .ZN(new_n1176));
  OR4_X1    g0976(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1080), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1067), .ZN(new_n1179));
  OR4_X1    g0979(.A1(G387), .A2(new_n1177), .A3(G375), .A4(new_n1179), .ZN(G407));
  INV_X1    g0980(.A(new_n1179), .ZN(new_n1181));
  INV_X1    g0981(.A(G213), .ZN(new_n1182));
  OR3_X1    g0982(.A1(new_n1182), .A2(KEYINPUT121), .A3(G343), .ZN(new_n1183));
  OAI21_X1  g0983(.A(KEYINPUT121), .B1(new_n1182), .B2(G343), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1181), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(G407), .B(G213), .C1(G375), .C2(new_n1187), .ZN(G409));
  INV_X1    g0988(.A(KEYINPUT61), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT60), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1155), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n964), .A3(new_n1077), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1155), .A2(new_n1190), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1173), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(G384), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(KEYINPUT123), .B2(new_n1185), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1186), .A2(G2897), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1196), .B(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1150), .A2(new_n1151), .B1(new_n1113), .B2(new_n1109), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1148), .B(new_n964), .C1(new_n1200), .C2(KEYINPUT57), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(G378), .A2(new_n1201), .A3(new_n1140), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1152), .A2(new_n906), .A3(new_n1114), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1140), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1181), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1186), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1189), .B1(new_n1199), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1005), .A2(new_n1027), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1030), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n1209), .B2(new_n1028), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1176), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1175), .B1(new_n965), .B2(new_n1003), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1210), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1212), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(G390), .A3(new_n1176), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(G387), .A2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n927), .A2(new_n1213), .A3(new_n1215), .A4(new_n958), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1067), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1178), .A2(KEYINPUT117), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1220), .B1(new_n1221), .B2(new_n1089), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1205), .B1(G375), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(new_n1185), .A3(new_n1195), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT63), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1219), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1207), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT122), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1224), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1206), .A2(KEYINPUT122), .A3(new_n1195), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n1225), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1227), .A2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1223), .A2(KEYINPUT62), .A3(new_n1185), .A4(new_n1195), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT124), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1206), .A2(KEYINPUT124), .A3(KEYINPUT62), .A4(new_n1195), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT62), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1229), .A2(new_n1238), .A3(new_n1230), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1207), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT125), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1232), .B1(new_n1240), .B2(new_n1242), .ZN(G405));
  NOR2_X1   g1043(.A1(G375), .A2(new_n1222), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1179), .B1(new_n1201), .B2(new_n1140), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1244), .A2(new_n1195), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1195), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G375), .A2(new_n1181), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1247), .B1(new_n1248), .B2(new_n1202), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1219), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1250), .A2(KEYINPUT127), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT127), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1195), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1248), .A2(new_n1202), .A3(new_n1247), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1252), .B1(new_n1255), .B2(new_n1219), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(new_n1241), .A3(new_n1254), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT126), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1251), .A2(new_n1256), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1250), .A2(KEYINPUT127), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1255), .A2(new_n1252), .A3(new_n1219), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1261), .A2(new_n1262), .B1(new_n1258), .B2(new_n1257), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1260), .A2(new_n1263), .ZN(G402));
endmodule


