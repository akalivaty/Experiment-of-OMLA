//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987;
  XOR2_X1   g000(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n202));
  OAI21_X1  g001(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g004(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n207), .A2(new_n208), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT66), .A3(KEYINPUT23), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT66), .B1(new_n215), .B2(KEYINPUT23), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n202), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT67), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n223), .A3(KEYINPUT23), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n208), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT68), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n213), .A2(KEYINPUT25), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n224), .A2(new_n230), .A3(new_n208), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n205), .A2(KEYINPUT69), .A3(new_n206), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT69), .B1(new_n205), .B2(new_n206), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n231), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n220), .B1(new_n229), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  INV_X1    g037(.A(G190gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n204), .B1(new_n240), .B2(KEYINPUT28), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n221), .A2(new_n223), .A3(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n244), .A2(new_n208), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G183gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT27), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT27), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G183gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n250), .A3(new_n239), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n241), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n236), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G134gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G127gat), .ZN(new_n258));
  INV_X1    g057(.A(G127gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G134gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G120gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(KEYINPUT1), .ZN(new_n263));
  INV_X1    g062(.A(G120gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G113gat), .ZN(new_n265));
  INV_X1    g064(.A(G113gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G120gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n274), .B(KEYINPUT64), .Z(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n227), .B1(new_n225), .B2(KEYINPUT68), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n207), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n232), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n231), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n254), .B1(new_n281), .B2(new_n220), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n263), .A2(new_n271), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n273), .A2(new_n276), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT34), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT34), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n273), .A2(new_n284), .A3(new_n287), .A4(new_n276), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G15gat), .B(G43gat), .Z(new_n290));
  XNOR2_X1  g089(.A(G71gat), .B(G99gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n256), .A2(new_n272), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n282), .A2(new_n283), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n275), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT33), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n276), .B1(new_n273), .B2(new_n284), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n292), .B1(new_n300), .B2(KEYINPUT33), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(new_n286), .A3(new_n288), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n304), .B2(new_n300), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n299), .A2(new_n302), .A3(KEYINPUT32), .A4(new_n296), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G228gat), .ZN(new_n308));
  INV_X1    g107(.A(G233gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G211gat), .ZN(new_n312));
  INV_X1    g111(.A(G218gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G211gat), .A2(G218gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n318), .A3(new_n315), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(G197gat), .A2(G204gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G197gat), .A2(G204gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT22), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n321), .A2(new_n322), .B1(new_n323), .B2(new_n315), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n317), .A2(new_n324), .A3(new_n319), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330));
  AND2_X1   g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT77), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n337));
  NAND2_X1  g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT78), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G141gat), .ZN(new_n344));
  INV_X1    g143(.A(G148gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347));
  NAND2_X1  g146(.A1(G141gat), .A2(G148gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n338), .A2(KEYINPUT2), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n343), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n340), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n350), .B1(new_n331), .B2(new_n332), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n346), .A2(new_n348), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n352), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n329), .B1(new_n330), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n353), .A2(new_n354), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(new_n340), .B2(new_n351), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n326), .A2(new_n330), .A3(new_n327), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(new_n356), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n311), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n360), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT85), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n343), .A2(new_n349), .A3(new_n350), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n333), .A2(new_n339), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n355), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n370), .B(new_n371), .C1(new_n360), .C2(new_n361), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n357), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT86), .B1(new_n374), .B2(KEYINPUT29), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n376), .A3(new_n330), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n328), .A3(new_n377), .ZN(new_n378));
  AND4_X1   g177(.A1(KEYINPUT87), .A2(new_n373), .A3(new_n378), .A4(new_n310), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n311), .B1(new_n366), .B2(new_n372), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT87), .B1(new_n380), .B2(new_n378), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n363), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G22gat), .ZN(new_n383));
  INV_X1    g182(.A(G22gat), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n384), .B(new_n363), .C1(new_n379), .C2(new_n381), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(KEYINPUT88), .A3(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(G78gat), .B(G106gat), .Z(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G50gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OR2_X1    g190(.A1(new_n379), .A2(new_n381), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT88), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n384), .A4(new_n363), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n386), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n383), .A2(KEYINPUT89), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n397), .A3(G22gat), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n396), .A2(new_n398), .A3(new_n390), .A4(new_n385), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n307), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT74), .ZN(new_n401));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT73), .B1(new_n282), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT73), .ZN(new_n404));
  INV_X1    g203(.A(new_n402), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n224), .A2(new_n208), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n406), .A2(new_n230), .B1(new_n279), .B2(new_n232), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n213), .A2(new_n208), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n408), .B(new_n207), .C1(new_n218), .C2(new_n217), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n407), .A2(new_n277), .B1(new_n409), .B2(new_n202), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n404), .B(new_n405), .C1(new_n410), .C2(new_n254), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n256), .A2(new_n330), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n403), .A2(new_n411), .B1(new_n412), .B2(new_n402), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n401), .B1(new_n413), .B2(new_n329), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n402), .B1(new_n282), .B2(KEYINPUT29), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n404), .B1(new_n256), .B2(new_n405), .ZN(new_n416));
  AOI211_X1 g215(.A(KEYINPUT73), .B(new_n402), .C1(new_n236), .C2(new_n255), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(KEYINPUT74), .A3(new_n328), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n282), .A2(new_n402), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n402), .B2(new_n412), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n329), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n414), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT76), .ZN(new_n424));
  XOR2_X1   g223(.A(G8gat), .B(G36gat), .Z(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT75), .ZN(new_n426));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  AND3_X1   g227(.A1(new_n423), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n424), .B1(new_n423), .B2(new_n428), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G225gat), .A2(G233gat), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n272), .B1(new_n360), .B2(new_n364), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n432), .B1(new_n433), .B2(new_n374), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(KEYINPUT5), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT82), .B1(new_n369), .B2(new_n272), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n360), .A2(new_n437), .A3(new_n283), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(KEYINPUT4), .A3(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n440));
  NAND3_X1  g239(.A1(new_n360), .A2(new_n283), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444));
  AOI211_X1 g243(.A(new_n444), .B(new_n440), .C1(new_n360), .C2(new_n283), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n283), .A2(new_n352), .A3(new_n355), .ZN(new_n446));
  INV_X1    g245(.A(new_n440), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT81), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT4), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n446), .A2(KEYINPUT82), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n437), .B1(new_n360), .B2(new_n283), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n434), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n369), .A2(new_n272), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n436), .A2(new_n438), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n432), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT5), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n443), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G1gat), .B(G29gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(KEYINPUT0), .ZN(new_n462));
  XNOR2_X1  g261(.A(G57gat), .B(G85gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n443), .B(new_n464), .C1(new_n454), .C2(new_n459), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n460), .A2(KEYINPUT6), .A3(new_n465), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n428), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n414), .A2(new_n419), .A3(new_n422), .A4(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT30), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n428), .A2(new_n474), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n414), .A2(new_n419), .A3(new_n422), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n471), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT83), .B1(new_n431), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n403), .A2(new_n411), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n329), .B1(new_n480), .B2(new_n415), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n422), .B1(new_n481), .B2(KEYINPUT74), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n413), .A2(new_n401), .A3(new_n329), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n428), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT76), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n423), .A2(new_n424), .A3(new_n428), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n414), .A2(new_n419), .A3(new_n422), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n470), .A2(new_n469), .B1(new_n489), .B2(new_n476), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n487), .A2(new_n488), .A3(new_n475), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n400), .A2(new_n479), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT35), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n475), .A2(new_n477), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n471), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n400), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n433), .A2(new_n374), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(new_n439), .B2(new_n441), .ZN(new_n503));
  OR3_X1    g302(.A1(new_n503), .A2(KEYINPUT39), .A3(new_n432), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n456), .A2(new_n457), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n505), .B(KEYINPUT39), .C1(new_n503), .C2(new_n432), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n464), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n509), .A2(KEYINPUT91), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(KEYINPUT91), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n507), .A2(new_n508), .B1(new_n460), .B2(new_n465), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT37), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n421), .B2(new_n328), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n418), .A2(new_n329), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n414), .A2(new_n419), .A3(new_n515), .A4(new_n422), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT92), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n428), .A4(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(new_n423), .B2(KEYINPUT37), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(new_n428), .A3(new_n521), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(new_n497), .A3(new_n473), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n395), .A2(new_n399), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n514), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n479), .A2(new_n491), .ZN(new_n532));
  INV_X1    g331(.A(new_n530), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT71), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n535), .A2(KEYINPUT71), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n307), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n305), .A2(KEYINPUT71), .A3(new_n535), .A4(new_n306), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT90), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n531), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n540), .B1(new_n532), .B2(new_n533), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT90), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n501), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G29gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT14), .B(G29gat), .Z(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(G36gat), .ZN(new_n551));
  INV_X1    g350(.A(G43gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(G50gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT94), .B(G50gat), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(new_n552), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n551), .B1(KEYINPUT15), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n552), .A2(G50gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(KEYINPUT15), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n559), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n551), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n563), .A2(KEYINPUT17), .ZN(new_n564));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565));
  INV_X1    g364(.A(G1gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT16), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n568), .B1(G1gat), .B2(new_n565), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G8gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n563), .A2(KEYINPUT17), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n564), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n563), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT95), .B1(new_n575), .B2(new_n570), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n571), .A2(new_n563), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n573), .B(new_n574), .C1(new_n576), .C2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT18), .ZN(new_n582));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G197gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT11), .B(G169gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  XOR2_X1   g385(.A(new_n586), .B(KEYINPUT12), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n576), .A2(new_n578), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n589), .B1(new_n575), .B2(new_n570), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n574), .B(KEYINPUT13), .Z(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT18), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n579), .A2(new_n580), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n582), .A2(new_n588), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT97), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n581), .A2(KEYINPUT18), .B1(new_n590), .B2(new_n591), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n597), .A2(new_n598), .A3(new_n588), .A4(new_n594), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n594), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n596), .A2(new_n599), .B1(new_n600), .B2(new_n587), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n547), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT98), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G71gat), .B(G78gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n605), .A2(new_n606), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n606), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(KEYINPUT99), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(new_n259), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n571), .B1(new_n613), .B2(new_n614), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(new_n334), .ZN(new_n622));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  OR2_X1    g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G85gat), .A2(G92gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT7), .ZN(new_n629));
  INV_X1    g428(.A(G99gat), .ZN(new_n630));
  INV_X1    g429(.A(G106gat), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT8), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT101), .B(G92gat), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n629), .B(new_n632), .C1(G85gat), .C2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G99gat), .B(G106gat), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n633), .A2(G85gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n635), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n637), .A2(new_n638), .A3(new_n629), .A4(new_n632), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n564), .A2(new_n572), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  AND2_X1   g441(.A1(G232gat), .A2(G233gat), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n575), .A2(new_n642), .B1(KEYINPUT41), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G190gat), .B(G218gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n643), .A2(KEYINPUT41), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT100), .ZN(new_n649));
  XNOR2_X1  g448(.A(G134gat), .B(G162gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n647), .A2(new_n652), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(G120gat), .B(G148gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT104), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n642), .A2(KEYINPUT10), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n613), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n609), .A2(new_n612), .A3(new_n640), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n636), .A2(new_n610), .A3(new_n639), .A4(new_n611), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(KEYINPUT102), .A3(new_n666), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n662), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(G230gat), .A2(G233gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT105), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n665), .A2(new_n672), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n660), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(KEYINPUT106), .B(new_n660), .C1(new_n674), .C2(new_n675), .ZN(new_n679));
  INV_X1    g478(.A(new_n672), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT103), .B1(new_n671), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT102), .B1(new_n665), .B2(new_n666), .ZN(new_n682));
  AOI211_X1 g481(.A(new_n668), .B(KEYINPUT10), .C1(new_n663), .C2(new_n664), .ZN(new_n683));
  OAI22_X1  g482(.A1(new_n682), .A2(new_n683), .B1(new_n613), .B2(new_n661), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n685), .A3(new_n672), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n675), .A2(new_n660), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n678), .A2(new_n679), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n627), .A2(new_n655), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n602), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n471), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n566), .ZN(G1324gat));
  NAND3_X1  g493(.A1(new_n602), .A2(new_n495), .A3(new_n691), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT16), .B(G8gat), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(G8gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n698), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(G1325gat));
  OAI21_X1  g501(.A(G15gat), .B1(new_n692), .B2(new_n541), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n307), .A2(G15gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n692), .B2(new_n704), .ZN(G1326gat));
  NAND3_X1  g504(.A1(new_n602), .A2(new_n533), .A3(new_n691), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT107), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT43), .B(G22gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  INV_X1    g508(.A(new_n627), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n689), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n655), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n602), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n548), .A3(new_n497), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT45), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n514), .A2(new_n529), .A3(new_n530), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n545), .A2(new_n718), .B1(new_n493), .B2(new_n499), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n719), .B2(new_n655), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n711), .A2(new_n601), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n655), .A2(new_n717), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n720), .B(new_n721), .C1(new_n547), .C2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n546), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n718), .B1(new_n545), .B2(KEYINPUT90), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n500), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n722), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n730), .A2(KEYINPUT108), .A3(new_n720), .A4(new_n721), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n726), .A2(new_n497), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n716), .B1(new_n548), .B2(new_n732), .ZN(G1328gat));
  INV_X1    g532(.A(G36gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n726), .A2(new_n495), .A3(new_n731), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n736), .B2(new_n735), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n713), .A2(G36gat), .A3(new_n496), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT46), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(G1329gat));
  NOR3_X1   g540(.A1(new_n713), .A2(G43gat), .A3(new_n307), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n540), .A3(new_n731), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(G43gat), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n724), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n552), .B1(new_n747), .B2(new_n540), .ZN(new_n748));
  OAI22_X1  g547(.A1(KEYINPUT47), .A2(new_n744), .B1(new_n746), .B2(new_n748), .ZN(G1330gat));
  NOR2_X1   g548(.A1(new_n530), .A2(new_n554), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n602), .A2(new_n712), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n554), .B1(new_n724), .B2(new_n530), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n752), .A2(KEYINPUT48), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n726), .A2(new_n533), .A3(new_n731), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n554), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n752), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n751), .B1(new_n756), .B2(new_n554), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n761), .A2(KEYINPUT110), .A3(KEYINPUT48), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n754), .B1(new_n760), .B2(new_n762), .ZN(G1331gat));
  INV_X1    g562(.A(new_n601), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n678), .A2(new_n679), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n687), .A2(new_n688), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n627), .A2(new_n655), .A3(new_n767), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n719), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n471), .B(KEYINPUT111), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g572(.A(new_n496), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n775), .B(new_n776), .Z(G1333gat));
  INV_X1    g576(.A(new_n307), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n769), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(G71gat), .B1(new_n779), .B2(KEYINPUT112), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(KEYINPUT112), .B2(new_n779), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n769), .A2(G71gat), .A3(new_n540), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n533), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g585(.A1(new_n730), .A2(new_n720), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n627), .A2(new_n764), .A3(new_n689), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n471), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n719), .A2(new_n655), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n627), .A2(new_n764), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n791), .A2(KEYINPUT51), .A3(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n689), .A2(G85gat), .A3(new_n471), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n790), .A2(new_n799), .ZN(G1336gat));
  NAND3_X1  g599(.A1(new_n787), .A2(new_n495), .A3(new_n788), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT113), .B1(new_n801), .B2(new_n633), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(KEYINPUT52), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n496), .A2(new_n689), .A3(G92gat), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n801), .A2(new_n633), .B1(new_n797), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n803), .B(new_n805), .ZN(G1337gat));
  OAI21_X1  g605(.A(G99gat), .B1(new_n789), .B2(new_n541), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n797), .A2(new_n630), .A3(new_n778), .A4(new_n767), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1338gat));
  OAI21_X1  g608(.A(G106gat), .B1(new_n789), .B2(new_n530), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n797), .A2(new_n631), .A3(new_n533), .A4(new_n767), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n812), .B(new_n815), .ZN(G1339gat));
  NAND2_X1  g615(.A1(new_n691), .A2(new_n601), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  INV_X1    g617(.A(new_n673), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT54), .B1(new_n684), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n681), .B2(new_n686), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n684), .A2(new_n819), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n660), .B1(new_n822), .B2(KEYINPUT54), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n818), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n671), .B2(new_n673), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n684), .A2(new_n685), .A3(new_n672), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n685), .B1(new_n684), .B2(new_n672), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n659), .B1(new_n674), .B2(new_n825), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(KEYINPUT55), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n824), .A2(new_n831), .A3(new_n766), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n596), .A2(new_n599), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n589), .A2(new_n573), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n834), .A2(new_n574), .B1(new_n590), .B2(new_n591), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n586), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n832), .A2(new_n837), .A3(new_n655), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n596), .A2(new_n599), .B1(new_n586), .B2(new_n835), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n767), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n840), .B1(new_n601), .B2(new_n832), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n838), .B1(new_n841), .B2(new_n655), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n817), .B1(new_n842), .B2(new_n627), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n771), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n844), .A2(new_n400), .A3(new_n496), .ZN(new_n845));
  AOI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n764), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n843), .A2(new_n530), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n495), .A2(new_n471), .A3(new_n307), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n601), .A2(new_n266), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT115), .ZN(G1340gat));
  AOI21_X1  g651(.A(G120gat), .B1(new_n845), .B2(new_n767), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n689), .A2(new_n264), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n849), .B2(new_n854), .ZN(G1341gat));
  INV_X1    g654(.A(new_n849), .ZN(new_n856));
  OAI21_X1  g655(.A(G127gat), .B1(new_n856), .B2(new_n710), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n845), .A2(new_n259), .A3(new_n627), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1342gat));
  INV_X1    g658(.A(new_n655), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n257), .A3(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n856), .B2(new_n655), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n533), .A2(KEYINPUT57), .ZN(new_n866));
  INV_X1    g665(.A(new_n838), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n837), .A2(new_n689), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n601), .B1(new_n832), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n824), .A2(new_n831), .A3(KEYINPUT116), .A4(new_n766), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n867), .B1(new_n872), .B2(new_n860), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n710), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n866), .B1(new_n874), .B2(new_n817), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n843), .A2(new_n533), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n690), .A2(new_n764), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n881), .B1(new_n873), .B2(new_n710), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT117), .B1(new_n882), .B2(new_n866), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n877), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n540), .A2(new_n471), .A3(new_n495), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n764), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n884), .A2(KEYINPUT118), .A3(new_n764), .A4(new_n885), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n888), .A2(G141gat), .A3(new_n889), .ZN(new_n890));
  AND4_X1   g689(.A1(new_n533), .A2(new_n844), .A3(new_n496), .A4(new_n541), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n344), .A3(new_n764), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n886), .A2(G141gat), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(new_n892), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n890), .A2(new_n894), .B1(new_n896), .B2(new_n893), .ZN(G1344gat));
  NOR2_X1   g696(.A1(new_n345), .A2(KEYINPUT59), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n884), .A2(new_n885), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n689), .ZN(new_n900));
  XNOR2_X1  g699(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n832), .A2(new_n869), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n764), .A3(new_n871), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n860), .B1(new_n903), .B2(new_n840), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT120), .B1(new_n904), .B2(new_n838), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n906), .B(new_n867), .C1(new_n872), .C2(new_n860), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n710), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n817), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n530), .A2(KEYINPUT57), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n911), .A2(new_n767), .A3(new_n885), .A4(new_n912), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT121), .B(new_n901), .C1(new_n913), .C2(G148gat), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n627), .B1(new_n873), .B2(KEYINPUT120), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n881), .B1(new_n916), .B2(new_n907), .ZN(new_n917));
  INV_X1    g716(.A(new_n910), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n767), .B(new_n912), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n885), .ZN(new_n920));
  OAI21_X1  g719(.A(G148gat), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n901), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n915), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n900), .B1(new_n914), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n891), .A2(new_n345), .A3(new_n767), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1345gat));
  OAI21_X1  g725(.A(G155gat), .B1(new_n899), .B2(new_n710), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n891), .A2(new_n334), .A3(new_n627), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1346gat));
  OAI21_X1  g728(.A(G162gat), .B1(new_n899), .B2(new_n655), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n891), .A2(new_n335), .A3(new_n860), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1347gat));
  AND2_X1   g731(.A1(new_n843), .A2(new_n471), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n933), .A2(new_n400), .A3(new_n495), .ZN(new_n934));
  AOI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n764), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n771), .A2(new_n496), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n847), .A2(new_n778), .A3(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(new_n209), .A3(new_n601), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT122), .ZN(G1348gat));
  AOI21_X1  g739(.A(G176gat), .B1(new_n934), .B2(new_n767), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT123), .Z(new_n942));
  NOR3_X1   g741(.A1(new_n937), .A2(new_n210), .A3(new_n689), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(G1349gat));
  OR3_X1    g743(.A1(new_n937), .A2(KEYINPUT124), .A3(new_n710), .ZN(new_n945));
  OAI21_X1  g744(.A(KEYINPUT124), .B1(new_n937), .B2(new_n710), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(G183gat), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n934), .A2(new_n238), .A3(new_n627), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g748(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1350gat));
  OAI21_X1  g753(.A(G190gat), .B1(new_n937), .B2(new_n655), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT61), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n934), .A2(new_n239), .A3(new_n860), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1351gat));
  NOR3_X1   g757(.A1(new_n540), .A2(new_n496), .A3(new_n530), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n933), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n764), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n911), .A2(new_n912), .ZN(new_n965));
  INV_X1    g764(.A(new_n936), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n966), .A2(new_n540), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n764), .A2(G197gat), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(G1352gat));
  NOR3_X1   g770(.A1(new_n960), .A2(G204gat), .A3(new_n689), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT62), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n919), .A2(new_n540), .A3(new_n966), .ZN(new_n974));
  INV_X1    g773(.A(G204gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(G1353gat));
  NAND3_X1  g775(.A1(new_n963), .A2(new_n312), .A3(new_n627), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n965), .A2(new_n627), .A3(new_n967), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n978), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  NOR3_X1   g781(.A1(new_n968), .A2(new_n313), .A3(new_n655), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n961), .A2(new_n860), .A3(new_n962), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n984), .A2(new_n985), .A3(new_n313), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(new_n984), .B2(new_n313), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n983), .A2(new_n986), .A3(new_n987), .ZN(G1355gat));
endmodule


