

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  NOR2_X1 U324 ( .A1(n433), .A2(n523), .ZN(n434) );
  XNOR2_X1 U325 ( .A(KEYINPUT101), .B(n463), .ZN(n549) );
  XOR2_X1 U326 ( .A(n333), .B(n332), .Z(n292) );
  XOR2_X1 U327 ( .A(n357), .B(n356), .Z(n293) );
  XNOR2_X1 U328 ( .A(n334), .B(n292), .ZN(n339) );
  XNOR2_X1 U329 ( .A(n404), .B(KEYINPUT47), .ZN(n405) );
  XNOR2_X1 U330 ( .A(n339), .B(n352), .ZN(n340) );
  XNOR2_X1 U331 ( .A(n406), .B(n405), .ZN(n411) );
  XOR2_X1 U332 ( .A(n355), .B(n341), .Z(n470) );
  NOR2_X1 U333 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U334 ( .A(n358), .B(n293), .ZN(n361) );
  AND2_X1 U335 ( .A1(n492), .A2(n476), .ZN(n477) );
  XNOR2_X1 U336 ( .A(n477), .B(KEYINPUT37), .ZN(n522) );
  XNOR2_X1 U337 ( .A(n366), .B(n365), .ZN(n584) );
  XOR2_X1 U338 ( .A(n453), .B(n452), .Z(n534) );
  XNOR2_X1 U339 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n480) );
  XNOR2_X1 U341 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XNOR2_X1 U342 ( .A(n481), .B(n480), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n295) );
  XNOR2_X1 U344 ( .A(G92GAT), .B(KEYINPUT77), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n308) );
  XOR2_X1 U346 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n297) );
  XNOR2_X1 U347 ( .A(G218GAT), .B(KEYINPUT81), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U349 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n299) );
  XNOR2_X1 U350 ( .A(G106GAT), .B(G162GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U352 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U353 ( .A(G134GAT), .B(KEYINPUT80), .Z(n424) );
  XOR2_X1 U354 ( .A(G99GAT), .B(G85GAT), .Z(n357) );
  XOR2_X1 U355 ( .A(G190GAT), .B(KEYINPUT82), .Z(n343) );
  XOR2_X1 U356 ( .A(n357), .B(n343), .Z(n303) );
  NAND2_X1 U357 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n424), .B(n304), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n315) );
  XOR2_X1 U362 ( .A(G29GAT), .B(G36GAT), .Z(n310) );
  XNOR2_X1 U363 ( .A(G50GAT), .B(G43GAT), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U365 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n312) );
  XNOR2_X1 U366 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n380) );
  XNOR2_X1 U369 ( .A(n315), .B(n380), .ZN(n489) );
  INV_X1 U370 ( .A(KEYINPUT74), .ZN(n316) );
  NAND2_X1 U371 ( .A1(n316), .A2(KEYINPUT75), .ZN(n319) );
  INV_X1 U372 ( .A(KEYINPUT75), .ZN(n317) );
  NAND2_X1 U373 ( .A1(n317), .A2(KEYINPUT74), .ZN(n318) );
  NAND2_X1 U374 ( .A1(n319), .A2(n318), .ZN(n321) );
  XNOR2_X1 U375 ( .A(G78GAT), .B(G148GAT), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n323) );
  XOR2_X1 U377 ( .A(G106GAT), .B(G204GAT), .Z(n322) );
  XOR2_X1 U378 ( .A(n323), .B(n322), .Z(n355) );
  XOR2_X1 U379 ( .A(G155GAT), .B(KEYINPUT3), .Z(n325) );
  XNOR2_X1 U380 ( .A(KEYINPUT94), .B(KEYINPUT2), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U382 ( .A(n326), .B(KEYINPUT95), .Z(n328) );
  XNOR2_X1 U383 ( .A(KEYINPUT93), .B(G162GAT), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n432) );
  XOR2_X1 U385 ( .A(G141GAT), .B(G22GAT), .Z(n371) );
  XOR2_X1 U386 ( .A(KEYINPUT96), .B(KEYINPUT24), .Z(n330) );
  NAND2_X1 U387 ( .A1(G228GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n371), .B(n331), .ZN(n334) );
  XOR2_X1 U390 ( .A(KEYINPUT91), .B(KEYINPUT23), .Z(n333) );
  XNOR2_X1 U391 ( .A(G50GAT), .B(KEYINPUT22), .ZN(n332) );
  INV_X1 U392 ( .A(G197GAT), .ZN(n338) );
  XOR2_X1 U393 ( .A(KEYINPUT92), .B(G218GAT), .Z(n336) );
  XNOR2_X1 U394 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n352) );
  XOR2_X1 U397 ( .A(n432), .B(n340), .Z(n341) );
  XNOR2_X1 U398 ( .A(G176GAT), .B(G92GAT), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n342), .B(G64GAT), .ZN(n359) );
  XOR2_X1 U400 ( .A(n359), .B(n343), .Z(n347) );
  XOR2_X1 U401 ( .A(G169GAT), .B(G8GAT), .Z(n374) );
  XOR2_X1 U402 ( .A(G183GAT), .B(KEYINPUT19), .Z(n345) );
  XNOR2_X1 U403 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n449) );
  XNOR2_X1 U405 ( .A(n374), .B(n449), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U407 ( .A(G204GAT), .B(KEYINPUT98), .Z(n349) );
  NAND2_X1 U408 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U410 ( .A(n351), .B(n350), .Z(n354) );
  XNOR2_X1 U411 ( .A(G36GAT), .B(n352), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n526) );
  INV_X1 U413 ( .A(KEYINPUT41), .ZN(n367) );
  XOR2_X1 U414 ( .A(G57GAT), .B(KEYINPUT13), .Z(n387) );
  XNOR2_X1 U415 ( .A(n355), .B(n387), .ZN(n358) );
  XOR2_X1 U416 ( .A(KEYINPUT76), .B(KEYINPUT33), .Z(n356) );
  XOR2_X1 U417 ( .A(G120GAT), .B(G71GAT), .Z(n439) );
  XNOR2_X1 U418 ( .A(n439), .B(n359), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n366) );
  XOR2_X1 U420 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n363) );
  NAND2_X1 U421 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U423 ( .A(KEYINPUT31), .B(n364), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n367), .B(n584), .ZN(n510) );
  XOR2_X1 U425 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n369) );
  XNOR2_X1 U426 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n379) );
  XNOR2_X1 U428 ( .A(G15GAT), .B(G1GAT), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n370), .B(KEYINPUT71), .ZN(n391) );
  XOR2_X1 U430 ( .A(n371), .B(n391), .Z(n373) );
  NAND2_X1 U431 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n373), .B(n372), .ZN(n375) );
  XOR2_X1 U433 ( .A(n375), .B(n374), .Z(n377) );
  XNOR2_X1 U434 ( .A(G113GAT), .B(G197GAT), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n581) );
  NOR2_X1 U438 ( .A1(n510), .A2(n581), .ZN(n383) );
  INV_X1 U439 ( .A(KEYINPUT46), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n403) );
  XOR2_X1 U441 ( .A(G71GAT), .B(G127GAT), .Z(n385) );
  XNOR2_X1 U442 ( .A(G22GAT), .B(G183GAT), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U444 ( .A(n387), .B(n386), .Z(n389) );
  NAND2_X1 U445 ( .A1(G231GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U447 ( .A(n390), .B(KEYINPUT15), .Z(n393) );
  XNOR2_X1 U448 ( .A(n391), .B(KEYINPUT12), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n401) );
  XOR2_X1 U450 ( .A(G211GAT), .B(G155GAT), .Z(n395) );
  XNOR2_X1 U451 ( .A(G8GAT), .B(G78GAT), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U453 ( .A(KEYINPUT14), .B(KEYINPUT83), .Z(n397) );
  XNOR2_X1 U454 ( .A(G64GAT), .B(KEYINPUT84), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U456 ( .A(n399), .B(n398), .Z(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n561) );
  INV_X1 U458 ( .A(n489), .ZN(n565) );
  NOR2_X1 U459 ( .A1(n561), .A2(n565), .ZN(n402) );
  NAND2_X1 U460 ( .A1(n403), .A2(n402), .ZN(n406) );
  XOR2_X1 U461 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n404) );
  XOR2_X1 U462 ( .A(KEYINPUT72), .B(n581), .Z(n568) );
  XNOR2_X1 U463 ( .A(KEYINPUT36), .B(n489), .ZN(n485) );
  INV_X1 U464 ( .A(n561), .ZN(n588) );
  NOR2_X1 U465 ( .A1(n485), .A2(n588), .ZN(n407) );
  XNOR2_X1 U466 ( .A(KEYINPUT45), .B(n407), .ZN(n408) );
  NAND2_X1 U467 ( .A1(n408), .A2(n584), .ZN(n409) );
  NOR2_X1 U468 ( .A1(n568), .A2(n409), .ZN(n410) );
  NOR2_X1 U469 ( .A1(n411), .A2(n410), .ZN(n412) );
  XOR2_X1 U470 ( .A(KEYINPUT48), .B(n412), .Z(n548) );
  NAND2_X1 U471 ( .A1(n526), .A2(n548), .ZN(n413) );
  XNOR2_X1 U472 ( .A(KEYINPUT54), .B(n413), .ZN(n433) );
  XOR2_X1 U473 ( .A(G85GAT), .B(G120GAT), .Z(n415) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(G141GAT), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U476 ( .A(KEYINPUT6), .B(G57GAT), .Z(n417) );
  XNOR2_X1 U477 ( .A(G1GAT), .B(G148GAT), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U479 ( .A(n419), .B(n418), .Z(n430) );
  XOR2_X1 U480 ( .A(KEYINPUT97), .B(KEYINPUT4), .Z(n421) );
  XNOR2_X1 U481 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n428) );
  XOR2_X1 U483 ( .A(G127GAT), .B(KEYINPUT0), .Z(n423) );
  XNOR2_X1 U484 ( .A(G113GAT), .B(KEYINPUT86), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n448) );
  XOR2_X1 U486 ( .A(n424), .B(n448), .Z(n426) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n523) );
  XNOR2_X1 U492 ( .A(n434), .B(KEYINPUT64), .ZN(n482) );
  NAND2_X1 U493 ( .A1(n470), .A2(n482), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n435), .B(KEYINPUT55), .ZN(n454) );
  XOR2_X1 U495 ( .A(G190GAT), .B(G134GAT), .Z(n437) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G99GAT), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U498 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n453) );
  XOR2_X1 U501 ( .A(KEYINPUT88), .B(KEYINPUT90), .Z(n443) );
  XNOR2_X1 U502 ( .A(G169GAT), .B(G176GAT), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U504 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n445) );
  XNOR2_X1 U505 ( .A(G15GAT), .B(KEYINPUT87), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U507 ( .A(n447), .B(n446), .Z(n451) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n452) );
  NAND2_X1 U510 ( .A1(n454), .A2(n534), .ZN(n572) );
  NOR2_X1 U511 ( .A1(n489), .A2(n572), .ZN(n458) );
  XNOR2_X1 U512 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n456) );
  INV_X1 U513 ( .A(G190GAT), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n568), .A2(n584), .ZN(n494) );
  NAND2_X1 U515 ( .A1(n534), .A2(n526), .ZN(n459) );
  NAND2_X1 U516 ( .A1(n459), .A2(n470), .ZN(n460) );
  XOR2_X1 U517 ( .A(KEYINPUT25), .B(n460), .Z(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(KEYINPUT102), .ZN(n465) );
  XNOR2_X1 U519 ( .A(n526), .B(KEYINPUT27), .ZN(n468) );
  NOR2_X1 U520 ( .A1(n534), .A2(n470), .ZN(n462) );
  XOR2_X1 U521 ( .A(KEYINPUT26), .B(n462), .Z(n463) );
  NAND2_X1 U522 ( .A1(n468), .A2(n549), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U524 ( .A(KEYINPUT103), .B(n466), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n523), .A2(n467), .ZN(n474) );
  NAND2_X1 U526 ( .A1(n468), .A2(n523), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n469), .B(KEYINPUT99), .ZN(n550) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT28), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT66), .ZN(n501) );
  NAND2_X1 U530 ( .A1(n550), .A2(n501), .ZN(n536) );
  NOR2_X1 U531 ( .A1(n534), .A2(n536), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT100), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT104), .B(n475), .Z(n492) );
  NOR2_X1 U534 ( .A1(n561), .A2(n485), .ZN(n476) );
  OR2_X1 U535 ( .A1(n494), .A2(n522), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT107), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT38), .B(n479), .ZN(n508) );
  NAND2_X1 U538 ( .A1(n508), .A2(n534), .ZN(n481) );
  NAND2_X1 U539 ( .A1(n549), .A2(n482), .ZN(n484) );
  INV_X1 U540 ( .A(KEYINPUT125), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n587) );
  NOR2_X1 U542 ( .A1(n485), .A2(n587), .ZN(n486) );
  XNOR2_X1 U543 ( .A(KEYINPUT62), .B(n486), .ZN(n488) );
  INV_X1 U544 ( .A(G218GAT), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n488), .B(n487), .ZN(G1355GAT) );
  NAND2_X1 U546 ( .A1(n561), .A2(n489), .ZN(n490) );
  XNOR2_X1 U547 ( .A(n490), .B(KEYINPUT85), .ZN(n491) );
  XNOR2_X1 U548 ( .A(KEYINPUT16), .B(n491), .ZN(n493) );
  NAND2_X1 U549 ( .A1(n493), .A2(n492), .ZN(n511) );
  NOR2_X1 U550 ( .A1(n494), .A2(n511), .ZN(n502) );
  NAND2_X1 U551 ( .A1(n523), .A2(n502), .ZN(n495) );
  XNOR2_X1 U552 ( .A(n495), .B(KEYINPUT34), .ZN(n496) );
  XNOR2_X1 U553 ( .A(G1GAT), .B(n496), .ZN(G1324GAT) );
  NAND2_X1 U554 ( .A1(n502), .A2(n526), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n497), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT105), .B(KEYINPUT35), .Z(n499) );
  NAND2_X1 U557 ( .A1(n502), .A2(n534), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U559 ( .A(G15GAT), .B(n500), .Z(G1326GAT) );
  INV_X1 U560 ( .A(n501), .ZN(n531) );
  NAND2_X1 U561 ( .A1(n531), .A2(n502), .ZN(n503) );
  XNOR2_X1 U562 ( .A(n503), .B(KEYINPUT106), .ZN(n504) );
  XNOR2_X1 U563 ( .A(G22GAT), .B(n504), .ZN(G1327GAT) );
  XOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT39), .Z(n506) );
  NAND2_X1 U565 ( .A1(n508), .A2(n523), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NAND2_X1 U567 ( .A1(n508), .A2(n526), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n507), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U569 ( .A1(n508), .A2(n531), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U571 ( .A(n510), .ZN(n557) );
  NAND2_X1 U572 ( .A1(n581), .A2(n557), .ZN(n521) );
  NOR2_X1 U573 ( .A1(n521), .A2(n511), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n523), .A2(n518), .ZN(n514) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(KEYINPUT42), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  XOR2_X1 U578 ( .A(G64GAT), .B(KEYINPUT109), .Z(n516) );
  NAND2_X1 U579 ( .A1(n518), .A2(n526), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n518), .A2(n534), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U584 ( .A1(n518), .A2(n531), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n525) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n530), .A2(n523), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  XOR2_X1 U590 ( .A(G92GAT), .B(KEYINPUT111), .Z(n528) );
  NAND2_X1 U591 ( .A1(n530), .A2(n526), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n530), .A2(n534), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n532), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NAND2_X1 U598 ( .A1(n534), .A2(n548), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n568), .A2(n545), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n539) );
  NAND2_X1 U603 ( .A1(n545), .A2(n557), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n540), .ZN(G1341GAT) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n544) );
  XOR2_X1 U607 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n542) );
  NAND2_X1 U608 ( .A1(n545), .A2(n561), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U612 ( .A1(n545), .A2(n565), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  INV_X1 U614 ( .A(n548), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U617 ( .A(KEYINPUT117), .B(n553), .Z(n564) );
  INV_X1 U618 ( .A(n581), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n564), .A2(n554), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT118), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  NAND2_X1 U623 ( .A1(n564), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  XOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT119), .Z(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1346GAT) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(KEYINPUT120), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n567), .B(n566), .ZN(G1347GAT) );
  INV_X1 U632 ( .A(n568), .ZN(n569) );
  NOR2_X1 U633 ( .A1(n569), .A2(n572), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n570), .B(KEYINPUT121), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n571), .B(G169GAT), .ZN(G1348GAT) );
  NOR2_X1 U636 ( .A1(n572), .A2(n510), .ZN(n577) );
  XOR2_X1 U637 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n574) );
  XNOR2_X1 U638 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT56), .B(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1349GAT) );
  NOR2_X1 U642 ( .A1(n588), .A2(n572), .ZN(n578) );
  XOR2_X1 U643 ( .A(G183GAT), .B(n578), .Z(G1350GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n583) );
  NOR2_X1 U647 ( .A1(n581), .A2(n587), .ZN(n582) );
  XOR2_X1 U648 ( .A(n583), .B(n582), .Z(G1352GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n587), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(G1354GAT) );
endmodule

