//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT68), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n453), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT72), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n463), .A2(KEYINPUT72), .A3(G101), .A4(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT71), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n470), .B2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(G2104), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n471), .A2(new_n473), .A3(new_n463), .A4(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n468), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n474), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n483));
  INV_X1    g058(.A(G125), .ZN(new_n484));
  NOR3_X1   g059(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT69), .B1(new_n486), .B2(G125), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n480), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n477), .B1(new_n488), .B2(G2105), .ZN(G160));
  NAND4_X1  g064(.A1(new_n471), .A2(new_n473), .A3(G2105), .A4(new_n474), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n463), .A2(G112), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n493));
  OAI22_X1  g068(.A1(new_n490), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n475), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(G136), .B2(new_n495), .ZN(G162));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n471), .A2(new_n473), .A3(new_n498), .A4(new_n474), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n497), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n499), .A2(KEYINPUT4), .B1(new_n486), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G126), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n463), .A2(G114), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  OAI22_X1  g079(.A1(new_n490), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n501), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(G75), .A2(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(G651), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT73), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n518), .A2(G50), .A3(G543), .A4(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n508), .A2(new_n509), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n512), .B(new_n520), .C1(new_n521), .C2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  INV_X1    g100(.A(new_n523), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n518), .A2(G543), .A3(new_n519), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n522), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n527), .A2(new_n530), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n538), .A2(new_n528), .B1(new_n523), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT74), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n514), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(new_n526), .A2(G81), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n514), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n529), .A2(G43), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g127(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  AOI22_X1  g131(.A1(new_n522), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(KEYINPUT76), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n514), .B1(new_n557), .B2(KEYINPUT76), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n558), .A2(new_n559), .B1(G91), .B2(new_n526), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n518), .A2(G53), .A3(G543), .A4(new_n519), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(G299));
  NAND2_X1  g138(.A1(new_n541), .A2(new_n543), .ZN(G301));
  NAND4_X1  g139(.A1(new_n518), .A2(G49), .A3(G543), .A4(new_n519), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n566));
  INV_X1    g141(.A(G87), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n565), .B(new_n566), .C1(new_n523), .C2(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT77), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G288));
  NAND4_X1  g145(.A1(new_n518), .A2(G86), .A3(new_n522), .A4(new_n519), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n518), .A2(G48), .A3(G543), .A4(new_n519), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n574));
  INV_X1    g149(.A(new_n509), .ZN(new_n575));
  NOR2_X1   g150(.A1(KEYINPUT5), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G61), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n574), .B1(new_n579), .B2(G651), .ZN(new_n580));
  AOI211_X1 g155(.A(KEYINPUT78), .B(new_n514), .C1(new_n577), .C2(new_n578), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n573), .B1(new_n580), .B2(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n514), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT79), .ZN(new_n585));
  AOI22_X1  g160(.A1(G47), .A2(new_n529), .B1(new_n526), .B2(G85), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G290));
  INV_X1    g162(.A(G92), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n523), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(new_n522), .ZN(new_n592));
  XNOR2_X1  g167(.A(KEYINPUT80), .B(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n529), .A2(G54), .B1(new_n594), .B2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT81), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n590), .A2(new_n598), .A3(new_n595), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  MUX2_X1   g177(.A(G301), .B(new_n601), .S(new_n602), .Z(G284));
  MUX2_X1   g178(.A(G301), .B(new_n601), .S(new_n602), .Z(G321));
  NAND2_X1  g179(.A1(G299), .A2(new_n602), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n602), .B2(G168), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n602), .B2(G168), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n600), .B1(new_n608), .B2(G860), .ZN(G148));
  OAI21_X1  g184(.A(KEYINPUT82), .B1(new_n550), .B2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n600), .A2(new_n608), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  MUX2_X1   g187(.A(KEYINPUT82), .B(new_n610), .S(new_n612), .Z(G323));
  XOR2_X1   g188(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n614));
  XNOR2_X1  g189(.A(G323), .B(new_n614), .ZN(G282));
  NOR2_X1   g190(.A1(new_n472), .A2(G2105), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n486), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  OR2_X1    g195(.A1(G99), .A2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n621), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n490), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(G135), .B2(new_n495), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(G2096), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n620), .A2(new_n627), .A3(new_n628), .ZN(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n642), .A2(G14), .A3(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT17), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT84), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n648), .B2(new_n645), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n650), .B2(new_n652), .ZN(new_n654));
  INV_X1    g229(.A(new_n645), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n651), .A3(new_n647), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n646), .A2(new_n651), .A3(new_n648), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n667), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n669), .B(new_n672), .C1(new_n664), .C2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G23), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n568), .B(KEYINPUT86), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT33), .B(G1976), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n684), .B(new_n685), .Z(new_n686));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n681), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n681), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT88), .Z(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(G1971), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n681), .A2(G6), .ZN(new_n693));
  INV_X1    g268(.A(G305), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(new_n681), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT32), .B(G1981), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n691), .A2(G1971), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n692), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n686), .A2(new_n687), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n688), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT34), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  MUX2_X1   g279(.A(G24), .B(G290), .S(G16), .Z(new_n705));
  INV_X1    g280(.A(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G25), .ZN(new_n709));
  OR2_X1    g284(.A1(G95), .A2(G2105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n710), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n711));
  INV_X1    g286(.A(G119), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n490), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G131), .B2(new_n495), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n709), .B1(new_n714), .B2(new_n708), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n703), .A2(new_n704), .A3(new_n707), .A4(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G4), .A2(G16), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n600), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT89), .B(G1348), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n681), .A2(G19), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT90), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n550), .B2(new_n681), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1341), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n708), .A2(G27), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G164), .B2(new_n708), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2078), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G11), .ZN(new_n732));
  INV_X1    g307(.A(G28), .ZN(new_n733));
  AOI21_X1  g308(.A(G29), .B1(new_n733), .B2(KEYINPUT30), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(KEYINPUT94), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(KEYINPUT94), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(KEYINPUT30), .B2(new_n733), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n732), .B1(new_n735), .B2(new_n737), .C1(new_n626), .C2(new_n708), .ZN(new_n738));
  INV_X1    g313(.A(G2072), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n708), .A2(G33), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT25), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G139), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OAI221_X1 g320(.A(new_n743), .B1(new_n475), .B2(new_n744), .C1(new_n745), .C2(new_n463), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n740), .B1(new_n746), .B2(G29), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n738), .B1(new_n739), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n739), .B2(new_n747), .ZN(new_n749));
  NOR4_X1   g324(.A1(new_n724), .A2(new_n728), .A3(new_n731), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n708), .A2(G26), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n495), .A2(G140), .ZN(new_n754));
  INV_X1    g329(.A(new_n490), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G128), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n463), .A2(G116), .ZN(new_n757));
  OAI21_X1  g332(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n754), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT91), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n753), .B1(new_n760), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2067), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n750), .B(new_n762), .C1(new_n722), .C2(new_n723), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT26), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n766), .A2(new_n767), .B1(G105), .B2(new_n616), .ZN(new_n768));
  INV_X1    g343(.A(G129), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n490), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G141), .B2(new_n495), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT93), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(new_n708), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n708), .B2(G32), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n681), .A2(G5), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G171), .B2(new_n681), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n774), .A2(new_n775), .B1(G1961), .B2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2090), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n708), .A2(G35), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT95), .Z(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G162), .B2(new_n708), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT29), .Z(new_n783));
  OAI221_X1 g358(.A(new_n778), .B1(new_n779), .B2(new_n783), .C1(new_n775), .C2(new_n774), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n681), .A2(G21), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G168), .B2(new_n681), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n786), .A2(G1966), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(G1966), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT24), .ZN(new_n789));
  INV_X1    g364(.A(G34), .ZN(new_n790));
  AOI21_X1  g365(.A(G29), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G160), .B2(new_n708), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G2084), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n788), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n787), .B(new_n796), .C1(new_n795), .C2(new_n794), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n681), .A2(G20), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT23), .Z(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G299), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1956), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n777), .A2(G1961), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n783), .A2(new_n779), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n797), .A2(new_n801), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n720), .A2(new_n763), .A3(new_n784), .A4(new_n804), .ZN(G311));
  OR4_X1    g380(.A1(new_n720), .A2(new_n763), .A3(new_n784), .A4(new_n804), .ZN(G150));
  NAND2_X1  g381(.A1(new_n600), .A2(G559), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT38), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n526), .A2(G93), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT96), .B(G55), .Z(new_n811));
  OAI221_X1 g386(.A(new_n809), .B1(new_n514), .B2(new_n810), .C1(new_n528), .C2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n550), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n808), .B(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n816), .A2(new_n817), .A3(G860), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n812), .A2(G860), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n820));
  XOR2_X1   g395(.A(new_n819), .B(new_n820), .Z(new_n821));
  OR2_X1    g396(.A1(new_n818), .A2(new_n821), .ZN(G145));
  NAND2_X1  g397(.A1(new_n495), .A2(G142), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n755), .A2(G130), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n825));
  INV_X1    g400(.A(G118), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n825), .A2(KEYINPUT99), .B1(new_n826), .B2(G2105), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(KEYINPUT99), .B2(new_n825), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n823), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(new_n618), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n714), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n486), .A2(new_n500), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n501), .A2(KEYINPUT98), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n505), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n760), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n771), .A2(new_n746), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n772), .B2(new_n746), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n840), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n832), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n831), .B(KEYINPUT100), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(new_n843), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n626), .B(G160), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G162), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(G37), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n847), .A2(new_n843), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n850), .B1(new_n854), .B2(new_n848), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g432(.A1(new_n812), .A2(new_n602), .ZN(new_n858));
  XNOR2_X1  g433(.A(G290), .B(new_n694), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n683), .B(G166), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT103), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT42), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n865));
  INV_X1    g440(.A(new_n861), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n864), .B(new_n865), .C1(KEYINPUT42), .C2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n865), .B2(new_n864), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n596), .A2(G299), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n596), .A2(G299), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT41), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n611), .B(new_n813), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n871), .B(KEYINPUT102), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n868), .B(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n858), .B1(new_n878), .B2(new_n602), .ZN(G295));
  OAI21_X1  g454(.A(new_n858), .B1(new_n878), .B2(new_n602), .ZN(G331));
  NAND2_X1  g455(.A1(G171), .A2(G168), .ZN(new_n881));
  NAND2_X1  g456(.A1(G301), .A2(G286), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n814), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n813), .A3(new_n882), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(KEYINPUT106), .A3(new_n885), .ZN(new_n886));
  OR3_X1    g461(.A1(new_n883), .A2(KEYINPUT106), .A3(new_n814), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n870), .A3(new_n869), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n885), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n872), .A2(new_n890), .A3(KEYINPUT105), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n884), .A2(new_n885), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n873), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n889), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n863), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT107), .B1(new_n897), .B2(G37), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n895), .A2(new_n896), .ZN(new_n899));
  AOI21_X1  g474(.A(G37), .B1(new_n895), .B2(new_n896), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT43), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n899), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n893), .A2(new_n876), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT108), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n888), .A2(new_n873), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n896), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AND4_X1   g483(.A1(KEYINPUT43), .A2(new_n904), .A3(new_n853), .A4(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT44), .B1(new_n903), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(new_n898), .B2(new_n902), .ZN(new_n913));
  AND4_X1   g488(.A1(new_n912), .A2(new_n904), .A3(new_n853), .A4(new_n908), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n915), .ZN(G397));
  XOR2_X1   g491(.A(new_n760), .B(G2067), .Z(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n771), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n503), .A2(new_n504), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n919), .B1(new_n755), .B2(G126), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n833), .A2(KEYINPUT98), .A3(new_n834), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT98), .B1(new_n833), .B2(new_n834), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G1384), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n925), .A2(KEYINPUT109), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(KEYINPUT109), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n477), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n483), .B1(new_n482), .B2(new_n484), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n486), .A2(KEYINPUT69), .A3(G125), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n479), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n930), .B(G40), .C1(new_n933), .C2(new_n463), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n918), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT127), .Z(new_n937));
  INV_X1    g512(.A(G1996), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n939), .B(KEYINPUT46), .Z(new_n940));
  NOR2_X1   g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT47), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n772), .A2(new_n938), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n917), .B(new_n943), .C1(new_n938), .C2(new_n771), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n714), .A2(new_n716), .ZN(new_n945));
  OAI22_X1  g520(.A1(new_n944), .A2(new_n945), .B1(G2067), .B2(new_n760), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n935), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n714), .B(new_n716), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n935), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n935), .A2(new_n706), .A3(new_n585), .A4(new_n586), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n952));
  OAI22_X1  g527(.A1(new_n949), .A2(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n947), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n942), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G8), .ZN(new_n957));
  NOR2_X1   g532(.A1(G168), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n925), .A2(new_n927), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n927), .A2(G1384), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(G164), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(KEYINPUT116), .B(new_n962), .C1(new_n501), .C2(new_n505), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n934), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(G1966), .B1(new_n960), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G40), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n968), .B(new_n477), .C1(new_n488), .C2(G2105), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n795), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n839), .B2(G1384), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n920), .A2(new_n835), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(KEYINPUT50), .A3(new_n924), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n970), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT119), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1966), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT116), .B1(new_n973), .B2(new_n962), .ZN(new_n978));
  INV_X1    g553(.A(new_n965), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n969), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT45), .B1(new_n923), .B2(new_n924), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT50), .B1(new_n923), .B2(new_n924), .ZN(new_n983));
  INV_X1    g558(.A(new_n974), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n795), .B(new_n969), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT119), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n982), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n959), .B1(new_n976), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n967), .A2(new_n975), .A3(KEYINPUT119), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n986), .B1(new_n982), .B2(new_n985), .ZN(new_n992));
  OAI21_X1  g567(.A(G8), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT120), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n958), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n957), .B1(new_n976), .B2(new_n987), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT120), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n990), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(G8), .B1(new_n967), .B2(new_n975), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(new_n990), .A3(new_n959), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n989), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1976), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT52), .B1(G288), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n839), .A2(G1384), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n957), .B1(new_n1005), .B2(new_n969), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n683), .A2(G1976), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1007), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n969), .A2(new_n924), .A3(new_n923), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G8), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT52), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1981), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n579), .A2(G651), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n573), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT111), .B1(G305), .B2(G1981), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n580), .A2(new_n581), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n1013), .A4(new_n573), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1015), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1006), .B1(new_n1020), .B2(KEYINPUT49), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n1022), .B(new_n1015), .C1(new_n1016), .C2(new_n1019), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1008), .B(new_n1012), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n925), .A2(KEYINPUT50), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n924), .B1(new_n501), .B2(new_n505), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1028), .B2(KEYINPUT50), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n973), .A2(KEYINPUT114), .A3(new_n971), .A4(new_n924), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1026), .A2(new_n779), .A3(new_n969), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n923), .A2(new_n962), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1028), .A2(new_n927), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n969), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1971), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G8), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G303), .A2(G8), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1039), .A2(KEYINPUT115), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n957), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1044), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n779), .B(new_n969), .C1(new_n983), .C2(new_n984), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1037), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1044), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1042), .A2(KEYINPUT110), .A3(new_n1043), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1051), .A2(G8), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1025), .A2(new_n1046), .A3(new_n1049), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT124), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1059));
  AOI211_X1 g634(.A(new_n957), .B(new_n1059), .C1(new_n1037), .C2(new_n1050), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(new_n1024), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1061), .A2(KEYINPUT124), .A3(new_n1049), .A4(new_n1046), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(G2078), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n960), .A2(new_n966), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n969), .B1(new_n983), .B2(new_n984), .ZN(new_n1068));
  INV_X1    g643(.A(G1961), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G2078), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1033), .A2(new_n1071), .A3(new_n969), .A4(new_n1034), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1072), .A2(KEYINPUT121), .A3(new_n1065), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT121), .B1(new_n1072), .B2(new_n1065), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1067), .B(new_n1070), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G171), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n930), .A2(G40), .A3(new_n1066), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n488), .A2(KEYINPUT123), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n463), .B1(new_n488), .B2(KEYINPUT123), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n929), .A2(new_n1033), .A3(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n1070), .C1(new_n1074), .C2(new_n1073), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(G171), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1064), .B1(new_n1080), .B2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT58), .B(G1341), .Z(new_n1089));
  NAND2_X1  g664(.A1(new_n1010), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1035), .B2(G1996), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n550), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT59), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1094), .A3(new_n550), .ZN(new_n1095));
  INV_X1    g670(.A(G1348), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1068), .A2(new_n1096), .ZN(new_n1097));
  OR3_X1    g672(.A1(new_n1010), .A2(KEYINPUT118), .A3(G2067), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT118), .B1(new_n1010), .B2(G2067), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n597), .A2(new_n1100), .A3(new_n599), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n601), .A2(new_n1100), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1093), .A2(new_n1095), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n562), .B2(KEYINPUT117), .ZN(new_n1106));
  XNOR2_X1  g681(.A(G299), .B(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n934), .B1(new_n925), .B2(KEYINPUT50), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1956), .B1(new_n1109), .B2(new_n1031), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1033), .A2(new_n969), .A3(new_n1034), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1108), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1026), .A2(new_n969), .A3(new_n1031), .ZN(new_n1115));
  INV_X1    g690(.A(G1956), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1107), .B1(new_n1117), .B2(new_n1112), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1105), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1108), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT61), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1104), .A2(new_n1119), .A3(new_n1120), .A4(new_n1123), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n601), .B1(new_n1125), .B2(new_n1097), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1122), .B1(new_n1126), .B2(new_n1118), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1075), .B2(G171), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1070), .A2(new_n1067), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1130), .A2(KEYINPUT125), .A3(G301), .A4(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1064), .B1(new_n1086), .B2(G171), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1124), .A2(new_n1127), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1002), .A2(new_n1063), .A3(new_n1088), .A4(new_n1135), .ZN(new_n1136));
  OR3_X1    g711(.A1(new_n1024), .A2(G286), .A3(new_n999), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1044), .B1(new_n1051), .B2(G8), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT63), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1025), .A2(new_n1060), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n569), .A2(new_n1003), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(KEYINPUT112), .Z(new_n1143));
  NOR2_X1   g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1016), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1019), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT113), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT113), .ZN(new_n1149));
  OAI221_X1 g724(.A(new_n1149), .B1(new_n1145), .B2(new_n1146), .C1(new_n1141), .C2(new_n1143), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1006), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1139), .A2(new_n1140), .A3(new_n1151), .ZN(new_n1152));
  NOR4_X1   g727(.A1(new_n1056), .A2(KEYINPUT63), .A3(G286), .A4(new_n999), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1058), .A2(new_n1080), .A3(new_n1062), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n959), .B1(new_n996), .B2(KEYINPUT120), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n994), .B(new_n957), .C1(new_n976), .C2(new_n987), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT51), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n988), .B1(new_n1158), .B2(new_n1000), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1155), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g736(.A(KEYINPUT62), .B(new_n988), .C1(new_n1158), .C2(new_n1000), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1136), .B(new_n1154), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n1164));
  XNOR2_X1  g739(.A(G290), .B(new_n706), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n949), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n935), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1163), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1164), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n956), .B1(new_n1168), .B2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g745(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1172));
  OAI211_X1 g746(.A(new_n856), .B(new_n1172), .C1(new_n913), .C2(new_n914), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


