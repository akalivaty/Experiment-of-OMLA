//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G128), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n190), .A2(new_n191), .A3(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT64), .B1(new_n198), .B2(new_n189), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(KEYINPUT0), .A3(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n203));
  AND4_X1   g017(.A1(new_n203), .A2(new_n193), .A3(new_n195), .A4(G128), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g021(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n194), .C2(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(G128), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n204), .B1(new_n209), .B2(new_n196), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n202), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G224), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G953), .ZN(new_n215));
  XOR2_X1   g029(.A(new_n213), .B(new_n215), .Z(new_n216));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n217));
  INV_X1    g031(.A(G116), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G119), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT68), .A3(G116), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(G119), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT5), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n220), .A3(G116), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G113), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT2), .B(G113), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n230), .A2(new_n219), .A3(new_n221), .A4(new_n222), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n232));
  INV_X1    g046(.A(G107), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(G104), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT77), .A2(G107), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT77), .A2(G107), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(G104), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n234), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G104), .ZN(new_n241));
  AOI21_X1  g055(.A(G101), .B1(new_n241), .B2(G107), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n235), .B2(new_n236), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n233), .A2(G104), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n240), .A2(new_n242), .B1(new_n245), .B2(G101), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n228), .A2(new_n231), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G110), .B(G122), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n241), .A2(G107), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT77), .B(G107), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n238), .ZN(new_n254));
  INV_X1    g068(.A(G101), .ZN(new_n255));
  OR2_X1    g069(.A1(KEYINPUT78), .A2(KEYINPUT4), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT78), .A2(KEYINPUT4), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n254), .A2(KEYINPUT79), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT79), .B1(new_n254), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n223), .A2(new_n229), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n231), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n255), .B1(new_n240), .B2(new_n251), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n252), .B(new_n242), .C1(new_n253), .C2(new_n238), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT4), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n250), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n254), .A2(new_n258), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT79), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n254), .A2(KEYINPUT79), .A3(new_n258), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n274), .B1(new_n240), .B2(new_n242), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n254), .A2(G101), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n275), .A2(new_n276), .B1(new_n262), .B2(new_n231), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n273), .A2(new_n277), .A3(KEYINPUT84), .ZN(new_n278));
  AOI211_X1 g092(.A(new_n247), .B(new_n249), .C1(new_n268), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n247), .B1(new_n268), .B2(new_n278), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT85), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n248), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OAI22_X1  g098(.A1(new_n279), .A2(new_n280), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n268), .A2(new_n278), .ZN(new_n286));
  INV_X1    g100(.A(new_n247), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT6), .A3(new_n283), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n216), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n213), .A2(new_n292), .A3(new_n215), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n215), .A2(new_n292), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n212), .B2(new_n202), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n246), .B1(new_n228), .B2(new_n231), .ZN(new_n297));
  INV_X1    g111(.A(new_n225), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT86), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n227), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n299), .B2(new_n298), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n246), .A2(new_n231), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n297), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  XOR2_X1   g117(.A(new_n248), .B(KEYINPUT8), .Z(new_n304));
  OAI21_X1  g118(.A(new_n296), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n291), .B1(new_n305), .B2(new_n279), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n188), .B1(new_n290), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n216), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n286), .A2(new_n287), .A3(new_n248), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n309), .A2(KEYINPUT6), .B1(new_n288), .B2(new_n283), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n281), .A2(new_n280), .A3(new_n284), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n303), .A2(new_n304), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n313), .A2(new_n295), .A3(new_n293), .ZN(new_n314));
  AOI21_X1  g128(.A(G902), .B1(new_n314), .B2(new_n309), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n315), .A3(new_n187), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n307), .A2(new_n316), .A3(KEYINPUT87), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n290), .A2(new_n306), .A3(new_n188), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT87), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(G214), .B1(G237), .B2(G902), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G131), .ZN(new_n325));
  INV_X1    g139(.A(G137), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G134), .ZN(new_n327));
  INV_X1    g141(.A(G134), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G137), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n325), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n208), .A2(G128), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT67), .B1(new_n193), .B2(KEYINPUT1), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n196), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n204), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n335));
  NOR2_X1   g149(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n327), .B2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n326), .A2(KEYINPUT65), .A3(KEYINPUT11), .A4(G134), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n337), .A2(new_n325), .A3(new_n329), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT66), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n338), .A2(new_n329), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT66), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n341), .A2(new_n342), .A3(new_n325), .A4(new_n337), .ZN(new_n343));
  AOI221_X4 g157(.A(new_n330), .B1(new_n333), .B2(new_n334), .C1(new_n340), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n343), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n337), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G131), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n201), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n263), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n333), .A2(new_n334), .ZN(new_n350));
  INV_X1    g164(.A(new_n330), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n263), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n340), .A2(new_n343), .B1(G131), .B2(new_n346), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n352), .B(new_n353), .C1(new_n354), .C2(new_n201), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT28), .ZN(new_n357));
  NOR2_X1   g171(.A1(G237), .A2(G953), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G210), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(KEYINPUT27), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT26), .B(G101), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT28), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n357), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(G902), .B1(new_n365), .B2(KEYINPUT29), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n365), .A2(KEYINPUT29), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n344), .B2(new_n348), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n352), .B(KEYINPUT30), .C1(new_n354), .C2(new_n201), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n263), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT69), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT69), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n369), .A2(new_n373), .A3(new_n370), .A4(new_n263), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n362), .B1(new_n375), .B2(new_n355), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n366), .B1(new_n367), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G472), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT32), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n355), .A2(new_n362), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT31), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n362), .B1(new_n357), .B2(new_n364), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n380), .B1(new_n372), .B2(new_n374), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT31), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(G472), .A2(G902), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n379), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n389), .ZN(new_n391));
  AOI211_X1 g205(.A(KEYINPUT32), .B(new_n391), .C1(new_n383), .C2(new_n387), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n378), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT16), .ZN(new_n394));
  INV_X1    g208(.A(G140), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n211), .B2(KEYINPUT71), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT71), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(G125), .A3(G140), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n394), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT72), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(new_n395), .A3(G125), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT72), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G146), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  OR2_X1    g219(.A1(new_n399), .A2(new_n403), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n399), .A2(new_n400), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n192), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(G119), .B(G128), .Z(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT24), .B(G110), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT23), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n220), .B2(G128), .ZN(new_n414));
  INV_X1    g228(.A(G128), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT23), .A3(G119), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n414), .B(new_n416), .C1(G119), .C2(new_n415), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n412), .B1(G110), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n409), .A2(new_n418), .ZN(new_n419));
  OR3_X1    g233(.A1(new_n417), .A2(KEYINPUT73), .A3(G110), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT73), .B1(new_n417), .B2(G110), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n410), .A2(new_n411), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G125), .B(G140), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n192), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n405), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT22), .B(G137), .ZN(new_n428));
  INV_X1    g242(.A(G221), .ZN(new_n429));
  INV_X1    g243(.A(G234), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n429), .A2(new_n430), .A3(G953), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n428), .B(new_n431), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n419), .A2(new_n426), .A3(new_n432), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n291), .A3(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n434), .A2(new_n291), .A3(new_n435), .A4(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G217), .B1(new_n430), .B2(G902), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT70), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(G902), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT75), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n434), .A2(new_n435), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT76), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n447), .A2(KEYINPUT76), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n444), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(G475), .A2(G902), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n396), .A2(new_n398), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n425), .B(KEYINPUT89), .C1(new_n192), .C2(new_n452), .ZN(new_n453));
  OR3_X1    g267(.A1(new_n452), .A2(KEYINPUT89), .A3(new_n192), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(new_n194), .ZN(new_n456));
  NOR2_X1   g270(.A1(KEYINPUT88), .A2(G143), .ZN(new_n457));
  OAI211_X1 g271(.A(G214), .B(new_n358), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n358), .A2(G214), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n455), .B2(new_n194), .ZN(new_n460));
  AND2_X1   g274(.A1(KEYINPUT18), .A2(G131), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n461), .B1(new_n458), .B2(new_n460), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n453), .B(new_n454), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n458), .A2(new_n460), .A3(new_n325), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n325), .B1(new_n458), .B2(new_n460), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT19), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n424), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n467), .B2(new_n452), .ZN(new_n469));
  OAI22_X1  g283(.A1(new_n465), .A2(new_n466), .B1(G146), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n192), .B1(new_n406), .B2(new_n407), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT90), .ZN(new_n473));
  XNOR2_X1  g287(.A(G113), .B(G122), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(new_n241), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n458), .A2(new_n460), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G131), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n458), .A2(new_n460), .A3(new_n325), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n466), .A2(KEYINPUT17), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n482), .A2(new_n408), .A3(new_n405), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n475), .A3(new_n464), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n477), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n473), .B1(new_n472), .B2(new_n476), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n451), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT20), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT20), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n490), .B(new_n451), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n484), .A2(new_n464), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n476), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n485), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n291), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n489), .A2(new_n491), .B1(G475), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G953), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G952), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(G234), .B2(G237), .ZN(new_n500));
  AOI211_X1 g314(.A(new_n291), .B(new_n498), .C1(G234), .C2(G237), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT21), .B(G898), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n218), .B2(G122), .ZN(new_n505));
  INV_X1    g319(.A(G122), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT91), .A3(G116), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n218), .A2(G122), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n253), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n237), .A3(new_n509), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT92), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n511), .A2(KEYINPUT92), .A3(new_n512), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT93), .B1(new_n415), .B2(G143), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT93), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n194), .A3(G128), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n517), .A2(new_n519), .B1(new_n415), .B2(G143), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT13), .B1(new_n415), .B2(G143), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(new_n328), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n520), .B(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n515), .A2(new_n516), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n520), .B(new_n328), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n509), .B(KEYINPUT14), .ZN(new_n526));
  INV_X1    g340(.A(new_n508), .ZN(new_n527));
  OAI21_X1  g341(.A(G107), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n512), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT9), .B(G234), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(G217), .A3(new_n498), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n524), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n533), .B1(new_n524), .B2(new_n529), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n291), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(G478), .ZN(new_n539));
  INV_X1    g353(.A(G478), .ZN(new_n540));
  OAI221_X1 g354(.A(new_n291), .B1(KEYINPUT15), .B2(new_n540), .C1(new_n535), .C2(new_n536), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n497), .A2(new_n503), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n429), .B1(new_n531), .B2(new_n291), .ZN(new_n544));
  INV_X1    g358(.A(G469), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(new_n291), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT77), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n233), .ZN(new_n548));
  NAND2_X1  g362(.A1(KEYINPUT77), .A2(G107), .ZN(new_n549));
  AOI21_X1  g363(.A(G104), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n244), .ZN(new_n551));
  OAI21_X1  g365(.A(G101), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n265), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT10), .B1(new_n210), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT80), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n555), .B(KEYINPUT1), .C1(new_n194), .C2(G146), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G128), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n193), .B2(KEYINPUT1), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n196), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n334), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT10), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n246), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n276), .A2(KEYINPUT4), .A3(new_n265), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n564), .B(new_n565), .C1(new_n260), .C2(new_n259), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n563), .A2(new_n566), .A3(new_n354), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n354), .B1(new_n563), .B2(new_n566), .ZN(new_n568));
  XNOR2_X1  g382(.A(G110), .B(G140), .ZN(new_n569));
  INV_X1    g383(.A(G227), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(G953), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n569), .B(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n567), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n563), .A2(new_n566), .A3(new_n354), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT82), .B1(new_n246), .B2(new_n350), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n246), .A2(new_n560), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT82), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n210), .A2(new_n553), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT81), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT12), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n354), .A2(new_n580), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n579), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n583), .B1(new_n579), .B2(new_n584), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n574), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n573), .B1(new_n587), .B2(new_n572), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n546), .B1(new_n588), .B2(G469), .ZN(new_n589));
  INV_X1    g403(.A(new_n572), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n590), .B(new_n574), .C1(new_n585), .C2(new_n586), .ZN(new_n591));
  OAI211_X1 g405(.A(KEYINPUT83), .B(new_n572), .C1(new_n567), .C2(new_n568), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n563), .A2(new_n566), .ZN(new_n594));
  INV_X1    g408(.A(new_n354), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n574), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT83), .B1(new_n597), .B2(new_n572), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n545), .B(new_n291), .C1(new_n593), .C2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n544), .B1(new_n589), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n543), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n324), .A2(new_n393), .A3(new_n450), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT94), .B(G101), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G3));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n187), .B1(new_n312), .B2(new_n315), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n322), .B1(new_n318), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT33), .B1(new_n535), .B2(new_n536), .ZN(new_n608));
  INV_X1    g422(.A(new_n536), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n534), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n540), .A2(G902), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT95), .B(G478), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n612), .A2(new_n613), .B1(new_n537), .B2(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n496), .A2(new_n616), .A3(new_n503), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n605), .B1(new_n607), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n323), .B1(new_n307), .B2(new_n316), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(KEYINPUT96), .A3(new_n617), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n375), .A2(new_n386), .A3(new_n381), .ZN(new_n623));
  INV_X1    g437(.A(new_n384), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n385), .A2(new_n386), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n389), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(G902), .B1(new_n383), .B2(new_n387), .ZN(new_n628));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n627), .B(new_n450), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n589), .A2(new_n599), .ZN(new_n631));
  INV_X1    g445(.A(new_n544), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n622), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NAND2_X1  g451(.A1(new_n496), .A2(new_n542), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n503), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n620), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n433), .A2(KEYINPUT36), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n427), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n427), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n446), .A3(new_n647), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n444), .A2(KEYINPUT97), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT97), .B1(new_n444), .B2(new_n648), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n644), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n444), .A2(new_n648), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n444), .A2(KEYINPUT97), .A3(new_n648), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT98), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n391), .B1(new_n383), .B2(new_n387), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n388), .A2(new_n291), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n658), .B1(new_n659), .B2(G472), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n324), .A2(new_n601), .A3(new_n657), .A4(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  XOR2_X1   g477(.A(KEYINPUT99), .B(G900), .Z(new_n664));
  AND2_X1   g478(.A1(new_n501), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n500), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n496), .A2(new_n542), .A3(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n607), .A2(new_n633), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n393), .A3(new_n657), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XNOR2_X1  g488(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n670), .B(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n633), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n321), .B(KEYINPUT38), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n649), .A2(new_n650), .ZN(new_n682));
  INV_X1    g496(.A(new_n542), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n496), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(new_n322), .A3(new_n684), .ZN(new_n685));
  NOR4_X1   g499(.A1(new_n679), .A2(new_n680), .A3(new_n681), .A4(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n362), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n375), .B2(new_n355), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n291), .B1(new_n356), .B2(new_n362), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g506(.A(KEYINPUT101), .B(G472), .C1(new_n688), .C2(new_n689), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n390), .B2(new_n392), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT102), .Z(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n686), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n686), .A2(new_n697), .A3(KEYINPUT104), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n194), .ZN(G45));
  NAND2_X1  g517(.A1(new_n307), .A2(new_n316), .ZN(new_n704));
  INV_X1    g518(.A(new_n670), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n496), .A2(new_n616), .A3(new_n705), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n322), .A2(new_n704), .A3(new_n600), .A4(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n393), .A2(new_n657), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  INV_X1    g523(.A(new_n450), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n627), .A2(KEYINPUT32), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n658), .A2(new_n379), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n710), .B1(new_n713), .B2(new_n378), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n291), .B1(new_n593), .B2(new_n598), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G469), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n632), .A3(new_n599), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n714), .A2(new_n622), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND4_X1  g535(.A1(new_n393), .A2(new_n450), .A3(new_n640), .A4(new_n718), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NOR2_X1   g539(.A1(new_n607), .A2(new_n717), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n393), .A2(new_n657), .A3(new_n543), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  INV_X1    g542(.A(new_n630), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n684), .B(new_n322), .C1(new_n318), .C2(new_n606), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n717), .A2(new_n503), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  INV_X1    g548(.A(new_n682), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n726), .A2(new_n660), .A3(new_n735), .A4(new_n706), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n323), .B1(new_n317), .B2(new_n320), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n393), .A2(new_n450), .A3(new_n600), .A4(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n706), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n739), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n633), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n714), .A3(KEYINPUT42), .A4(new_n706), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  NOR2_X1   g561(.A1(new_n740), .A2(new_n671), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT106), .B(G134), .Z(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G36));
  NAND2_X1  g564(.A1(new_n588), .A2(KEYINPUT45), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(KEYINPUT107), .Z(new_n752));
  OAI21_X1  g566(.A(G469), .B1(new_n588), .B2(KEYINPUT45), .ZN(new_n753));
  OAI22_X1  g567(.A1(new_n752), .A2(new_n753), .B1(new_n545), .B2(new_n291), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n599), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n754), .A2(new_n755), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n632), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n739), .B(KEYINPUT111), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n759), .A2(new_n676), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n496), .B(KEYINPUT108), .ZN(new_n762));
  INV_X1    g576(.A(new_n616), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(KEYINPUT43), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT43), .B1(new_n763), .B2(new_n496), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n735), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT110), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n769), .A2(new_n772), .A3(KEYINPUT44), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n761), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  NOR4_X1   g592(.A1(new_n743), .A2(new_n393), .A3(new_n450), .A4(new_n741), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n759), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n759), .A2(new_n780), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  NAND2_X1  g598(.A1(new_n716), .A2(new_n599), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT49), .Z(new_n786));
  NOR3_X1   g600(.A1(new_n616), .A2(new_n323), .A3(new_n544), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n450), .A2(new_n786), .A3(new_n762), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n696), .A2(new_n680), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n651), .A2(new_n656), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n713), .B2(new_n378), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n770), .A2(new_n682), .A3(new_n741), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n791), .A2(new_n672), .B1(new_n792), .B2(new_n726), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n652), .A2(new_n705), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n600), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n730), .A2(new_n795), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n791), .A2(new_n707), .B1(new_n695), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n695), .A2(new_n796), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n673), .A2(new_n708), .A3(new_n736), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT114), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT52), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n799), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n719), .A2(new_n602), .A3(new_n733), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n634), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n317), .A2(new_n320), .A3(new_n322), .A4(new_n617), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n810), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n634), .A2(new_n324), .A3(new_n639), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n661), .A3(new_n727), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n809), .A2(new_n724), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n748), .B1(new_n742), .B2(new_n745), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n497), .A2(new_n542), .A3(new_n705), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n791), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n744), .B1(new_n823), .B2(new_n792), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n820), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n807), .A2(new_n826), .A3(KEYINPUT53), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n793), .A2(new_n797), .A3(KEYINPUT113), .A4(KEYINPUT52), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n829), .B1(new_n801), .B2(new_n805), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n806), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n827), .B1(KEYINPUT53), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT54), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n826), .A2(KEYINPUT53), .A3(new_n831), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT53), .B1(new_n807), .B2(new_n826), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n743), .A2(new_n717), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n450), .A2(new_n696), .A3(new_n500), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n496), .A3(new_n616), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n668), .B1(new_n766), .B2(new_n768), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n844), .A2(new_n841), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n660), .A3(new_n735), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n844), .A2(new_n729), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n680), .A2(new_n323), .A3(new_n718), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OR3_X1    g665(.A1(new_n849), .A2(new_n848), .A3(new_n850), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n849), .A2(new_n760), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n759), .B(new_n780), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n785), .A2(new_n632), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT115), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n854), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT51), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n853), .A2(KEYINPUT51), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n842), .A2(new_n497), .A3(new_n763), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n845), .A2(new_n714), .ZN(new_n863));
  XOR2_X1   g677(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n849), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n499), .B1(new_n866), .B2(new_n726), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n845), .A2(KEYINPUT116), .A3(KEYINPUT48), .A4(new_n714), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n862), .A2(new_n865), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n861), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n840), .A2(new_n859), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(G952), .A2(G953), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n789), .B1(new_n871), .B2(new_n872), .ZN(G75));
  NOR2_X1   g687(.A1(new_n498), .A2(G952), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(G210), .A2(G902), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n799), .A2(new_n802), .A3(new_n805), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n805), .B1(new_n799), .B2(new_n802), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n808), .A2(new_n818), .A3(new_n815), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n821), .A3(new_n724), .A4(new_n824), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n877), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n826), .A2(KEYINPUT53), .A3(new_n831), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n876), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n285), .A2(new_n289), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT117), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n216), .B(KEYINPUT55), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n885), .A2(KEYINPUT120), .A3(KEYINPUT56), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n891));
  INV_X1    g705(.A(new_n876), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n835), .B2(new_n836), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n889), .A2(KEYINPUT56), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n875), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n897), .B1(new_n885), .B2(new_n898), .ZN(new_n899));
  AOI211_X1 g713(.A(KEYINPUT118), .B(new_n876), .C1(new_n883), .C2(new_n884), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n889), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT119), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n903), .B(new_n889), .C1(new_n899), .C2(new_n900), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n896), .B1(new_n902), .B2(new_n904), .ZN(G51));
  NAND2_X1  g719(.A1(new_n883), .A2(new_n884), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n838), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n546), .B(KEYINPUT57), .Z(new_n908));
  OAI22_X1  g722(.A1(new_n907), .A2(new_n908), .B1(new_n598), .B2(new_n593), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n837), .A2(new_n291), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n752), .A2(new_n753), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n874), .B1(new_n909), .B2(new_n912), .ZN(G54));
  NAND3_X1  g727(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n486), .A2(new_n487), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .A4(new_n915), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n917), .A2(new_n875), .A3(new_n918), .ZN(G60));
  XOR2_X1   g733(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n920));
  NOR2_X1   g734(.A1(new_n540), .A2(new_n291), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n612), .B1(new_n840), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n612), .A2(new_n922), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n875), .B1(new_n907), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n925), .ZN(G63));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n646), .A2(new_n647), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT60), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n929), .B(new_n932), .C1(new_n835), .C2(new_n836), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n875), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n931), .B1(new_n883), .B2(new_n884), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n434), .A2(new_n435), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n927), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT122), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n927), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n934), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT123), .B1(new_n935), .B2(new_n937), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n946), .B(new_n927), .C1(new_n934), .C2(new_n938), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n940), .A2(new_n945), .A3(new_n947), .ZN(G66));
  OAI21_X1  g762(.A(G953), .B1(new_n502), .B2(new_n214), .ZN(new_n949));
  INV_X1    g763(.A(new_n820), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(new_n950), .B2(G953), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n887), .B1(G898), .B2(new_n498), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT124), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n951), .B(new_n953), .ZN(G69));
  NAND2_X1  g768(.A1(new_n369), .A2(new_n370), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(new_n469), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n700), .A2(new_n701), .A3(new_n708), .A4(new_n793), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n638), .B1(new_n496), .B2(new_n616), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n714), .A2(new_n677), .A3(new_n739), .A4(new_n959), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT125), .Z(new_n961));
  AND3_X1   g775(.A1(new_n783), .A2(new_n777), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n958), .A2(new_n498), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n956), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n570), .A2(G900), .A3(G953), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n783), .A2(new_n777), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n759), .A2(new_n676), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n714), .A2(new_n731), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AND4_X1   g785(.A1(new_n708), .A2(new_n971), .A3(new_n821), .A4(new_n793), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT126), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n968), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n967), .B1(new_n977), .B2(G953), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n966), .B1(new_n978), .B2(new_n956), .ZN(G72));
  NAND3_X1  g793(.A1(new_n375), .A2(new_n355), .A3(new_n687), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n974), .A2(new_n950), .A3(new_n976), .ZN(new_n981));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT63), .Z(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT127), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n980), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n688), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n958), .A2(new_n950), .A3(new_n962), .A4(new_n963), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n984), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n376), .A2(new_n385), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n833), .A2(new_n983), .A3(new_n989), .ZN(new_n990));
  NOR4_X1   g804(.A1(new_n985), .A2(new_n988), .A3(new_n990), .A4(new_n874), .ZN(G57));
endmodule


