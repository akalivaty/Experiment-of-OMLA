

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582;

  XOR2_X1 U324 ( .A(KEYINPUT100), .B(n467), .Z(n515) );
  XNOR2_X1 U325 ( .A(n401), .B(KEYINPUT48), .ZN(n402) );
  XNOR2_X1 U326 ( .A(n403), .B(n402), .ZN(n527) );
  NOR2_X1 U327 ( .A1(n437), .A2(n515), .ZN(n565) );
  XOR2_X1 U328 ( .A(KEYINPUT36), .B(n561), .Z(n579) );
  XOR2_X1 U329 ( .A(n354), .B(n353), .Z(n561) );
  XNOR2_X1 U330 ( .A(n458), .B(G176GAT), .ZN(n459) );
  XNOR2_X1 U331 ( .A(n460), .B(n459), .ZN(G1349GAT) );
  XOR2_X1 U332 ( .A(G99GAT), .B(KEYINPUT72), .Z(n293) );
  XNOR2_X1 U333 ( .A(G85GAT), .B(G106GAT), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n341) );
  XOR2_X1 U335 ( .A(KEYINPUT13), .B(G78GAT), .Z(n295) );
  XNOR2_X1 U336 ( .A(G57GAT), .B(G71GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n375) );
  XNOR2_X1 U338 ( .A(n341), .B(n375), .ZN(n310) );
  XOR2_X1 U339 ( .A(G148GAT), .B(KEYINPUT71), .Z(n315) );
  XOR2_X1 U340 ( .A(KEYINPUT73), .B(n315), .Z(n299) );
  XOR2_X1 U341 ( .A(G204GAT), .B(G176GAT), .Z(n297) );
  XNOR2_X1 U342 ( .A(G92GAT), .B(G64GAT), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n407) );
  XNOR2_X1 U344 ( .A(G120GAT), .B(n407), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U346 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n301) );
  NAND2_X1 U347 ( .A1(G230GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U349 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U350 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n305) );
  XNOR2_X1 U351 ( .A(KEYINPUT75), .B(KEYINPUT33), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n306), .B(KEYINPUT77), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n310), .B(n309), .ZN(n572) );
  NAND2_X1 U356 ( .A1(n572), .A2(KEYINPUT41), .ZN(n314) );
  INV_X1 U357 ( .A(n572), .ZN(n312) );
  INV_X1 U358 ( .A(KEYINPUT41), .ZN(n311) );
  NAND2_X1 U359 ( .A1(n312), .A2(n311), .ZN(n313) );
  NAND2_X1 U360 ( .A1(n314), .A2(n313), .ZN(n548) );
  XNOR2_X1 U361 ( .A(KEYINPUT112), .B(n548), .ZN(n533) );
  XOR2_X1 U362 ( .A(G155GAT), .B(G22GAT), .Z(n388) );
  XOR2_X1 U363 ( .A(n315), .B(n388), .Z(n317) );
  XNOR2_X1 U364 ( .A(G106GAT), .B(G50GAT), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n326) );
  XOR2_X1 U366 ( .A(G197GAT), .B(KEYINPUT95), .Z(n319) );
  XNOR2_X1 U367 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n412) );
  XOR2_X1 U369 ( .A(G204GAT), .B(n412), .Z(n324) );
  XOR2_X1 U370 ( .A(KEYINPUT2), .B(G162GAT), .Z(n321) );
  XNOR2_X1 U371 ( .A(KEYINPUT96), .B(G141GAT), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U373 ( .A(KEYINPUT3), .B(n322), .Z(n430) );
  XNOR2_X1 U374 ( .A(n430), .B(G211GAT), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U376 ( .A(n326), .B(n325), .Z(n328) );
  NAND2_X1 U377 ( .A1(G228GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n336) );
  XOR2_X1 U379 ( .A(KEYINPUT22), .B(KEYINPUT94), .Z(n330) );
  XNOR2_X1 U380 ( .A(G78GAT), .B(KEYINPUT97), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U382 ( .A(KEYINPUT23), .B(KEYINPUT98), .Z(n332) );
  XNOR2_X1 U383 ( .A(KEYINPUT99), .B(KEYINPUT24), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U385 ( .A(n334), .B(n333), .Z(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n471) );
  XOR2_X1 U387 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n338) );
  XNOR2_X1 U388 ( .A(KEYINPUT80), .B(KEYINPUT10), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n354) );
  XOR2_X1 U390 ( .A(G50GAT), .B(G43GAT), .Z(n340) );
  XNOR2_X1 U391 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n357) );
  XNOR2_X1 U393 ( .A(n341), .B(n357), .ZN(n346) );
  XOR2_X1 U394 ( .A(KEYINPUT67), .B(KEYINPUT79), .Z(n343) );
  NAND2_X1 U395 ( .A1(G232GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U397 ( .A(n344), .B(KEYINPUT78), .Z(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U399 ( .A(KEYINPUT11), .B(G218GAT), .Z(n348) );
  XOR2_X1 U400 ( .A(G29GAT), .B(G134GAT), .Z(n429) );
  XOR2_X1 U401 ( .A(G190GAT), .B(G36GAT), .Z(n404) );
  XNOR2_X1 U402 ( .A(n429), .B(n404), .ZN(n347) );
  XOR2_X1 U403 ( .A(n348), .B(n347), .Z(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n352) );
  XNOR2_X1 U405 ( .A(G162GAT), .B(G92GAT), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n353) );
  INV_X1 U407 ( .A(n561), .ZN(n554) );
  XOR2_X1 U408 ( .A(G169GAT), .B(G22GAT), .Z(n356) );
  XNOR2_X1 U409 ( .A(G113GAT), .B(G141GAT), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n370) );
  XOR2_X1 U411 ( .A(G15GAT), .B(KEYINPUT70), .Z(n387) );
  XOR2_X1 U412 ( .A(n387), .B(G36GAT), .Z(n359) );
  XNOR2_X1 U413 ( .A(G29GAT), .B(n357), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U415 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n361) );
  NAND2_X1 U416 ( .A1(G229GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U418 ( .A(n363), .B(n362), .Z(n368) );
  XOR2_X1 U419 ( .A(KEYINPUT69), .B(G197GAT), .Z(n365) );
  XNOR2_X1 U420 ( .A(G1GAT), .B(G8GAT), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n366), .B(KEYINPUT29), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U424 ( .A(n370), .B(n369), .Z(n568) );
  INV_X1 U425 ( .A(n568), .ZN(n556) );
  NOR2_X1 U426 ( .A1(n556), .A2(n548), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n371), .B(KEYINPUT46), .ZN(n372) );
  NOR2_X1 U428 ( .A1(n554), .A2(n372), .ZN(n393) );
  XOR2_X1 U429 ( .A(KEYINPUT84), .B(KEYINPUT14), .Z(n374) );
  XNOR2_X1 U430 ( .A(KEYINPUT12), .B(KEYINPUT83), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n379) );
  XOR2_X1 U432 ( .A(n375), .B(KEYINPUT86), .Z(n377) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n392) );
  XOR2_X1 U436 ( .A(KEYINPUT85), .B(KEYINPUT82), .Z(n381) );
  XNOR2_X1 U437 ( .A(KEYINPUT87), .B(KEYINPUT81), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U439 ( .A(n382), .B(KEYINPUT15), .Z(n384) );
  XOR2_X1 U440 ( .A(G127GAT), .B(G1GAT), .Z(n422) );
  XNOR2_X1 U441 ( .A(n422), .B(G64GAT), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n386) );
  XNOR2_X1 U443 ( .A(G183GAT), .B(G211GAT), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n385), .B(G8GAT), .ZN(n416) );
  XOR2_X1 U445 ( .A(n386), .B(n416), .Z(n390) );
  XNOR2_X1 U446 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n575) );
  XNOR2_X1 U449 ( .A(n575), .B(KEYINPUT117), .ZN(n558) );
  NAND2_X1 U450 ( .A1(n393), .A2(n558), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n394), .B(KEYINPUT47), .ZN(n400) );
  XOR2_X1 U452 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n396) );
  NAND2_X1 U453 ( .A1(n575), .A2(n579), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  NAND2_X1 U455 ( .A1(n397), .A2(n556), .ZN(n398) );
  NOR2_X1 U456 ( .A1(n398), .A2(n572), .ZN(n399) );
  NOR2_X1 U457 ( .A1(n400), .A2(n399), .ZN(n403) );
  INV_X1 U458 ( .A(KEYINPUT64), .ZN(n401) );
  XOR2_X1 U459 ( .A(KEYINPUT101), .B(n404), .Z(n406) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U462 ( .A(n408), .B(n407), .Z(n414) );
  XOR2_X1 U463 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n410) );
  XNOR2_X1 U464 ( .A(KEYINPUT17), .B(G169GAT), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U466 ( .A(KEYINPUT19), .B(n411), .Z(n452) );
  XNOR2_X1 U467 ( .A(n452), .B(n412), .ZN(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U469 ( .A(n416), .B(n415), .ZN(n518) );
  NAND2_X1 U470 ( .A1(n527), .A2(n518), .ZN(n418) );
  XOR2_X1 U471 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n417) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n437) );
  XOR2_X1 U473 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n420) );
  XNOR2_X1 U474 ( .A(G155GAT), .B(G57GAT), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U476 ( .A(n421), .B(G148GAT), .Z(n424) );
  XNOR2_X1 U477 ( .A(n422), .B(G85GAT), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U479 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n426) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U482 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U485 ( .A(KEYINPUT0), .B(KEYINPUT89), .Z(n434) );
  XNOR2_X1 U486 ( .A(G120GAT), .B(G113GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U488 ( .A(KEYINPUT88), .B(n435), .Z(n456) );
  XNOR2_X1 U489 ( .A(n436), .B(n456), .ZN(n467) );
  NAND2_X1 U490 ( .A1(n471), .A2(n565), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n438), .B(KEYINPUT55), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n439), .B(KEYINPUT122), .ZN(n457) );
  XOR2_X1 U493 ( .A(G176GAT), .B(KEYINPUT90), .Z(n441) );
  XNOR2_X1 U494 ( .A(G127GAT), .B(G71GAT), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U496 ( .A(KEYINPUT20), .B(KEYINPUT92), .Z(n443) );
  XNOR2_X1 U497 ( .A(G183GAT), .B(KEYINPUT93), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U499 ( .A(n445), .B(n444), .Z(n454) );
  XOR2_X1 U500 ( .A(G190GAT), .B(G43GAT), .Z(n447) );
  XNOR2_X1 U501 ( .A(G134GAT), .B(G99GAT), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(G15GAT), .B(n448), .Z(n450) );
  NAND2_X1 U504 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n456), .B(n455), .ZN(n530) );
  INV_X1 U509 ( .A(n530), .ZN(n520) );
  NAND2_X1 U510 ( .A1(n457), .A2(n520), .ZN(n560) );
  NOR2_X1 U511 ( .A1(n533), .A2(n560), .ZN(n460) );
  XNOR2_X1 U512 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n458) );
  NOR2_X1 U513 ( .A1(n556), .A2(n572), .ZN(n491) );
  NAND2_X1 U514 ( .A1(n518), .A2(n520), .ZN(n461) );
  NAND2_X1 U515 ( .A1(n461), .A2(n471), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n462), .B(KEYINPUT25), .ZN(n463) );
  XNOR2_X1 U517 ( .A(n463), .B(KEYINPUT103), .ZN(n466) );
  XNOR2_X1 U518 ( .A(KEYINPUT27), .B(n518), .ZN(n469) );
  NOR2_X1 U519 ( .A1(n471), .A2(n520), .ZN(n464) );
  XNOR2_X1 U520 ( .A(n464), .B(KEYINPUT26), .ZN(n566) );
  NAND2_X1 U521 ( .A1(n469), .A2(n566), .ZN(n465) );
  NAND2_X1 U522 ( .A1(n466), .A2(n465), .ZN(n468) );
  NAND2_X1 U523 ( .A1(n468), .A2(n467), .ZN(n473) );
  NAND2_X1 U524 ( .A1(n515), .A2(n469), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT102), .ZN(n545) );
  XOR2_X1 U526 ( .A(n471), .B(KEYINPUT28), .Z(n524) );
  NOR2_X1 U527 ( .A1(n545), .A2(n524), .ZN(n528) );
  NAND2_X1 U528 ( .A1(n528), .A2(n530), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n473), .A2(n472), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT104), .B(n474), .Z(n487) );
  NAND2_X1 U531 ( .A1(n561), .A2(n575), .ZN(n475) );
  XNOR2_X1 U532 ( .A(KEYINPUT16), .B(n475), .ZN(n476) );
  NOR2_X1 U533 ( .A1(n487), .A2(n476), .ZN(n504) );
  AND2_X1 U534 ( .A1(n491), .A2(n504), .ZN(n483) );
  NAND2_X1 U535 ( .A1(n515), .A2(n483), .ZN(n477) );
  XNOR2_X1 U536 ( .A(KEYINPUT34), .B(n477), .ZN(n478) );
  XNOR2_X1 U537 ( .A(G1GAT), .B(n478), .ZN(G1324GAT) );
  NAND2_X1 U538 ( .A1(n518), .A2(n483), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n479), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT35), .B(KEYINPUT105), .Z(n481) );
  NAND2_X1 U541 ( .A1(n483), .A2(n520), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U543 ( .A(G15GAT), .B(n482), .Z(G1326GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n485) );
  NAND2_X1 U545 ( .A1(n483), .A2(n524), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(n486), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT109), .B(KEYINPUT39), .Z(n494) );
  NOR2_X1 U549 ( .A1(n575), .A2(n487), .ZN(n488) );
  XNOR2_X1 U550 ( .A(KEYINPUT108), .B(n488), .ZN(n489) );
  NAND2_X1 U551 ( .A1(n489), .A2(n579), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n490), .B(KEYINPUT37), .ZN(n514) );
  NAND2_X1 U553 ( .A1(n491), .A2(n514), .ZN(n492) );
  XOR2_X1 U554 ( .A(KEYINPUT38), .B(n492), .Z(n500) );
  NAND2_X1 U555 ( .A1(n500), .A2(n515), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U557 ( .A(G29GAT), .B(n495), .Z(G1328GAT) );
  NAND2_X1 U558 ( .A1(n500), .A2(n518), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(KEYINPUT110), .ZN(n497) );
  XNOR2_X1 U560 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n500), .A2(n520), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n498), .B(KEYINPUT40), .ZN(n499) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n500), .A2(n524), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n503) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT113), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(n506) );
  NOR2_X1 U569 ( .A1(n568), .A2(n533), .ZN(n513) );
  AND2_X1 U570 ( .A1(n513), .A2(n504), .ZN(n510) );
  NAND2_X1 U571 ( .A1(n515), .A2(n510), .ZN(n505) );
  XOR2_X1 U572 ( .A(n506), .B(n505), .Z(G1332GAT) );
  NAND2_X1 U573 ( .A1(n518), .A2(n510), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n507), .B(KEYINPUT114), .ZN(n508) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n510), .A2(n520), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n509), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U579 ( .A1(n510), .A2(n524), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  XOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT115), .Z(n517) );
  AND2_X1 U582 ( .A1(n514), .A2(n513), .ZN(n523) );
  NAND2_X1 U583 ( .A1(n523), .A2(n515), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n518), .A2(n523), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n520), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(KEYINPUT116), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(n522), .ZN(G1338GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n541), .A2(n568), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT118), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  INV_X1 U598 ( .A(n541), .ZN(n537) );
  NOR2_X1 U599 ( .A1(n533), .A2(n537), .ZN(n535) );
  XNOR2_X1 U600 ( .A(KEYINPUT119), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n536), .Z(G1341GAT) );
  NOR2_X1 U603 ( .A1(n558), .A2(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT120), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n540), .Z(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n554), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n566), .A2(n527), .ZN(n544) );
  NOR2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n553), .A2(n568), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(G141GAT), .ZN(G1344GAT) );
  INV_X1 U614 ( .A(n553), .ZN(n547) );
  NOR2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n553), .A2(n575), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n560), .ZN(n557) );
  XOR2_X1 U624 ( .A(G169GAT), .B(n557), .Z(G1348GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n558), .ZN(n559) );
  XOR2_X1 U626 ( .A(G183GAT), .B(n559), .Z(G1350GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U628 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(n567), .B(KEYINPUT124), .Z(n580) );
  AND2_X1 U633 ( .A1(n580), .A2(n568), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n572), .A2(n580), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n577) );
  NAND2_X1 U641 ( .A1(n575), .A2(n580), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

