

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751;

  XNOR2_X1 U373 ( .A(n714), .B(n715), .ZN(n356) );
  INV_X1 U374 ( .A(n717), .ZN(n353) );
  AND2_X1 U375 ( .A1(n404), .A2(n557), .ZN(n403) );
  XNOR2_X1 U376 ( .A(n570), .B(n434), .ZN(n659) );
  OR2_X1 U377 ( .A1(n694), .A2(G902), .ZN(n437) );
  XNOR2_X1 U378 ( .A(n502), .B(n501), .ZN(n399) );
  XNOR2_X1 U379 ( .A(n446), .B(n445), .ZN(n400) );
  BUF_X1 U380 ( .A(G137), .Z(n351) );
  XNOR2_X2 U381 ( .A(n464), .B(KEYINPUT89), .ZN(n617) );
  XNOR2_X2 U382 ( .A(n651), .B(KEYINPUT83), .ZN(n587) );
  XNOR2_X2 U383 ( .A(n539), .B(n538), .ZN(n676) );
  XNOR2_X2 U384 ( .A(n536), .B(KEYINPUT105), .ZN(n548) );
  NOR2_X2 U385 ( .A1(n676), .A2(n540), .ZN(n541) );
  XNOR2_X2 U386 ( .A(n453), .B(n452), .ZN(n718) );
  XNOR2_X2 U387 ( .A(n400), .B(n447), .ZN(n453) );
  NOR2_X2 U388 ( .A1(n393), .A2(n392), .ZN(n391) );
  NAND2_X2 U389 ( .A1(n615), .A2(n751), .ZN(n612) );
  INV_X1 U390 ( .A(n352), .ZN(G54) );
  NAND2_X1 U391 ( .A1(n354), .A2(n353), .ZN(n352) );
  XNOR2_X1 U392 ( .A(n697), .B(n355), .ZN(n354) );
  INV_X1 U393 ( .A(n698), .ZN(n355) );
  NOR2_X1 U394 ( .A1(n356), .A2(n717), .ZN(G66) );
  XNOR2_X1 U395 ( .A(G143), .B(G113), .ZN(n510) );
  INV_X2 U396 ( .A(G953), .ZN(n728) );
  OR2_X2 U397 ( .A1(n431), .A2(n430), .ZN(n404) );
  AND2_X2 U398 ( .A1(n681), .A2(n617), .ZN(n416) );
  INV_X1 U399 ( .A(KEYINPUT3), .ZN(n445) );
  AND2_X1 U400 ( .A1(n401), .A2(n406), .ZN(n405) );
  XNOR2_X1 U401 ( .A(n531), .B(KEYINPUT22), .ZN(n550) );
  NAND2_X1 U402 ( .A1(n382), .A2(n385), .ZN(n583) );
  XNOR2_X1 U403 ( .A(n413), .B(n412), .ZN(n530) );
  NOR2_X1 U404 ( .A1(n585), .A2(n360), .ZN(n413) );
  NOR2_X1 U405 ( .A1(n555), .A2(KEYINPUT44), .ZN(n357) );
  INV_X1 U406 ( .A(n597), .ZN(n358) );
  NOR2_X1 U407 ( .A1(n555), .A2(KEYINPUT44), .ZN(n431) );
  XNOR2_X1 U408 ( .A(n470), .B(n471), .ZN(n585) );
  AND2_X2 U409 ( .A1(n416), .A2(n414), .ZN(n359) );
  NOR2_X1 U410 ( .A1(n586), .A2(n585), .ZN(n638) );
  INV_X1 U411 ( .A(G469), .ZN(n436) );
  NAND2_X1 U412 ( .A1(n749), .A2(n632), .ZN(n556) );
  NOR2_X1 U413 ( .A1(G953), .A2(G237), .ZN(n508) );
  XNOR2_X1 U414 ( .A(n432), .B(KEYINPUT69), .ZN(n478) );
  XNOR2_X1 U415 ( .A(G134), .B(G131), .ZN(n432) );
  NAND2_X1 U416 ( .A1(n399), .A2(n655), .ZN(n658) );
  INV_X1 U417 ( .A(KEYINPUT87), .ZN(n371) );
  XOR2_X1 U418 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n457) );
  INV_X1 U419 ( .A(KEYINPUT91), .ZN(n455) );
  INV_X1 U420 ( .A(KEYINPUT93), .ZN(n477) );
  XNOR2_X1 U421 ( .A(G110), .B(G107), .ZN(n721) );
  XOR2_X1 U422 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n521) );
  XNOR2_X1 U423 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n520) );
  XNOR2_X1 U424 ( .A(n527), .B(KEYINPUT9), .ZN(n425) );
  XNOR2_X1 U425 ( .A(G116), .B(G134), .ZN(n518) );
  XOR2_X1 U426 ( .A(G122), .B(G107), .Z(n519) );
  XNOR2_X1 U427 ( .A(n428), .B(n507), .ZN(n427) );
  XNOR2_X1 U428 ( .A(n466), .B(KEYINPUT79), .ZN(n467) );
  INV_X1 U429 ( .A(n583), .ZN(n390) );
  AND2_X1 U430 ( .A1(n637), .A2(n647), .ZN(n426) );
  NOR2_X1 U431 ( .A1(n708), .A2(G902), .ZN(n528) );
  XNOR2_X1 U432 ( .A(n435), .B(KEYINPUT65), .ZN(n434) );
  INV_X1 U433 ( .A(KEYINPUT1), .ZN(n435) );
  AND2_X1 U434 ( .A1(n638), .A2(n588), .ZN(n420) );
  NAND2_X1 U435 ( .A1(G234), .A2(G237), .ZN(n472) );
  XNOR2_X1 U436 ( .A(n422), .B(n421), .ZN(n651) );
  INV_X1 U437 ( .A(KEYINPUT103), .ZN(n421) );
  NOR2_X1 U438 ( .A1(n637), .A2(n633), .ZN(n422) );
  INV_X1 U439 ( .A(KEYINPUT48), .ZN(n439) );
  XOR2_X1 U440 ( .A(G137), .B(G140), .Z(n490) );
  XNOR2_X1 U441 ( .A(n509), .B(n506), .ZN(n428) );
  XOR2_X1 U442 ( .A(G140), .B(G131), .Z(n511) );
  XOR2_X1 U443 ( .A(G104), .B(G122), .Z(n513) );
  XOR2_X1 U444 ( .A(KEYINPUT77), .B(G104), .Z(n480) );
  XNOR2_X1 U445 ( .A(n478), .B(n433), .ZN(n734) );
  XNOR2_X1 U446 ( .A(n490), .B(KEYINPUT94), .ZN(n433) );
  NOR2_X1 U447 ( .A1(G902), .A2(G237), .ZN(n465) );
  XNOR2_X1 U448 ( .A(G902), .B(KEYINPUT15), .ZN(n464) );
  XOR2_X1 U449 ( .A(KEYINPUT21), .B(n488), .Z(n655) );
  NAND2_X1 U450 ( .A1(n389), .A2(n398), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n517), .B(n516), .ZN(n543) );
  XNOR2_X1 U452 ( .A(n449), .B(n351), .ZN(n443) );
  INV_X1 U453 ( .A(KEYINPUT45), .ZN(n560) );
  XNOR2_X1 U454 ( .A(n372), .B(n371), .ZN(n559) );
  XNOR2_X1 U455 ( .A(G119), .B(G128), .ZN(n494) );
  XNOR2_X1 U456 ( .A(n381), .B(n490), .ZN(n493) );
  XNOR2_X1 U457 ( .A(n463), .B(n462), .ZN(n688) );
  XNOR2_X1 U458 ( .A(n718), .B(n454), .ZN(n463) );
  INV_X1 U459 ( .A(KEYINPUT0), .ZN(n412) );
  NAND2_X1 U460 ( .A1(n396), .A2(n581), .ZN(n395) );
  AND2_X1 U461 ( .A1(n383), .A2(n367), .ZN(n382) );
  NOR2_X1 U462 ( .A1(n387), .A2(KEYINPUT30), .ZN(n386) );
  XNOR2_X1 U463 ( .A(n526), .B(n424), .ZN(n708) );
  XNOR2_X1 U464 ( .A(n525), .B(n425), .ZN(n424) );
  XNOR2_X1 U465 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U466 ( .A1(G952), .A2(n728), .ZN(n717) );
  XNOR2_X1 U467 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n576) );
  INV_X1 U468 ( .A(KEYINPUT40), .ZN(n369) );
  NOR2_X1 U469 ( .A1(n659), .A2(n598), .ZN(n599) );
  XNOR2_X1 U470 ( .A(n377), .B(KEYINPUT36), .ZN(n598) );
  OR2_X1 U471 ( .A1(n602), .A2(n597), .ZN(n377) );
  XNOR2_X1 U472 ( .A(KEYINPUT32), .B(n553), .ZN(n749) );
  NOR2_X1 U473 ( .A1(n550), .A2(n659), .ZN(n551) );
  AND2_X1 U474 ( .A1(n542), .A2(n423), .ZN(n633) );
  INV_X1 U475 ( .A(KEYINPUT64), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n686), .B(n373), .ZN(G75) );
  XNOR2_X1 U477 ( .A(n374), .B(KEYINPUT53), .ZN(n373) );
  INV_X1 U478 ( .A(KEYINPUT117), .ZN(n374) );
  NOR2_X1 U479 ( .A1(n564), .A2(n476), .ZN(n360) );
  NOR2_X1 U480 ( .A1(n567), .A2(n399), .ZN(n361) );
  XNOR2_X1 U481 ( .A(KEYINPUT95), .B(KEYINPUT5), .ZN(n362) );
  AND2_X1 U482 ( .A1(n596), .A2(n361), .ZN(n363) );
  AND2_X1 U483 ( .A1(n532), .A2(n659), .ZN(n364) );
  XNOR2_X1 U484 ( .A(n597), .B(n573), .ZN(n646) );
  NAND2_X1 U485 ( .A1(n655), .A2(n574), .ZN(n365) );
  OR2_X1 U486 ( .A1(n593), .A2(n418), .ZN(n366) );
  INV_X1 U487 ( .A(KEYINPUT76), .ZN(n581) );
  OR2_X1 U488 ( .A1(n647), .A2(n388), .ZN(n367) );
  BUF_X1 U489 ( .A(n681), .Z(n368) );
  BUF_X1 U490 ( .A(n359), .Z(n713) );
  NAND2_X1 U491 ( .A1(n679), .A2(n415), .ZN(n414) );
  NAND2_X1 U492 ( .A1(n391), .A2(n390), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n453), .B(n442), .ZN(n450) );
  XNOR2_X2 U494 ( .A(n370), .B(n369), .ZN(n750) );
  NAND2_X1 U495 ( .A1(n609), .A2(n637), .ZN(n370) );
  XNOR2_X1 U496 ( .A(n429), .B(n427), .ZN(n515) );
  INV_X1 U497 ( .A(n543), .ZN(n423) );
  INV_X1 U498 ( .A(n550), .ZN(n532) );
  NOR2_X2 U499 ( .A1(G902), .A2(n618), .ZN(n451) );
  XNOR2_X1 U500 ( .A(n409), .B(n408), .ZN(n407) );
  NOR2_X2 U501 ( .A1(n704), .A2(n717), .ZN(n706) );
  NAND2_X1 U502 ( .A1(n548), .A2(n547), .ZN(n372) );
  NOR2_X2 U503 ( .A1(n621), .A2(n717), .ZN(n375) );
  NOR2_X2 U504 ( .A1(n691), .A2(n717), .ZN(n376) );
  XNOR2_X2 U505 ( .A(n546), .B(KEYINPUT35), .ZN(n555) );
  INV_X2 U506 ( .A(n533), .ZN(n662) );
  XNOR2_X2 U507 ( .A(n451), .B(G472), .ZN(n533) );
  NOR2_X2 U508 ( .A1(n750), .A2(n746), .ZN(n584) );
  NAND2_X1 U509 ( .A1(n384), .A2(KEYINPUT30), .ZN(n383) );
  NAND2_X1 U510 ( .A1(n748), .A2(n600), .ZN(n601) );
  XNOR2_X1 U511 ( .A(n599), .B(KEYINPUT113), .ZN(n748) );
  XNOR2_X1 U512 ( .A(n375), .B(n623), .ZN(G57) );
  XNOR2_X1 U513 ( .A(n376), .B(n693), .ZN(G51) );
  AND2_X2 U514 ( .A1(n378), .A2(n608), .ZN(n615) );
  XNOR2_X1 U515 ( .A(n379), .B(n439), .ZN(n378) );
  NAND2_X1 U516 ( .A1(n440), .A2(n380), .ZN(n379) );
  XNOR2_X1 U517 ( .A(n584), .B(KEYINPUT46), .ZN(n380) );
  XNOR2_X1 U518 ( .A(n512), .B(n381), .ZN(n429) );
  XNOR2_X1 U519 ( .A(n381), .B(n736), .ZN(n741) );
  XNOR2_X2 U520 ( .A(n489), .B(KEYINPUT10), .ZN(n381) );
  INV_X1 U521 ( .A(n438), .ZN(n384) );
  NAND2_X1 U522 ( .A1(n438), .A2(n386), .ZN(n385) );
  INV_X1 U523 ( .A(n647), .ZN(n387) );
  INV_X1 U524 ( .A(KEYINPUT30), .ZN(n388) );
  OR2_X2 U525 ( .A1(n579), .A2(n395), .ZN(n394) );
  INV_X1 U526 ( .A(n392), .ZN(n397) );
  NAND2_X1 U527 ( .A1(n579), .A2(KEYINPUT76), .ZN(n389) );
  NAND2_X1 U528 ( .A1(n397), .A2(n394), .ZN(n582) );
  NAND2_X1 U529 ( .A1(n394), .A2(n646), .ZN(n393) );
  INV_X1 U530 ( .A(n580), .ZN(n396) );
  NAND2_X1 U531 ( .A1(n580), .A2(KEYINPUT76), .ZN(n398) );
  INV_X1 U532 ( .A(n399), .ZN(n554) );
  XNOR2_X1 U533 ( .A(n554), .B(KEYINPUT104), .ZN(n549) );
  NAND2_X1 U534 ( .A1(n402), .A2(n357), .ZN(n401) );
  NOR2_X1 U535 ( .A1(n556), .A2(KEYINPUT73), .ZN(n402) );
  NAND2_X1 U536 ( .A1(n556), .A2(KEYINPUT73), .ZN(n406) );
  NAND2_X1 U537 ( .A1(n405), .A2(n403), .ZN(n558) );
  NAND2_X1 U538 ( .A1(n407), .A2(n554), .ZN(n632) );
  NAND2_X1 U539 ( .A1(n532), .A2(n410), .ZN(n409) );
  NOR2_X1 U540 ( .A1(n438), .A2(n411), .ZN(n410) );
  INV_X1 U541 ( .A(n659), .ZN(n411) );
  XNOR2_X1 U542 ( .A(n448), .B(n443), .ZN(n442) );
  NOR2_X1 U543 ( .A1(n601), .A2(n366), .ZN(n440) );
  NOR2_X2 U544 ( .A1(n688), .A2(n617), .ZN(n468) );
  XNOR2_X2 U545 ( .A(G143), .B(G128), .ZN(n527) );
  XNOR2_X1 U546 ( .A(n493), .B(n444), .ZN(n498) );
  NOR2_X2 U547 ( .A1(n570), .A2(n658), .ZN(n578) );
  INV_X1 U548 ( .A(KEYINPUT2), .ZN(n415) );
  XNOR2_X2 U549 ( .A(n612), .B(n611), .ZN(n740) );
  NAND2_X1 U550 ( .A1(n729), .A2(n417), .ZN(n681) );
  XNOR2_X1 U551 ( .A(n616), .B(KEYINPUT85), .ZN(n417) );
  XNOR2_X2 U552 ( .A(n561), .B(n560), .ZN(n729) );
  NAND2_X1 U553 ( .A1(n419), .A2(n636), .ZN(n418) );
  NAND2_X1 U554 ( .A1(n587), .A2(n420), .ZN(n419) );
  INV_X1 U555 ( .A(n637), .ZN(n640) );
  NAND2_X1 U556 ( .A1(n426), .A2(n363), .ZN(n602) );
  NOR2_X2 U557 ( .A1(n423), .A2(n542), .ZN(n637) );
  INV_X1 U558 ( .A(KEYINPUT73), .ZN(n430) );
  XNOR2_X2 U559 ( .A(n437), .B(n436), .ZN(n570) );
  AND2_X1 U560 ( .A1(n438), .A2(n361), .ZN(n569) );
  XNOR2_X2 U561 ( .A(n662), .B(KEYINPUT106), .ZN(n438) );
  NOR2_X1 U562 ( .A1(n583), .A2(n582), .ZN(n591) );
  XNOR2_X2 U563 ( .A(n441), .B(KEYINPUT39), .ZN(n609) );
  NOR2_X2 U564 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X2 U565 ( .A(G116), .B(G113), .ZN(n446) );
  XNOR2_X1 U566 ( .A(n734), .B(n483), .ZN(n484) );
  XNOR2_X2 U567 ( .A(G146), .B(G125), .ZN(n489) );
  AND2_X1 U568 ( .A1(n524), .A2(G221), .ZN(n444) );
  XNOR2_X1 U569 ( .A(n456), .B(n455), .ZN(n458) );
  XNOR2_X1 U570 ( .A(n478), .B(n362), .ZN(n448) );
  INV_X1 U571 ( .A(n645), .ZN(n608) );
  XNOR2_X1 U572 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U573 ( .A(n513), .B(KEYINPUT16), .ZN(n452) );
  XNOR2_X1 U574 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U575 ( .A(n459), .B(n481), .ZN(n461) );
  XNOR2_X1 U576 ( .A(n530), .B(n477), .ZN(n540) );
  INV_X1 U577 ( .A(KEYINPUT84), .ZN(n611) );
  XNOR2_X1 U578 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U579 ( .A(n500), .B(KEYINPUT25), .ZN(n501) );
  XNOR2_X1 U580 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U581 ( .A(n622), .B(KEYINPUT88), .ZN(n623) );
  XNOR2_X1 U582 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U583 ( .A(n577), .B(n576), .ZN(n746) );
  XNOR2_X1 U584 ( .A(KEYINPUT4), .B(n527), .ZN(n735) );
  XNOR2_X1 U585 ( .A(G101), .B(n735), .ZN(n460) );
  XNOR2_X1 U586 ( .A(G146), .B(n460), .ZN(n485) );
  XOR2_X1 U587 ( .A(G119), .B(KEYINPUT90), .Z(n447) );
  NAND2_X1 U588 ( .A1(n508), .A2(G210), .ZN(n449) );
  XNOR2_X1 U589 ( .A(n450), .B(n485), .ZN(n618) );
  INV_X1 U590 ( .A(KEYINPUT19), .ZN(n471) );
  INV_X1 U591 ( .A(n489), .ZN(n454) );
  NAND2_X1 U592 ( .A1(G224), .A2(n728), .ZN(n456) );
  XNOR2_X1 U593 ( .A(KEYINPUT71), .B(n721), .ZN(n481) );
  XNOR2_X1 U594 ( .A(n465), .B(KEYINPUT75), .ZN(n469) );
  AND2_X1 U595 ( .A1(G210), .A2(n469), .ZN(n466) );
  XNOR2_X2 U596 ( .A(n468), .B(n467), .ZN(n607) );
  NAND2_X1 U597 ( .A1(G214), .A2(n469), .ZN(n647) );
  NAND2_X1 U598 ( .A1(n607), .A2(n647), .ZN(n470) );
  XOR2_X1 U599 ( .A(KEYINPUT14), .B(KEYINPUT92), .Z(n473) );
  XOR2_X1 U600 ( .A(n473), .B(n472), .Z(n474) );
  NAND2_X1 U601 ( .A1(G952), .A2(n474), .ZN(n674) );
  NOR2_X1 U602 ( .A1(G953), .A2(n674), .ZN(n564) );
  AND2_X1 U603 ( .A1(n474), .A2(G953), .ZN(n475) );
  NAND2_X1 U604 ( .A1(G902), .A2(n475), .ZN(n562) );
  NOR2_X1 U605 ( .A1(G898), .A2(n562), .ZN(n476) );
  NOR2_X1 U606 ( .A1(n662), .A2(n540), .ZN(n503) );
  NAND2_X1 U607 ( .A1(G227), .A2(n728), .ZN(n479) );
  XNOR2_X1 U608 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U609 ( .A(n485), .B(n484), .ZN(n694) );
  INV_X1 U610 ( .A(n617), .ZN(n486) );
  NAND2_X1 U611 ( .A1(G234), .A2(n486), .ZN(n487) );
  XNOR2_X1 U612 ( .A(KEYINPUT20), .B(n487), .ZN(n499) );
  NAND2_X1 U613 ( .A1(G221), .A2(n499), .ZN(n488) );
  XOR2_X1 U614 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n492) );
  NAND2_X1 U615 ( .A1(G234), .A2(n728), .ZN(n491) );
  XNOR2_X1 U616 ( .A(n492), .B(n491), .ZN(n524) );
  XOR2_X1 U617 ( .A(KEYINPUT24), .B(G110), .Z(n495) );
  XNOR2_X1 U618 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U619 ( .A(n496), .B(KEYINPUT23), .Z(n497) );
  XNOR2_X1 U620 ( .A(n498), .B(n497), .ZN(n712) );
  NOR2_X1 U621 ( .A1(G902), .A2(n712), .ZN(n502) );
  NAND2_X1 U622 ( .A1(G217), .A2(n499), .ZN(n500) );
  NAND2_X1 U623 ( .A1(n503), .A2(n578), .ZN(n504) );
  XNOR2_X1 U624 ( .A(n504), .B(KEYINPUT96), .ZN(n625) );
  NOR2_X1 U625 ( .A1(n659), .A2(n658), .ZN(n537) );
  NAND2_X1 U626 ( .A1(n662), .A2(n537), .ZN(n667) );
  NOR2_X1 U627 ( .A1(n530), .A2(n667), .ZN(n505) );
  XNOR2_X1 U628 ( .A(KEYINPUT31), .B(n505), .ZN(n642) );
  NAND2_X1 U629 ( .A1(n625), .A2(n642), .ZN(n529) );
  XNOR2_X1 U630 ( .A(KEYINPUT13), .B(G475), .ZN(n517) );
  XOR2_X1 U631 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n507) );
  XNOR2_X1 U632 ( .A(KEYINPUT11), .B(KEYINPUT99), .ZN(n506) );
  NAND2_X1 U633 ( .A1(G214), .A2(n508), .ZN(n509) );
  XNOR2_X1 U634 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U635 ( .A(n513), .B(KEYINPUT97), .ZN(n514) );
  XNOR2_X1 U636 ( .A(n515), .B(n514), .ZN(n701) );
  NOR2_X1 U637 ( .A1(G902), .A2(n701), .ZN(n516) );
  XNOR2_X1 U638 ( .A(n519), .B(n518), .ZN(n523) );
  XNOR2_X1 U639 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U640 ( .A(n523), .B(n522), .Z(n526) );
  NAND2_X1 U641 ( .A1(G217), .A2(n524), .ZN(n525) );
  XOR2_X1 U642 ( .A(G478), .B(n528), .Z(n542) );
  NAND2_X1 U643 ( .A1(n529), .A2(n587), .ZN(n535) );
  NOR2_X1 U644 ( .A1(n543), .A2(n542), .ZN(n574) );
  OR2_X2 U645 ( .A1(n530), .A2(n365), .ZN(n531) );
  XNOR2_X1 U646 ( .A(KEYINPUT6), .B(n533), .ZN(n596) );
  NOR2_X1 U647 ( .A1(n596), .A2(n549), .ZN(n534) );
  NAND2_X1 U648 ( .A1(n364), .A2(n534), .ZN(n624) );
  NAND2_X1 U649 ( .A1(n535), .A2(n624), .ZN(n536) );
  XOR2_X1 U650 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n539) );
  NAND2_X1 U651 ( .A1(n537), .A2(n596), .ZN(n538) );
  XNOR2_X1 U652 ( .A(n541), .B(KEYINPUT34), .ZN(n545) );
  NAND2_X1 U653 ( .A1(n543), .A2(n542), .ZN(n589) );
  XOR2_X1 U654 ( .A(n589), .B(KEYINPUT78), .Z(n544) );
  NAND2_X1 U655 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U656 ( .A1(n555), .A2(KEYINPUT44), .ZN(n547) );
  INV_X1 U657 ( .A(n549), .ZN(n656) );
  NOR2_X1 U658 ( .A1(n596), .A2(n656), .ZN(n552) );
  NAND2_X1 U659 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U660 ( .A1(n556), .A2(KEYINPUT44), .ZN(n557) );
  NOR2_X1 U661 ( .A1(G900), .A2(n562), .ZN(n563) );
  NOR2_X1 U662 ( .A1(n564), .A2(n563), .ZN(n580) );
  INV_X1 U663 ( .A(n655), .ZN(n565) );
  NOR2_X1 U664 ( .A1(n580), .A2(n565), .ZN(n566) );
  XOR2_X1 U665 ( .A(KEYINPUT70), .B(n566), .Z(n567) );
  XNOR2_X1 U666 ( .A(KEYINPUT28), .B(KEYINPUT111), .ZN(n568) );
  XNOR2_X1 U667 ( .A(n569), .B(n568), .ZN(n572) );
  XNOR2_X1 U668 ( .A(KEYINPUT110), .B(n570), .ZN(n571) );
  OR2_X1 U669 ( .A1(n572), .A2(n571), .ZN(n586) );
  INV_X1 U670 ( .A(n607), .ZN(n597) );
  XNOR2_X1 U671 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n573) );
  NAND2_X1 U672 ( .A1(n646), .A2(n647), .ZN(n650) );
  INV_X1 U673 ( .A(n574), .ZN(n649) );
  NOR2_X1 U674 ( .A1(n650), .A2(n649), .ZN(n575) );
  XNOR2_X1 U675 ( .A(n575), .B(KEYINPUT41), .ZN(n675) );
  NOR2_X1 U676 ( .A1(n586), .A2(n675), .ZN(n577) );
  XNOR2_X1 U677 ( .A(n578), .B(KEYINPUT109), .ZN(n579) );
  XNOR2_X1 U678 ( .A(KEYINPUT67), .B(KEYINPUT47), .ZN(n588) );
  NOR2_X1 U679 ( .A1(n597), .A2(n589), .ZN(n590) );
  NAND2_X1 U680 ( .A1(n591), .A2(n590), .ZN(n636) );
  AND2_X1 U681 ( .A1(KEYINPUT47), .A2(n651), .ZN(n592) );
  NOR2_X1 U682 ( .A1(KEYINPUT82), .A2(n592), .ZN(n593) );
  NAND2_X1 U683 ( .A1(n651), .A2(KEYINPUT82), .ZN(n594) );
  NAND2_X1 U684 ( .A1(n594), .A2(n638), .ZN(n595) );
  NAND2_X1 U685 ( .A1(n595), .A2(KEYINPUT47), .ZN(n600) );
  XNOR2_X1 U686 ( .A(n602), .B(KEYINPUT107), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n603), .A2(n659), .ZN(n604) );
  XNOR2_X1 U688 ( .A(n604), .B(KEYINPUT108), .ZN(n605) );
  XOR2_X1 U689 ( .A(KEYINPUT43), .B(n605), .Z(n606) );
  NOR2_X1 U690 ( .A1(n358), .A2(n606), .ZN(n645) );
  NAND2_X1 U691 ( .A1(n609), .A2(n633), .ZN(n610) );
  XNOR2_X1 U692 ( .A(n610), .B(KEYINPUT114), .ZN(n751) );
  NAND2_X1 U693 ( .A1(KEYINPUT2), .A2(n751), .ZN(n613) );
  XOR2_X1 U694 ( .A(KEYINPUT80), .B(n613), .Z(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n359), .A2(G472), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n618), .B(KEYINPUT62), .ZN(n619) );
  XNOR2_X1 U698 ( .A(n620), .B(n619), .ZN(n621) );
  INV_X1 U699 ( .A(KEYINPUT63), .ZN(n622) );
  XNOR2_X1 U700 ( .A(G101), .B(n624), .ZN(G3) );
  BUF_X1 U701 ( .A(n625), .Z(n627) );
  NOR2_X1 U702 ( .A1(n627), .A2(n640), .ZN(n626) );
  XOR2_X1 U703 ( .A(G104), .B(n626), .Z(G6) );
  INV_X1 U704 ( .A(n633), .ZN(n643) );
  NOR2_X1 U705 ( .A1(n643), .A2(n627), .ZN(n631) );
  XOR2_X1 U706 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n629) );
  XNOR2_X1 U707 ( .A(G107), .B(KEYINPUT27), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n631), .B(n630), .ZN(G9) );
  XNOR2_X1 U710 ( .A(n632), .B(G110), .ZN(G12) );
  XOR2_X1 U711 ( .A(G128), .B(KEYINPUT29), .Z(n635) );
  NAND2_X1 U712 ( .A1(n638), .A2(n633), .ZN(n634) );
  XNOR2_X1 U713 ( .A(n635), .B(n634), .ZN(G30) );
  XNOR2_X1 U714 ( .A(G143), .B(n636), .ZN(G45) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n639), .B(G146), .ZN(G48) );
  NOR2_X1 U717 ( .A1(n640), .A2(n642), .ZN(n641) );
  XOR2_X1 U718 ( .A(G113), .B(n641), .Z(G15) );
  NOR2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U720 ( .A(G116), .B(n644), .Z(G18) );
  XOR2_X1 U721 ( .A(G140), .B(n645), .Z(G42) );
  NOR2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n653) );
  NOR2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U726 ( .A1(n676), .A2(n654), .ZN(n671) );
  NOR2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U728 ( .A(KEYINPUT49), .B(n657), .ZN(n665) );
  XOR2_X1 U729 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n661) );
  NAND2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U735 ( .A(KEYINPUT51), .B(n668), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n669), .A2(n675), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(KEYINPUT52), .ZN(n673) );
  NOR2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n678) );
  NOR2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n684) );
  XNOR2_X1 U742 ( .A(KEYINPUT81), .B(KEYINPUT2), .ZN(n680) );
  NAND2_X1 U743 ( .A1(n740), .A2(n729), .ZN(n679) );
  NAND2_X1 U744 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X1 U745 ( .A1(n682), .A2(n368), .ZN(n683) );
  NAND2_X1 U746 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U747 ( .A1(G953), .A2(n685), .ZN(n686) );
  NAND2_X1 U748 ( .A1(n359), .A2(G210), .ZN(n690) );
  XOR2_X1 U749 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n687) );
  XNOR2_X1 U750 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U751 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U752 ( .A(KEYINPUT118), .B(KEYINPUT56), .ZN(n692) );
  XNOR2_X1 U753 ( .A(n692), .B(KEYINPUT86), .ZN(n693) );
  XNOR2_X1 U754 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n696) );
  XNOR2_X1 U755 ( .A(n694), .B(KEYINPUT57), .ZN(n695) );
  XNOR2_X1 U756 ( .A(n696), .B(n695), .ZN(n698) );
  NAND2_X1 U757 ( .A1(n713), .A2(G469), .ZN(n697) );
  NAND2_X1 U758 ( .A1(n359), .A2(G475), .ZN(n703) );
  XOR2_X1 U759 ( .A(KEYINPUT59), .B(KEYINPUT120), .Z(n700) );
  XNOR2_X1 U760 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U761 ( .A(KEYINPUT60), .B(KEYINPUT66), .ZN(n705) );
  XNOR2_X1 U762 ( .A(n706), .B(n705), .ZN(G60) );
  NAND2_X1 U763 ( .A1(n713), .A2(G478), .ZN(n710) );
  INV_X1 U764 ( .A(KEYINPUT121), .ZN(n707) );
  NOR2_X1 U765 ( .A1(n717), .A2(n711), .ZN(G63) );
  XNOR2_X1 U766 ( .A(n712), .B(KEYINPUT122), .ZN(n715) );
  NAND2_X1 U767 ( .A1(G217), .A2(n713), .ZN(n714) );
  BUF_X1 U768 ( .A(n718), .Z(n719) );
  XOR2_X1 U769 ( .A(n719), .B(KEYINPUT124), .Z(n720) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U771 ( .A(n722), .B(G101), .ZN(n724) );
  NOR2_X1 U772 ( .A1(n728), .A2(G898), .ZN(n723) );
  NOR2_X1 U773 ( .A1(n724), .A2(n723), .ZN(n733) );
  XOR2_X1 U774 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n726) );
  NAND2_X1 U775 ( .A1(G224), .A2(G953), .ZN(n725) );
  XNOR2_X1 U776 ( .A(n726), .B(n725), .ZN(n727) );
  NAND2_X1 U777 ( .A1(n727), .A2(G898), .ZN(n731) );
  NAND2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U780 ( .A(n733), .B(n732), .ZN(G69) );
  XNOR2_X1 U781 ( .A(n734), .B(n735), .ZN(n736) );
  XOR2_X1 U782 ( .A(KEYINPUT126), .B(n741), .Z(n737) );
  XNOR2_X1 U783 ( .A(G227), .B(n737), .ZN(n738) );
  NAND2_X1 U784 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U785 ( .A1(n739), .A2(G953), .ZN(n745) );
  XOR2_X1 U786 ( .A(n741), .B(n740), .Z(n742) );
  NOR2_X1 U787 ( .A1(G953), .A2(n742), .ZN(n743) );
  XNOR2_X1 U788 ( .A(KEYINPUT125), .B(n743), .ZN(n744) );
  NAND2_X1 U789 ( .A1(n745), .A2(n744), .ZN(G72) );
  XOR2_X1 U790 ( .A(n746), .B(n351), .Z(G39) );
  XOR2_X1 U791 ( .A(G125), .B(KEYINPUT37), .Z(n747) );
  XNOR2_X1 U792 ( .A(n748), .B(n747), .ZN(G27) );
  XOR2_X1 U793 ( .A(n555), .B(G122), .Z(G24) );
  XNOR2_X1 U794 ( .A(n749), .B(G119), .ZN(G21) );
  XOR2_X1 U795 ( .A(n750), .B(G131), .Z(G33) );
  XNOR2_X1 U796 ( .A(G134), .B(n751), .ZN(G36) );
endmodule

