//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n193), .A2(KEYINPUT64), .A3(G143), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT64), .B1(new_n193), .B2(G143), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n190), .B(new_n192), .C1(new_n194), .C2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n190), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT0), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(new_n191), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n190), .B(new_n206), .C1(new_n194), .C2(new_n195), .ZN(new_n207));
  INV_X1    g021(.A(new_n206), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n191), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n200), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n204), .B1(new_n203), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G953), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G224), .ZN(new_n214));
  XOR2_X1   g028(.A(new_n214), .B(KEYINPUT79), .Z(new_n215));
  XNOR2_X1  g029(.A(new_n212), .B(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT5), .ZN(new_n217));
  INV_X1    g031(.A(G119), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G116), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n220));
  INV_X1    g034(.A(G116), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G119), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(G119), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n218), .A2(KEYINPUT67), .A3(G116), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(G113), .B(new_n219), .C1(new_n225), .C2(new_n217), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT2), .B(G113), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G107), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G104), .ZN(new_n231));
  INV_X1    g045(.A(G104), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(G107), .ZN(new_n233));
  OAI21_X1  g047(.A(G101), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n230), .A3(G104), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n235), .A2(new_n230), .A3(KEYINPUT75), .A4(G104), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n231), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G101), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT3), .B1(new_n232), .B2(G107), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT74), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(KEYINPUT74), .B(KEYINPUT3), .C1(new_n232), .C2(G107), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n229), .A2(new_n234), .A3(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n240), .A2(new_n241), .A3(new_n246), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n241), .B1(new_n240), .B2(new_n246), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n231), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT75), .B1(new_n233), .B2(new_n235), .ZN(new_n254));
  INV_X1    g068(.A(new_n239), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n245), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n230), .A2(G104), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT74), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n251), .B(G101), .C1(new_n256), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n225), .A2(new_n227), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n228), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n248), .B1(new_n252), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g079(.A(G110), .B(G122), .Z(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n250), .A2(new_n251), .B1(new_n228), .B2(new_n262), .ZN(new_n268));
  OAI21_X1  g082(.A(G101), .B1(new_n256), .B2(new_n260), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT4), .A3(new_n247), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n266), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n248), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n267), .A2(KEYINPUT6), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT78), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n271), .B2(new_n248), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n247), .A2(new_n234), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n268), .A2(new_n270), .B1(new_n279), .B2(new_n229), .ZN(new_n280));
  NOR4_X1   g094(.A1(new_n280), .A2(KEYINPUT78), .A3(KEYINPUT6), .A4(new_n272), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n216), .B(new_n274), .C1(new_n278), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT80), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n265), .A2(new_n277), .A3(new_n266), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT78), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n276), .A2(new_n275), .A3(new_n277), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT80), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n216), .A4(new_n274), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G210), .B1(G237), .B2(G902), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(KEYINPUT81), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n214), .A2(KEYINPUT7), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n212), .B(new_n294), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n279), .A2(new_n229), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n296), .A2(new_n248), .ZN(new_n297));
  XOR2_X1   g111(.A(new_n266), .B(KEYINPUT8), .Z(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n295), .B(new_n273), .C1(new_n297), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n290), .A2(new_n293), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n277), .B1(new_n265), .B2(new_n266), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n285), .A2(new_n286), .B1(new_n273), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n288), .B1(new_n306), .B2(new_n216), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n282), .A2(KEYINPUT80), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n303), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n292), .B(KEYINPUT82), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n304), .A2(KEYINPUT83), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT83), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n290), .A2(new_n312), .A3(new_n293), .A4(new_n303), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n188), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT11), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  AOI22_X1  g131(.A1(KEYINPUT65), .A2(new_n316), .B1(new_n317), .B2(G137), .ZN(new_n318));
  OAI22_X1  g132(.A1(KEYINPUT65), .A2(new_n316), .B1(new_n317), .B2(G137), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT65), .ZN(new_n320));
  INV_X1    g134(.A(G137), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT11), .A4(G134), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G131), .ZN(new_n324));
  INV_X1    g138(.A(G131), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n318), .A2(new_n319), .A3(new_n325), .A4(new_n322), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n211), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n193), .A2(G143), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT64), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n189), .B2(G146), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n193), .A2(KEYINPUT64), .A3(G143), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n332), .A2(new_n192), .B1(new_n198), .B2(new_n200), .ZN(new_n333));
  AND4_X1   g147(.A1(new_n325), .A2(new_n318), .A3(new_n319), .A4(new_n322), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n317), .A2(G137), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n321), .A2(G134), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n325), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n333), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n263), .B1(new_n327), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n324), .A2(new_n326), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n207), .A2(new_n210), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n228), .A2(new_n262), .ZN(new_n343));
  INV_X1    g157(.A(new_n337), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n202), .A2(new_n326), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n315), .B1(new_n339), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n346), .A2(new_n315), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT26), .B(G101), .Z(new_n349));
  NOR2_X1   g163(.A1(G237), .A2(G953), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G210), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n349), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT29), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n347), .A2(new_n348), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT70), .B1(new_n356), .B2(G902), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n343), .B1(new_n342), .B2(new_n345), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n346), .A2(new_n315), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n354), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n364));
  NAND2_X1  g178(.A1(KEYINPUT66), .A2(KEYINPUT30), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT66), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n365), .B(new_n368), .C1(new_n327), .C2(new_n338), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n342), .A2(new_n366), .A3(new_n367), .A4(new_n345), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n359), .B1(new_n371), .B2(new_n263), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n363), .B(new_n364), .C1(new_n372), .C2(new_n354), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT70), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT28), .B1(new_n359), .B2(new_n360), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n362), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n374), .B(new_n301), .C1(new_n376), .C2(new_n355), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n357), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G472), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT71), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(KEYINPUT71), .A3(G472), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n354), .B1(new_n361), .B2(new_n362), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n371), .A2(new_n263), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n354), .A3(new_n346), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT31), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n372), .A2(KEYINPUT31), .A3(new_n354), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n383), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(G472), .A2(G902), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT32), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT31), .B1(new_n372), .B2(new_n354), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n343), .B1(new_n369), .B2(new_n370), .ZN(new_n394));
  INV_X1    g208(.A(new_n354), .ZN(new_n395));
  NOR4_X1   g209(.A1(new_n394), .A2(new_n386), .A3(new_n395), .A4(new_n359), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n361), .A2(new_n362), .ZN(new_n397));
  OAI22_X1  g211(.A1(new_n393), .A2(new_n396), .B1(new_n397), .B2(new_n354), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT32), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(new_n390), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n381), .A2(new_n382), .B1(new_n392), .B2(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(G125), .A2(G140), .ZN(new_n402));
  NOR2_X1   g216(.A1(G125), .A2(G140), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT16), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OR3_X1    g218(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(G146), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT72), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n405), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n193), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n407), .B(new_n409), .ZN(new_n410));
  OR3_X1    g224(.A1(new_n218), .A2(KEYINPUT23), .A3(G128), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT23), .B1(new_n218), .B2(G128), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n411), .A2(new_n412), .B1(new_n218), .B2(G128), .ZN(new_n413));
  INV_X1    g227(.A(G110), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  XOR2_X1   g229(.A(G119), .B(G128), .Z(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT24), .B(G110), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n410), .B(new_n415), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n413), .A2(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n419), .A2(KEYINPUT73), .ZN(new_n420));
  INV_X1    g234(.A(G140), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n203), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(G125), .A2(G140), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n193), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n419), .A2(KEYINPUT73), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n420), .A2(new_n425), .A3(new_n406), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n213), .A2(G221), .A3(G234), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT22), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(G137), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n418), .A2(new_n427), .A3(new_n431), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n301), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT25), .ZN(new_n436));
  INV_X1    g250(.A(G217), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(G234), .B2(new_n301), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT25), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n433), .A2(new_n439), .A3(new_n301), .A4(new_n434), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n436), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n433), .A2(new_n434), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n438), .A2(G902), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n324), .A2(new_n326), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(KEYINPUT76), .ZN(new_n447));
  INV_X1    g261(.A(new_n198), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n196), .B1(new_n448), .B2(new_n332), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n247), .A2(new_n234), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n202), .B1(new_n247), .B2(new_n234), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT12), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT10), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n333), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n247), .A2(new_n234), .A3(new_n449), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n279), .A2(new_n456), .B1(new_n457), .B2(new_n455), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n270), .A2(new_n261), .A3(new_n341), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n446), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G110), .B(G140), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n213), .A2(G227), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n462), .B(new_n463), .Z(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n460), .A2(new_n464), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT77), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n446), .B1(new_n458), .B2(new_n459), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(KEYINPUT77), .A3(new_n464), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n473), .A3(G469), .ZN(new_n474));
  INV_X1    g288(.A(G469), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n452), .B(KEYINPUT12), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n467), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n464), .B1(new_n471), .B2(new_n460), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n475), .B(new_n301), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n475), .A2(new_n301), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n474), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT9), .B(G234), .Z(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G221), .B1(new_n484), .B2(G902), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n401), .A2(new_n445), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT15), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G478), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT88), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(G122), .ZN(new_n492));
  INV_X1    g306(.A(G122), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT88), .ZN(new_n494));
  OAI21_X1  g308(.A(G116), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n493), .B2(G116), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n221), .A2(KEYINPUT89), .A3(G122), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n495), .B1(KEYINPUT14), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT92), .B1(new_n499), .B2(KEYINPUT14), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n502), .B(new_n503), .C1(new_n497), .C2(new_n498), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n500), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT93), .B1(new_n505), .B2(new_n230), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n497), .A2(new_n498), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n493), .A2(KEYINPUT88), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n491), .A2(G122), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n221), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT90), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n495), .A2(new_n499), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT90), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n230), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n510), .B1(new_n507), .B2(new_n503), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n499), .A2(KEYINPUT14), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n502), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n499), .A2(KEYINPUT92), .A3(KEYINPUT14), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(G107), .ZN(new_n523));
  XNOR2_X1  g337(.A(G128), .B(G143), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(new_n317), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n317), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n526), .B1(new_n525), .B2(new_n527), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n506), .A2(new_n516), .A3(new_n523), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n524), .A2(KEYINPUT13), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n191), .A2(KEYINPUT13), .A3(G143), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(new_n317), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n532), .A2(new_n534), .B1(new_n317), .B2(new_n524), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n513), .A2(new_n515), .A3(new_n230), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n511), .A2(new_n512), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n514), .A2(KEYINPUT90), .ZN(new_n538));
  AOI21_X1  g352(.A(G107), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n535), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n484), .A2(new_n437), .A3(G953), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n531), .A2(new_n540), .A3(new_n542), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n490), .B1(new_n546), .B2(new_n301), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n531), .A2(new_n540), .A3(new_n542), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n542), .B1(new_n531), .B2(new_n540), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n301), .B(new_n490), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n488), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n301), .B1(new_n548), .B2(new_n549), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n489), .A3(G478), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(KEYINPUT94), .A3(new_n550), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n402), .B2(new_n403), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n422), .A2(KEYINPUT19), .A3(new_n423), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n193), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n406), .ZN(new_n561));
  INV_X1    g375(.A(G237), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n213), .A3(G214), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n189), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n350), .A2(G143), .A3(G214), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G131), .ZN(new_n567));
  AND4_X1   g381(.A1(G143), .A2(new_n562), .A3(new_n213), .A4(G214), .ZN(new_n568));
  AOI21_X1  g382(.A(G143), .B1(new_n350), .B2(G214), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n325), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n561), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n424), .B(G146), .ZN(new_n573));
  NAND2_X1  g387(.A1(KEYINPUT18), .A2(G131), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT84), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n566), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n574), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n570), .A2(KEYINPUT84), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n573), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT85), .B1(new_n572), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n573), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n577), .B1(new_n570), .B2(KEYINPUT84), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n566), .A2(new_n575), .A3(new_n574), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT85), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n571), .A2(new_n567), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n560), .A2(new_n406), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n584), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(G113), .B(G122), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(new_n232), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n580), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT86), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n591), .B(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n566), .A2(KEYINPUT17), .A3(G131), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n586), .B2(KEYINPUT17), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n584), .B(new_n595), .C1(new_n410), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(G475), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n301), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT87), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT20), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(G475), .B1(new_n593), .B2(new_n598), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT20), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n301), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n605), .B2(new_n301), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n607), .B1(new_n608), .B2(new_n602), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n410), .A2(new_n597), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n592), .B1(new_n610), .B2(new_n579), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n598), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n301), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n604), .A2(new_n609), .B1(G475), .B2(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n213), .A2(G952), .ZN(new_n615));
  NAND2_X1  g429(.A1(G234), .A2(G237), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT21), .B(G898), .Z(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n616), .A2(G902), .A3(G953), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n618), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n556), .A2(new_n614), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n314), .A2(new_n487), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G101), .ZN(G3));
  AOI21_X1  g442(.A(new_n293), .B1(new_n290), .B2(new_n303), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n188), .B1(new_n630), .B2(new_n304), .ZN(new_n631));
  OAI21_X1  g445(.A(G472), .B1(new_n389), .B2(G902), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n398), .A2(new_n390), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n482), .A2(new_n632), .A3(new_n633), .A4(new_n485), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n445), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n613), .A2(G475), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n606), .A2(new_n599), .A3(new_n600), .A4(new_n301), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n601), .A2(KEYINPUT20), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(KEYINPUT87), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n636), .B1(new_n639), .B2(new_n603), .ZN(new_n640));
  INV_X1    g454(.A(G478), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n546), .A2(new_n641), .A3(new_n301), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT33), .B1(new_n542), .B2(KEYINPUT95), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n548), .B2(new_n549), .ZN(new_n645));
  INV_X1    g459(.A(new_n644), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n544), .A2(new_n545), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n641), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n641), .A2(new_n301), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n643), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n640), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n623), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n631), .A2(new_n635), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT96), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n653), .B(new_n655), .ZN(G6));
  XOR2_X1   g470(.A(new_n623), .B(KEYINPUT98), .Z(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n292), .B(new_n302), .C1(new_n283), .C2(new_n289), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n187), .B(new_n658), .C1(new_n629), .C2(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n637), .A2(new_n608), .A3(KEYINPUT97), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT97), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n638), .B2(new_n607), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n664), .A2(new_n636), .A3(new_n555), .A4(new_n552), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n635), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  INV_X1    g483(.A(new_n634), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n432), .A2(KEYINPUT36), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT99), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n428), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n443), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n441), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n314), .A2(new_n626), .A3(new_n670), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT37), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n414), .ZN(G12));
  OAI211_X1 g492(.A(new_n187), .B(new_n675), .C1(new_n629), .C2(new_n659), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n621), .A2(G900), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n617), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n665), .A2(new_n486), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n382), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT71), .B1(new_n378), .B2(G472), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n389), .A2(KEYINPUT32), .A3(new_n391), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n399), .B1(new_n398), .B2(new_n390), .ZN(new_n688));
  OAI22_X1  g502(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n680), .A2(new_n684), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  INV_X1    g505(.A(G472), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n395), .B1(new_n359), .B2(new_n360), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n385), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n692), .B1(new_n694), .B2(new_n301), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n392), .B2(new_n400), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n675), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n682), .B(KEYINPUT100), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT39), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n482), .A2(new_n485), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT101), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n482), .A2(new_n702), .A3(new_n485), .A4(new_n699), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n701), .A2(KEYINPUT40), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT40), .B1(new_n701), .B2(new_n703), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n697), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n304), .A2(KEYINPUT83), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n309), .A2(new_n310), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n313), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT38), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n311), .A2(KEYINPUT38), .A3(new_n313), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n556), .A2(new_n614), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n711), .A2(new_n712), .A3(new_n187), .A4(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n706), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n189), .ZN(G45));
  NOR3_X1   g530(.A1(new_n651), .A2(new_n486), .A3(new_n683), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n680), .A2(new_n689), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  OAI21_X1  g533(.A(new_n301), .B1(new_n477), .B2(new_n478), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n475), .A2(KEYINPUT102), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n485), .A3(new_n724), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n401), .A2(new_n725), .A3(new_n445), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n631), .A3(new_n652), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT103), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT41), .B(G113), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  NAND2_X1  g544(.A1(new_n666), .A2(new_n726), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G116), .ZN(G18));
  INV_X1    g546(.A(new_n725), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n680), .A2(new_n626), .A3(new_n689), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  NAND2_X1  g549(.A1(new_n632), .A2(KEYINPUT105), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n376), .A2(KEYINPUT104), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n376), .A2(KEYINPUT104), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n395), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n393), .B2(new_n396), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n390), .ZN(new_n741));
  INV_X1    g555(.A(new_n445), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n743), .B(G472), .C1(new_n389), .C2(G902), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n736), .A2(new_n741), .A3(new_n742), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n725), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT106), .B1(new_n556), .B2(new_n614), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n640), .A2(new_n748), .A3(new_n555), .A4(new_n552), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n660), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n746), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT107), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  AND4_X1   g568(.A1(new_n675), .A2(new_n736), .A3(new_n741), .A4(new_n744), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n651), .A2(new_n683), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n631), .A3(new_n756), .A4(new_n733), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(KEYINPUT42), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n707), .A2(new_n708), .A3(new_n187), .A4(new_n313), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n762), .A2(new_n651), .A3(new_n683), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n761), .B1(new_n763), .B2(new_n487), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n311), .A2(new_n187), .A3(new_n313), .A4(new_n682), .ZN(new_n765));
  INV_X1    g579(.A(new_n486), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n689), .A2(new_n742), .A3(new_n766), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n765), .A2(new_n767), .A3(new_n651), .A4(new_n760), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT109), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  NOR2_X1   g585(.A1(new_n401), .A2(new_n445), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n762), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n684), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n460), .A2(KEYINPUT77), .A3(new_n464), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT77), .B1(new_n460), .B2(new_n464), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n778), .A2(new_n779), .A3(new_n470), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n464), .B1(new_n454), .B2(new_n460), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n466), .A2(new_n473), .A3(KEYINPUT45), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(G469), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n782), .A2(KEYINPUT110), .A3(new_n783), .A4(G469), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n480), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT46), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT46), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n479), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(KEYINPUT111), .A3(new_n485), .A4(new_n699), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n479), .B1(new_n788), .B2(KEYINPUT46), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n794), .B(new_n480), .C1(new_n786), .C2(new_n787), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n485), .B(new_n699), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n632), .A2(new_n633), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n650), .A2(new_n614), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT43), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n650), .A2(new_n614), .A3(KEYINPUT43), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(new_n675), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n762), .B1(new_n807), .B2(KEYINPUT44), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT112), .B1(new_n807), .B2(KEYINPUT44), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n675), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT44), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n799), .A2(new_n808), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT113), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  OAI21_X1  g631(.A(new_n485), .B1(new_n793), .B2(new_n795), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(KEYINPUT47), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n819), .A2(KEYINPUT47), .ZN(new_n823));
  OAI221_X1 g637(.A(new_n485), .B1(new_n820), .B2(new_n823), .C1(new_n793), .C2(new_n795), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n689), .A2(new_n742), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n822), .A2(new_n824), .A3(new_n763), .A4(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  OAI211_X1 g641(.A(new_n689), .B(new_n680), .C1(new_n684), .C2(new_n717), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n696), .A2(new_n675), .A3(new_n683), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n750), .A2(new_n766), .A3(new_n631), .A4(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n830), .A3(new_n757), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT116), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n828), .A2(new_n830), .A3(KEYINPUT52), .A4(new_n757), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n835), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n833), .A3(KEYINPUT116), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n727), .A2(new_n752), .A3(new_n734), .A4(new_n731), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n634), .A2(new_n651), .A3(new_n445), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n314), .A2(new_n658), .A3(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n676), .A2(new_n627), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n554), .A2(new_n550), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n640), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n709), .A2(new_n187), .A3(new_n658), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT115), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n314), .A2(new_n849), .A3(new_n658), .A4(new_n846), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n850), .A3(new_n635), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n840), .A2(new_n843), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n651), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n741), .A3(new_n736), .A4(new_n744), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n689), .A2(new_n636), .A3(new_n845), .A4(new_n664), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n762), .A2(new_n683), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n766), .A3(new_n675), .A4(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n775), .B(new_n858), .C1(new_n764), .C2(new_n768), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT53), .B1(new_n839), .B2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n848), .A2(new_n850), .A3(new_n635), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n727), .A2(new_n734), .A3(new_n752), .A4(new_n731), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n676), .A2(new_n627), .A3(new_n842), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n859), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n833), .A2(new_n835), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n861), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n837), .B1(KEYINPUT116), .B2(new_n833), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n837), .A2(new_n833), .A3(KEYINPUT116), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n860), .B(KEYINPUT53), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n868), .A2(new_n870), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n617), .B1(new_n804), .B2(new_n805), .ZN(new_n879));
  INV_X1    g693(.A(new_n745), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n631), .A3(new_n733), .A4(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n872), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n880), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n822), .A2(new_n824), .ZN(new_n884));
  INV_X1    g698(.A(new_n724), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n722), .ZN(new_n886));
  INV_X1    g700(.A(new_n485), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n762), .B(new_n883), .C1(new_n884), .C2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n890));
  OR3_X1    g704(.A1(new_n762), .A2(new_n890), .A3(new_n725), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n890), .B1(new_n762), .B2(new_n725), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n891), .A2(new_n618), .A3(new_n892), .ZN(new_n893));
  OR3_X1    g707(.A1(new_n643), .A2(new_n648), .A3(new_n649), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n696), .A2(new_n742), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n893), .A2(new_n614), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n804), .A2(new_n805), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(new_n755), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n711), .A2(new_n712), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n188), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n879), .A2(new_n733), .A3(new_n880), .ZN(new_n901));
  OR3_X1    g715(.A1(new_n900), .A2(KEYINPUT50), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT50), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n896), .A2(new_n898), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n906));
  OAI22_X1  g720(.A1(new_n889), .A2(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n893), .A2(new_n853), .A3(new_n895), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n905), .B(new_n906), .C1(new_n889), .C2(new_n904), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n892), .A2(new_n618), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(new_n772), .A3(new_n897), .A4(new_n891), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT120), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n893), .A2(new_n915), .A3(new_n772), .A4(new_n897), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(KEYINPUT48), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(KEYINPUT121), .B(KEYINPUT48), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n914), .A2(new_n916), .A3(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n920), .A2(new_n615), .A3(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n923), .ZN(new_n924));
  OAI22_X1  g738(.A1(new_n882), .A2(new_n924), .B1(G952), .B2(G953), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n887), .B(new_n802), .C1(new_n711), .C2(new_n712), .ZN(new_n926));
  INV_X1    g740(.A(new_n886), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n927), .A2(KEYINPUT49), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n188), .B1(new_n927), .B2(KEYINPUT49), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n926), .A2(new_n895), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n930), .ZN(G75));
  NOR2_X1   g745(.A1(new_n213), .A2(G952), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT122), .Z(new_n933));
  XNOR2_X1  g747(.A(new_n306), .B(new_n216), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT55), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n935), .A2(KEYINPUT56), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n301), .B1(new_n875), .B2(new_n876), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(new_n310), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n292), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI211_X1 g755(.A(new_n933), .B(new_n938), .C1(new_n941), .C2(new_n935), .ZN(G51));
  XNOR2_X1  g756(.A(new_n480), .B(KEYINPUT57), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n875), .A2(new_n877), .A3(new_n876), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n477), .A2(new_n478), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n937), .A2(new_n786), .A3(new_n787), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n932), .B1(new_n948), .B2(new_n949), .ZN(G54));
  NAND3_X1  g764(.A1(new_n937), .A2(KEYINPUT58), .A3(G475), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n598), .A3(new_n593), .ZN(new_n952));
  INV_X1    g766(.A(new_n932), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n937), .A2(KEYINPUT58), .A3(G475), .A4(new_n599), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G60));
  AND2_X1   g769(.A1(new_n645), .A2(new_n647), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n649), .B(KEYINPUT59), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n956), .B(new_n958), .C1(new_n944), .C2(new_n945), .ZN(new_n959));
  INV_X1    g773(.A(new_n933), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n957), .B1(new_n872), .B2(new_n878), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n959), .B(new_n960), .C1(new_n961), .C2(new_n956), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(G63));
  NAND2_X1  g777(.A1(new_n875), .A2(new_n876), .ZN(new_n964));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT123), .Z(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT60), .Z(new_n967));
  AOI21_X1  g781(.A(new_n442), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n967), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n875), .B2(new_n876), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n933), .B1(new_n972), .B2(new_n673), .ZN(new_n973));
  OAI21_X1  g787(.A(KEYINPUT124), .B1(new_n972), .B2(new_n442), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n970), .A2(KEYINPUT61), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n964), .A2(new_n673), .A3(new_n967), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n960), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n976), .B1(new_n978), .B2(new_n968), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n975), .A2(new_n979), .ZN(G66));
  INV_X1    g794(.A(G224), .ZN(new_n981));
  OAI21_X1  g795(.A(G953), .B1(new_n620), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n865), .B2(G953), .ZN(new_n983));
  INV_X1    g797(.A(G898), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n306), .B1(new_n984), .B2(G953), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT125), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n983), .B(new_n986), .ZN(G69));
  AOI21_X1  g801(.A(new_n213), .B1(G227), .B2(G900), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT127), .Z(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n815), .A2(new_n769), .A3(new_n826), .ZN(new_n993));
  INV_X1    g807(.A(new_n775), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n828), .A2(new_n757), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n773), .B1(new_n792), .B2(new_n798), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n750), .A2(new_n631), .ZN(new_n997));
  AOI211_X1 g811(.A(new_n994), .B(new_n995), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n993), .A2(new_n213), .A3(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n558), .A2(new_n559), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n371), .B(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(G900), .B2(G953), .ZN(new_n1003));
  INV_X1    g817(.A(new_n995), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n1004), .B(KEYINPUT62), .C1(new_n706), .C2(new_n714), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n715), .B2(new_n995), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n651), .B1(new_n640), .B2(new_n845), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n774), .A2(new_n703), .A3(new_n701), .A4(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n815), .A2(new_n1008), .A3(new_n826), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n213), .ZN(new_n1012));
  AOI22_X1  g826(.A1(new_n999), .A2(new_n1003), .B1(new_n1012), .B2(new_n1002), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n988), .A2(new_n989), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n992), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1014), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1003), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n996), .A2(new_n997), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1018), .A2(new_n775), .A3(new_n1004), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n815), .A2(new_n769), .A3(new_n826), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1017), .B1(new_n1021), .B2(new_n213), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1001), .B1(new_n1011), .B2(new_n213), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1016), .B(new_n991), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1015), .A2(new_n1024), .ZN(G72));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  INV_X1    g841(.A(new_n385), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n372), .A2(new_n354), .ZN(new_n1029));
  OAI221_X1 g843(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .C1(new_n861), .C2(new_n871), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1027), .B1(new_n1011), .B2(new_n852), .ZN(new_n1031));
  INV_X1    g845(.A(new_n372), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1031), .A2(new_n354), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1030), .A2(new_n953), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1021), .A2(new_n865), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n354), .B1(new_n1035), .B2(new_n1027), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1034), .B1(new_n372), .B2(new_n1036), .ZN(G57));
endmodule


