//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G224), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n189), .A2(KEYINPUT7), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G143), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n193), .B(new_n195), .C1(new_n196), .C2(new_n192), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT68), .B(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n192), .A2(G143), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(new_n196), .B2(new_n192), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n191), .B(new_n197), .C1(new_n200), .C2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT80), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT82), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n209), .A3(new_n192), .ZN(new_n210));
  INV_X1    g024(.A(new_n201), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n198), .A2(new_n199), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n215), .A3(new_n191), .A4(new_n197), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n204), .A2(new_n205), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n207), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n218), .B1(new_n220), .B2(new_n193), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT0), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT65), .B1(new_n222), .B2(new_n194), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n210), .B2(new_n211), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n225), .A2(KEYINPUT0), .A3(G128), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n221), .B1(new_n228), .B2(new_n218), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G125), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n217), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n204), .A2(new_n216), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT82), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n190), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n230), .A3(new_n190), .ZN(new_n235));
  INV_X1    g049(.A(G113), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT2), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT2), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G113), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G116), .B(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G119), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G116), .ZN(new_n245));
  INV_X1    g059(.A(G116), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G119), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT69), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n241), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT5), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n246), .A2(G119), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT5), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n236), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n243), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G104), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT3), .B1(new_n257), .B2(G107), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g073(.A(G107), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(G104), .ZN(new_n261));
  INV_X1    g075(.A(G101), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n257), .A2(G107), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n258), .A2(new_n261), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n257), .A2(G107), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n260), .A2(G104), .ZN(new_n266));
  OAI21_X1  g080(.A(G101), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n256), .A2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n245), .A2(new_n247), .A3(new_n250), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n250), .B1(new_n245), .B2(new_n247), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n237), .B(new_n239), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n242), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n258), .A2(new_n261), .A3(new_n263), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(G101), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(G101), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT4), .A3(new_n264), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n274), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(G110), .B(G122), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n270), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT81), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT5), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n255), .A2(new_n284), .B1(new_n240), .B2(new_n241), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(new_n268), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n256), .B2(new_n268), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n281), .B(KEYINPUT8), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n283), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n271), .A2(new_n272), .A3(new_n254), .ZN(new_n290));
  INV_X1    g104(.A(new_n255), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n242), .B(new_n268), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n285), .A2(new_n268), .ZN(new_n293));
  AND4_X1   g107(.A1(new_n283), .A2(new_n292), .A3(new_n288), .A4(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n235), .B(new_n282), .C1(new_n289), .C2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n187), .B1(new_n234), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT83), .ZN(new_n297));
  XOR2_X1   g111(.A(new_n281), .B(KEYINPUT79), .Z(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n270), .B2(new_n280), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT6), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n282), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n299), .A2(KEYINPUT6), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n232), .A2(new_n230), .A3(new_n189), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n189), .B1(new_n232), .B2(new_n230), .ZN(new_n304));
  OAI22_X1  g118(.A1(new_n301), .A2(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n306), .B(new_n187), .C1(new_n234), .C2(new_n295), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n297), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G210), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT84), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n297), .A2(new_n305), .A3(new_n311), .A4(new_n307), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT85), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(new_n319), .A3(new_n316), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT11), .ZN(new_n322));
  INV_X1    g136(.A(G134), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(G137), .ZN(new_n324));
  INV_X1    g138(.A(G137), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT11), .A3(G134), .ZN(new_n326));
  INV_X1    g140(.A(G131), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(G137), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n324), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n328), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n323), .A2(G137), .ZN(new_n331));
  OAI21_X1  g145(.A(G131), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n197), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n210), .A2(new_n211), .B1(new_n198), .B2(new_n199), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n329), .B(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n274), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n324), .A2(new_n326), .A3(new_n328), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G131), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT67), .A3(new_n329), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT67), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n340), .A3(G131), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n335), .B(new_n336), .C1(new_n229), .C2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n345));
  INV_X1    g159(.A(G210), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n346), .A2(G237), .A3(G953), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT26), .B(G101), .ZN(new_n349));
  XOR2_X1   g163(.A(new_n348), .B(new_n349), .Z(new_n350));
  NAND3_X1  g164(.A1(new_n343), .A2(new_n344), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n344), .B1(new_n343), .B2(new_n350), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n332), .A2(new_n329), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n214), .B2(new_n197), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n339), .A2(new_n341), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n193), .B1(new_n196), .B2(new_n192), .ZN(new_n359));
  INV_X1    g173(.A(new_n218), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI211_X1 g175(.A(new_n226), .B(new_n223), .C1(new_n210), .C2(new_n211), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(new_n360), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n357), .B1(new_n358), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n355), .B1(new_n364), .B2(KEYINPUT64), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n335), .B1(new_n229), .B2(new_n342), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT64), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT30), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n336), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT31), .B1(new_n354), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n368), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT30), .B1(new_n366), .B2(new_n367), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n274), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n343), .A2(new_n350), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT71), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n351), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT31), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n343), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n360), .B1(new_n224), .B2(new_n227), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n341), .B(new_n339), .C1(new_n380), .C2(new_n221), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n336), .B1(new_n381), .B2(new_n335), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT28), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT28), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n343), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n350), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n370), .A2(new_n378), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G472), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n187), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT32), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n383), .A2(KEYINPUT29), .A3(new_n385), .A4(new_n350), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n187), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT72), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT28), .B1(new_n364), .B2(new_n336), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n366), .A2(new_n274), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n343), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n400), .B2(KEYINPUT28), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT29), .B1(new_n401), .B2(new_n350), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n387), .B1(new_n369), .B2(new_n379), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n394), .A2(KEYINPUT72), .A3(new_n187), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n397), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G472), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n389), .A2(KEYINPUT32), .A3(new_n390), .A4(new_n187), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n393), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G217), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(G234), .B2(new_n187), .ZN(new_n411));
  INV_X1    g225(.A(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G125), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n191), .A2(G140), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT16), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT16), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n412), .A3(G125), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n192), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT73), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n415), .A2(G146), .A3(new_n417), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT68), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(G128), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n194), .A2(KEYINPUT68), .ZN(new_n425));
  OAI211_X1 g239(.A(KEYINPUT23), .B(G119), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n244), .A2(G128), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT23), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n244), .B2(G128), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G110), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n427), .B1(new_n198), .B2(new_n244), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT24), .B(G110), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n415), .A2(KEYINPUT73), .A3(G146), .A4(new_n417), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n422), .A2(new_n431), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G110), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n426), .A2(new_n437), .A3(new_n427), .A4(new_n429), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n432), .A2(new_n433), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT74), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n421), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n415), .A2(KEYINPUT74), .A3(G146), .A4(new_n417), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G125), .B(G140), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n192), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n440), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n436), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(G137), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n436), .A2(new_n447), .A3(new_n452), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT25), .B1(new_n456), .B2(new_n187), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n436), .A2(new_n447), .A3(new_n452), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n452), .B1(new_n436), .B2(new_n447), .ZN(new_n459));
  OAI211_X1 g273(.A(KEYINPUT25), .B(new_n187), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n411), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT76), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT76), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n464), .B(new_n411), .C1(new_n457), .C2(new_n461), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n456), .B(KEYINPUT77), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n411), .A2(G902), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n409), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(G237), .A2(G953), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(G143), .A3(G214), .ZN(new_n473));
  INV_X1    g287(.A(G214), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n474), .A2(G237), .A3(G953), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n473), .B1(new_n196), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(KEYINPUT87), .A3(G131), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT87), .B1(new_n476), .B2(G131), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT17), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n422), .A2(new_n435), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n476), .A2(G131), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n327), .B(new_n473), .C1(new_n196), .C2(new_n475), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n477), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n480), .B(new_n481), .C1(new_n486), .C2(KEYINPUT17), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n476), .A2(KEYINPUT18), .A3(G131), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n413), .A2(new_n414), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G146), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n446), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT18), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n492), .B(new_n473), .C1(new_n196), .C2(new_n475), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n488), .A2(new_n491), .A3(new_n485), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G113), .B(G122), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(new_n257), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n487), .A2(new_n497), .A3(new_n494), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n187), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G475), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n504));
  INV_X1    g318(.A(new_n494), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n489), .A2(KEYINPUT19), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT19), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n445), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n508), .A3(new_n192), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT88), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT88), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n506), .A2(new_n508), .A3(new_n511), .A4(new_n192), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n444), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n505), .B1(new_n513), .B2(new_n486), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n504), .B1(new_n514), .B2(new_n497), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n484), .A2(new_n485), .A3(new_n477), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n444), .A2(new_n510), .A3(new_n512), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n494), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT89), .A3(new_n498), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n515), .A2(new_n500), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT20), .ZN(new_n521));
  NOR2_X1   g335(.A1(G475), .A2(G902), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n520), .B2(new_n522), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n503), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT90), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n503), .B(new_n529), .C1(new_n523), .C2(new_n526), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n198), .A2(new_n206), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT13), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n219), .A2(G128), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n533), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT13), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT92), .A3(G134), .ZN(new_n538));
  XNOR2_X1  g352(.A(G116), .B(G122), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(new_n260), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n535), .A2(new_n531), .A3(G134), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n323), .B1(new_n534), .B2(new_n536), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n538), .B(new_n542), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n541), .A2(new_n260), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n246), .A2(KEYINPUT14), .A3(G122), .ZN(new_n549));
  INV_X1    g363(.A(new_n539), .ZN(new_n550));
  OAI211_X1 g364(.A(G107), .B(new_n549), .C1(new_n550), .C2(KEYINPUT14), .ZN(new_n551));
  INV_X1    g365(.A(new_n531), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n323), .B1(new_n552), .B2(new_n533), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n548), .B(new_n551), .C1(new_n543), .C2(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(KEYINPUT9), .B(G234), .Z(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n556), .A2(new_n410), .A3(G953), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n547), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n547), .B2(new_n554), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n187), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n561), .A3(G478), .ZN(new_n562));
  INV_X1    g376(.A(G478), .ZN(new_n563));
  OAI221_X1 g377(.A(new_n187), .B1(KEYINPUT15), .B2(new_n563), .C1(new_n558), .C2(new_n559), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G952), .ZN(new_n566));
  AOI211_X1 g380(.A(G953), .B(new_n566), .C1(G234), .C2(G237), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT21), .B(G898), .Z(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI211_X1 g383(.A(new_n187), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n528), .A2(new_n530), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G110), .B(G140), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n188), .A2(G227), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n574), .B(new_n575), .Z(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n279), .A2(new_n277), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n214), .B2(new_n197), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n578), .A2(new_n363), .B1(new_n580), .B2(new_n269), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n194), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n582));
  INV_X1    g396(.A(new_n193), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n219), .B2(G146), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n197), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n269), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n579), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n342), .B1(new_n581), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n269), .B(KEYINPUT10), .C1(new_n333), .C2(new_n334), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n279), .A2(new_n277), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n589), .B1(new_n229), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT10), .B1(new_n585), .B2(new_n269), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n591), .A2(new_n358), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n577), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n585), .A2(new_n269), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n214), .A2(new_n197), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n269), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n358), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT12), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n578), .A2(new_n363), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n600), .A2(new_n587), .A3(new_n342), .A4(new_n589), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n586), .B1(new_n596), .B2(new_n269), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT12), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n603), .A3(new_n358), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n599), .A2(new_n576), .A3(new_n601), .A4(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n594), .A2(KEYINPUT78), .A3(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n602), .A2(new_n603), .A3(new_n358), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n603), .B1(new_n602), .B2(new_n358), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT78), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n576), .A4(new_n601), .ZN(new_n611));
  INV_X1    g425(.A(G469), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n606), .A2(new_n611), .A3(new_n612), .A4(new_n187), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n187), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AND4_X1   g429(.A1(new_n577), .A2(new_n599), .A3(new_n601), .A4(new_n604), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n358), .B1(new_n591), .B2(new_n592), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n577), .B1(new_n617), .B2(new_n601), .ZN(new_n618));
  OAI21_X1  g432(.A(G469), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n613), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(G221), .B1(new_n556), .B2(G902), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n573), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n321), .A2(new_n471), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n558), .A2(new_n559), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n547), .A2(new_n554), .ZN(new_n628));
  INV_X1    g442(.A(new_n557), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n547), .A2(new_n554), .A3(new_n557), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT33), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(G478), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n560), .A2(G478), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n563), .A2(new_n187), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n520), .A2(new_n522), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n524), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n529), .B1(new_n642), .B2(new_n503), .ZN(new_n643));
  INV_X1    g457(.A(new_n530), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n638), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT93), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n308), .A2(new_n309), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n297), .A2(new_n305), .A3(new_n310), .A4(new_n307), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n316), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n571), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n390), .B1(new_n389), .B2(new_n187), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n391), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n620), .A2(new_n621), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n653), .A2(new_n469), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n646), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT34), .B(G104), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  NOR2_X1   g472(.A1(new_n639), .A2(new_n524), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n565), .B(new_n503), .C1(new_n659), .C2(new_n526), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n649), .A2(new_n571), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NOR2_X1   g478(.A1(new_n452), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n448), .B(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT94), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n666), .A2(new_n667), .A3(new_n467), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n666), .B2(new_n467), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n463), .A2(new_n465), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT95), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n463), .A2(KEYINPUT95), .A3(new_n465), .A4(new_n670), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n653), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n321), .A2(new_n623), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  INV_X1    g493(.A(new_n675), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n649), .A2(new_n654), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n567), .B1(new_n570), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n660), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n680), .A2(new_n681), .A3(new_n409), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XNOR2_X1  g500(.A(new_n683), .B(KEYINPUT39), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n654), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT97), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT40), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n680), .B1(new_n689), .B2(new_n690), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n315), .B(KEYINPUT38), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n354), .A2(new_n369), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n400), .B2(new_n387), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n695), .B2(G902), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n393), .A2(new_n408), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT96), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT96), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n393), .A2(new_n696), .A3(new_n699), .A4(new_n408), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n565), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n528), .B2(new_n530), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n701), .A2(new_n316), .A3(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n691), .A2(new_n692), .A3(new_n693), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n196), .ZN(G45));
  AOI211_X1 g520(.A(new_n683), .B(new_n637), .C1(new_n528), .C2(new_n530), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(new_n680), .A3(new_n681), .A4(new_n409), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  NAND3_X1  g523(.A1(new_n606), .A2(new_n187), .A3(new_n611), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n621), .A3(new_n613), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT98), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n711), .A2(KEYINPUT98), .A3(new_n621), .A4(new_n613), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n716), .A2(new_n409), .A3(new_n470), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n646), .A2(new_n650), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n661), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NOR3_X1   g536(.A1(new_n675), .A2(new_n649), .A3(new_n712), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(KEYINPUT99), .A3(new_n409), .A4(new_n573), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT99), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n647), .A2(new_n316), .A3(new_n648), .ZN(new_n726));
  INV_X1    g540(.A(new_n712), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n673), .A3(new_n674), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n573), .A2(new_n409), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  NAND2_X1  g546(.A1(new_n469), .A2(KEYINPUT100), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT100), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n463), .A2(new_n734), .A3(new_n465), .A4(new_n468), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT101), .B1(new_n736), .B2(new_n653), .ZN(new_n737));
  INV_X1    g551(.A(new_n391), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n651), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT101), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n733), .A4(new_n735), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n650), .A2(new_n716), .A3(new_n703), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  NOR2_X1   g559(.A1(new_n675), .A2(new_n649), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n739), .A3(new_n707), .A4(new_n727), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  INV_X1    g562(.A(new_n736), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n393), .A2(new_n750), .A3(new_n408), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n407), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n750), .B1(new_n393), .B2(new_n408), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n749), .B(KEYINPUT42), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n637), .B1(new_n528), .B2(new_n530), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n313), .A2(new_n316), .A3(new_n314), .ZN(new_n756));
  INV_X1    g570(.A(new_n683), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n755), .A2(new_n756), .A3(new_n622), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n622), .A2(new_n316), .A3(new_n313), .A4(new_n314), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n638), .B(new_n757), .C1(new_n643), .C2(new_n644), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT102), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n471), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n409), .A2(new_n470), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT102), .B1(new_n758), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n759), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n327), .ZN(G33));
  NAND4_X1  g584(.A1(new_n471), .A2(new_n622), .A3(new_n684), .A4(new_n756), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  INV_X1    g586(.A(KEYINPUT105), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n616), .A2(new_n618), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n612), .B1(new_n774), .B2(new_n775), .ZN(new_n777));
  OAI211_X1 g591(.A(KEYINPUT105), .B(KEYINPUT45), .C1(new_n616), .C2(new_n618), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n615), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT106), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n779), .A2(KEYINPUT106), .A3(KEYINPUT46), .A4(new_n615), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n613), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT107), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT46), .ZN(new_n787));
  INV_X1    g601(.A(new_n779), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n788), .B2(new_n614), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n782), .A2(KEYINPUT107), .A3(new_n613), .A4(new_n783), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n621), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n687), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT108), .Z(new_n794));
  NAND3_X1  g608(.A1(new_n638), .A2(new_n528), .A3(new_n530), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT43), .Z(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n653), .A3(new_n680), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  OR3_X1    g613(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n313), .A2(new_n316), .A3(new_n314), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n797), .B2(new_n799), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n798), .B1(new_n797), .B2(new_n799), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n794), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  INV_X1    g621(.A(KEYINPUT47), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(KEYINPUT110), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(KEYINPUT110), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n792), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n409), .A2(new_n470), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n761), .A2(new_n801), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n791), .A2(new_n621), .A3(new_n810), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  INV_X1    g633(.A(new_n567), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(new_n737), .B2(new_n741), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n693), .A2(new_n316), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n796), .A2(new_n821), .A3(new_n822), .A4(new_n727), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n819), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n801), .A2(new_n820), .A3(new_n712), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n470), .A2(new_n828), .A3(new_n698), .A4(new_n700), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n530), .A3(new_n528), .A4(new_n637), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n796), .A2(new_n676), .A3(new_n828), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT117), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n830), .A2(KEYINPUT117), .A3(new_n831), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n796), .A2(new_n821), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n756), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n711), .A2(new_n613), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n621), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n813), .B2(new_n816), .ZN(new_n838));
  OAI221_X1 g652(.A(new_n827), .B1(new_n832), .B2(new_n833), .C1(new_n835), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n796), .A2(new_n828), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT119), .Z(new_n843));
  NAND3_X1  g657(.A1(new_n834), .A2(new_n726), .A3(new_n727), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT118), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n844), .A2(KEYINPUT118), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n843), .A2(KEYINPUT48), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n566), .A2(G953), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n829), .A2(new_n646), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n839), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n816), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n791), .A2(new_n621), .B1(new_n811), .B2(new_n810), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT114), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n813), .A2(new_n854), .A3(new_n816), .ZN(new_n855));
  INV_X1    g669(.A(new_n837), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n835), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n830), .A2(new_n831), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n825), .A2(new_n826), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n825), .A2(KEYINPUT116), .A3(new_n826), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n857), .A2(KEYINPUT115), .A3(new_n858), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n850), .B1(new_n869), .B2(new_n819), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT113), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n321), .B(new_n623), .C1(new_n471), .C2(new_n676), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n528), .A2(new_n530), .A3(new_n565), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT111), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT111), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n528), .A2(new_n875), .A3(new_n530), .A4(new_n565), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n645), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n571), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n321), .A2(new_n877), .A3(new_n878), .A4(new_n655), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n659), .A2(new_n526), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(G475), .B2(new_n502), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n409), .A2(new_n702), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n755), .A2(new_n739), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n760), .A2(new_n683), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n680), .A3(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n872), .A2(new_n879), .A3(new_n886), .A4(new_n771), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n747), .A2(new_n685), .A3(new_n708), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n703), .A2(new_n726), .A3(new_n757), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n654), .A2(new_n671), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n701), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n888), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n681), .A2(new_n409), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n761), .A2(new_n675), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n675), .A2(new_n660), .A3(new_n683), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n701), .A2(new_n890), .A3(new_n891), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT52), .A4(new_n747), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n887), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n742), .A2(new_n743), .B1(new_n717), .B2(new_n661), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n731), .A3(new_n718), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n769), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n900), .A2(new_n903), .A3(KEYINPUT53), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT53), .B1(new_n900), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT54), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n901), .A2(new_n718), .A3(new_n731), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n763), .B1(new_n762), .B2(new_n471), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n758), .A2(new_n765), .A3(KEYINPUT102), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n768), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n759), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n907), .A2(new_n912), .A3(KEYINPUT112), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT112), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n769), .B2(new_n902), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n913), .A2(new_n915), .A3(KEYINPUT53), .A4(new_n900), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT53), .ZN(new_n917));
  AND4_X1   g731(.A1(new_n771), .A2(new_n872), .A3(new_n879), .A4(new_n886), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n747), .A2(new_n685), .A3(new_n708), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT52), .B1(new_n919), .B2(new_n898), .ZN(new_n920));
  AND4_X1   g734(.A1(KEYINPUT52), .A2(new_n897), .A3(new_n898), .A4(new_n747), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n907), .A2(new_n912), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n917), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n916), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n871), .B1(new_n906), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n906), .A2(new_n926), .A3(new_n871), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n870), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OR3_X1    g743(.A1(new_n842), .A2(KEYINPUT119), .A3(KEYINPUT48), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OAI22_X1  g745(.A1(new_n929), .A2(new_n931), .B1(G952), .B2(G953), .ZN(new_n932));
  INV_X1    g746(.A(new_n795), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n836), .B2(KEYINPUT49), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n693), .B(new_n934), .C1(KEYINPUT49), .C2(new_n836), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n698), .A2(new_n700), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n749), .A2(new_n621), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n935), .A2(new_n316), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n932), .A2(new_n938), .ZN(G75));
  AOI21_X1  g753(.A(new_n187), .B1(new_n916), .B2(new_n924), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT56), .B1(new_n940), .B2(G210), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n301), .A2(new_n302), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n303), .A2(new_n304), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n305), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT55), .Z(new_n946));
  XNOR2_X1  g760(.A(new_n941), .B(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n188), .A2(G952), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT120), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n949), .ZN(G51));
  INV_X1    g764(.A(KEYINPUT121), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n926), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n916), .A2(new_n924), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT54), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n916), .A2(new_n924), .A3(KEYINPUT121), .A4(new_n925), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n615), .A2(KEYINPUT57), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n615), .A2(KEYINPUT57), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n606), .A3(new_n611), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n940), .A2(new_n788), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n948), .B1(new_n960), .B2(new_n961), .ZN(G54));
  NAND3_X1  g776(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(new_n520), .Z(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(new_n948), .ZN(G60));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n627), .A2(new_n632), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n928), .A2(new_n927), .ZN(new_n968));
  XNOR2_X1  g782(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n636), .B(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n967), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n970), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n627), .A2(new_n632), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n956), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n949), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n966), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n949), .B1(new_n956), .B2(new_n973), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n928), .A2(new_n927), .A3(new_n972), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n978), .B(KEYINPUT123), .C1(new_n979), .C2(new_n967), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n977), .A2(new_n980), .ZN(G63));
  NAND2_X1  g795(.A1(G217), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT124), .Z(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT60), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n916), .B2(new_n924), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n949), .B1(new_n985), .B2(new_n666), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n466), .B2(new_n985), .ZN(new_n987));
  XNOR2_X1  g801(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G66));
  INV_X1    g803(.A(G224), .ZN(new_n990));
  OAI21_X1  g804(.A(G953), .B1(new_n569), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n907), .A2(new_n872), .A3(new_n879), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT126), .Z(new_n993));
  OAI21_X1  g807(.A(new_n991), .B1(new_n993), .B2(G953), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n942), .B1(G898), .B2(new_n188), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(G69));
  AOI21_X1  g810(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n705), .A2(new_n919), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(KEYINPUT62), .ZN(new_n1000));
  XOR2_X1   g814(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1001));
  NAND3_X1  g815(.A1(new_n705), .A2(new_n919), .A3(new_n1001), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n1000), .A2(new_n817), .A3(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n689), .A2(new_n471), .A3(new_n756), .A4(new_n877), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1003), .A2(new_n806), .A3(new_n1004), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n1005), .A2(new_n188), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n365), .A2(new_n368), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n506), .A2(new_n508), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1007), .B(new_n1008), .Z(new_n1009));
  NOR2_X1   g823(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n703), .A2(new_n726), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n804), .B1(new_n841), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n769), .B1(new_n794), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n919), .A2(new_n771), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1013), .A2(new_n188), .A3(new_n817), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(G900), .A2(G953), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1015), .A2(new_n1009), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n997), .B1(new_n1010), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n997), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1017), .B(new_n1020), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n1021), .ZN(G72));
  INV_X1    g836(.A(new_n948), .ZN(new_n1023));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT63), .Z(new_n1025));
  INV_X1    g839(.A(new_n403), .ZN(new_n1026));
  OAI221_X1 g840(.A(new_n1025), .B1(new_n1026), .B2(new_n694), .C1(new_n904), .C2(new_n905), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1025), .ZN(new_n1028));
  AND3_X1   g842(.A1(new_n1013), .A2(new_n817), .A3(new_n1014), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1028), .B1(new_n1029), .B2(new_n993), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n369), .A2(new_n379), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n387), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n1023), .B(new_n1027), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n993), .A2(new_n1003), .A3(new_n806), .A4(new_n1004), .ZN(new_n1034));
  AOI211_X1 g848(.A(new_n387), .B(new_n1031), .C1(new_n1034), .C2(new_n1025), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1033), .A2(new_n1035), .ZN(G57));
endmodule


