

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609;

  NOR2_X2 U326 ( .A1(n592), .A2(n555), .ZN(n471) );
  NOR2_X1 U327 ( .A1(n497), .A2(n496), .ZN(n509) );
  XNOR2_X1 U328 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n500) );
  XNOR2_X1 U329 ( .A(n458), .B(n457), .ZN(n461) );
  XOR2_X1 U330 ( .A(G204GAT), .B(G92GAT), .Z(n294) );
  XNOR2_X1 U331 ( .A(n448), .B(KEYINPUT47), .ZN(n449) );
  XNOR2_X1 U332 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U333 ( .A(n456), .B(KEYINPUT95), .ZN(n457) );
  INV_X1 U334 ( .A(KEYINPUT11), .ZN(n374) );
  XNOR2_X1 U335 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U336 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U337 ( .A(n462), .B(n294), .ZN(n463) );
  XNOR2_X1 U338 ( .A(n413), .B(n412), .ZN(n418) );
  XNOR2_X1 U339 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U340 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U341 ( .A(n501), .B(n500), .ZN(n543) );
  NOR2_X1 U342 ( .A1(n556), .A2(n479), .ZN(n588) );
  XOR2_X1 U343 ( .A(KEYINPUT115), .B(n471), .Z(n578) );
  INV_X1 U344 ( .A(G43GAT), .ZN(n504) );
  XNOR2_X1 U345 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U346 ( .A(n472), .B(G141GAT), .ZN(n473) );
  XNOR2_X1 U347 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U348 ( .A(n483), .B(n482), .ZN(G1349GAT) );
  XNOR2_X1 U349 ( .A(n507), .B(n506), .ZN(G1330GAT) );
  XOR2_X1 U350 ( .A(G78GAT), .B(G148GAT), .Z(n296) );
  XNOR2_X1 U351 ( .A(KEYINPUT76), .B(G204GAT), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n416) );
  INV_X1 U353 ( .A(KEYINPUT21), .ZN(n297) );
  NAND2_X1 U354 ( .A1(G211GAT), .A2(n297), .ZN(n300) );
  INV_X1 U355 ( .A(G211GAT), .ZN(n298) );
  NAND2_X1 U356 ( .A1(n298), .A2(KEYINPUT21), .ZN(n299) );
  NAND2_X1 U357 ( .A1(n300), .A2(n299), .ZN(n302) );
  XNOR2_X1 U358 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n455) );
  XNOR2_X1 U360 ( .A(n416), .B(n455), .ZN(n316) );
  XOR2_X1 U361 ( .A(KEYINPUT23), .B(KEYINPUT91), .Z(n304) );
  XNOR2_X1 U362 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U364 ( .A(G106GAT), .B(G218GAT), .Z(n306) );
  XOR2_X1 U365 ( .A(G50GAT), .B(G162GAT), .Z(n373) );
  XOR2_X1 U366 ( .A(G22GAT), .B(G155GAT), .Z(n379) );
  XNOR2_X1 U367 ( .A(n373), .B(n379), .ZN(n305) );
  XNOR2_X1 U368 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U369 ( .A(n308), .B(n307), .Z(n310) );
  NAND2_X1 U370 ( .A1(G228GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U371 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U372 ( .A(n311), .B(KEYINPUT89), .Z(n314) );
  XNOR2_X1 U373 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n312) );
  XNOR2_X1 U374 ( .A(n312), .B(KEYINPUT2), .ZN(n351) );
  XNOR2_X1 U375 ( .A(n351), .B(KEYINPUT90), .ZN(n313) );
  XNOR2_X1 U376 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n491) );
  XOR2_X1 U378 ( .A(G176GAT), .B(KEYINPUT86), .Z(n318) );
  XNOR2_X1 U379 ( .A(G113GAT), .B(KEYINPUT20), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n334) );
  XOR2_X1 U381 ( .A(G134GAT), .B(G99GAT), .Z(n320) );
  XNOR2_X1 U382 ( .A(G43GAT), .B(G190GAT), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U384 ( .A(n321), .B(KEYINPUT84), .Z(n323) );
  XOR2_X1 U385 ( .A(G120GAT), .B(G71GAT), .Z(n400) );
  XNOR2_X1 U386 ( .A(G169GAT), .B(n400), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U388 ( .A(KEYINPUT0), .B(KEYINPUT83), .Z(n344) );
  XOR2_X1 U389 ( .A(n344), .B(KEYINPUT85), .Z(n325) );
  NAND2_X1 U390 ( .A1(G227GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U391 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U392 ( .A(n327), .B(n326), .Z(n332) );
  XOR2_X1 U393 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n329) );
  XNOR2_X1 U394 ( .A(KEYINPUT87), .B(G183GAT), .ZN(n328) );
  XNOR2_X1 U395 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U396 ( .A(KEYINPUT18), .B(n330), .ZN(n465) );
  XOR2_X1 U397 ( .A(G15GAT), .B(G127GAT), .Z(n380) );
  XOR2_X1 U398 ( .A(n465), .B(n380), .Z(n331) );
  XNOR2_X1 U399 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n547) );
  INV_X1 U401 ( .A(n547), .ZN(n556) );
  NAND2_X1 U402 ( .A1(n491), .A2(n556), .ZN(n335) );
  XOR2_X1 U403 ( .A(n335), .B(KEYINPUT26), .Z(n484) );
  INV_X1 U404 ( .A(n484), .ZN(n592) );
  XOR2_X1 U405 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n337) );
  XNOR2_X1 U406 ( .A(G57GAT), .B(KEYINPUT6), .ZN(n336) );
  XNOR2_X1 U407 ( .A(n337), .B(n336), .ZN(n355) );
  XOR2_X1 U408 ( .A(G85GAT), .B(G155GAT), .Z(n339) );
  XNOR2_X1 U409 ( .A(G29GAT), .B(G162GAT), .ZN(n338) );
  XNOR2_X1 U410 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U411 ( .A(KEYINPUT92), .B(G148GAT), .Z(n341) );
  XNOR2_X1 U412 ( .A(G127GAT), .B(G120GAT), .ZN(n340) );
  XNOR2_X1 U413 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U414 ( .A(n343), .B(n342), .Z(n349) );
  XOR2_X1 U415 ( .A(G113GAT), .B(G1GAT), .Z(n430) );
  XOR2_X1 U416 ( .A(G134GAT), .B(KEYINPUT78), .Z(n365) );
  XOR2_X1 U417 ( .A(n365), .B(n344), .Z(n346) );
  NAND2_X1 U418 ( .A1(G225GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U419 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U420 ( .A(n430), .B(n347), .ZN(n348) );
  XNOR2_X1 U421 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U422 ( .A(n350), .B(KEYINPUT5), .Z(n353) );
  XNOR2_X1 U423 ( .A(n351), .B(KEYINPUT4), .ZN(n352) );
  XNOR2_X1 U424 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U425 ( .A(n355), .B(n354), .Z(n544) );
  INV_X1 U426 ( .A(n544), .ZN(n524) );
  XOR2_X1 U427 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n357) );
  XNOR2_X1 U428 ( .A(G43GAT), .B(G29GAT), .ZN(n356) );
  XNOR2_X1 U429 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U430 ( .A(KEYINPUT71), .B(n358), .ZN(n436) );
  INV_X1 U431 ( .A(G85GAT), .ZN(n359) );
  NAND2_X1 U432 ( .A1(n359), .A2(G92GAT), .ZN(n362) );
  INV_X1 U433 ( .A(G92GAT), .ZN(n360) );
  NAND2_X1 U434 ( .A1(n360), .A2(G85GAT), .ZN(n361) );
  NAND2_X1 U435 ( .A1(n362), .A2(n361), .ZN(n364) );
  XNOR2_X1 U436 ( .A(G99GAT), .B(G106GAT), .ZN(n363) );
  XNOR2_X1 U437 ( .A(n364), .B(n363), .ZN(n414) );
  XNOR2_X1 U438 ( .A(n414), .B(n365), .ZN(n367) );
  AND2_X1 U439 ( .A1(G232GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U440 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U441 ( .A(KEYINPUT9), .B(n368), .Z(n372) );
  XOR2_X1 U442 ( .A(KEYINPUT79), .B(G218GAT), .Z(n370) );
  XNOR2_X1 U443 ( .A(G36GAT), .B(G190GAT), .ZN(n369) );
  XNOR2_X1 U444 ( .A(n370), .B(n369), .ZN(n459) );
  XNOR2_X1 U445 ( .A(n459), .B(KEYINPUT10), .ZN(n371) );
  XNOR2_X1 U446 ( .A(n372), .B(n371), .ZN(n377) );
  XNOR2_X1 U447 ( .A(n373), .B(KEYINPUT65), .ZN(n375) );
  XOR2_X1 U448 ( .A(n436), .B(n378), .Z(n577) );
  XOR2_X1 U449 ( .A(KEYINPUT80), .B(n577), .Z(n567) );
  XNOR2_X1 U450 ( .A(n567), .B(KEYINPUT36), .ZN(n607) );
  XOR2_X1 U451 ( .A(n379), .B(G211GAT), .Z(n382) );
  XNOR2_X1 U452 ( .A(n380), .B(G78GAT), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n382), .B(n381), .ZN(n387) );
  XNOR2_X1 U454 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n383) );
  XNOR2_X1 U455 ( .A(n383), .B(KEYINPUT73), .ZN(n399) );
  XOR2_X1 U456 ( .A(n399), .B(KEYINPUT72), .Z(n385) );
  NAND2_X1 U457 ( .A1(G231GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U458 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U459 ( .A(n387), .B(n386), .Z(n389) );
  XNOR2_X1 U460 ( .A(G183GAT), .B(G71GAT), .ZN(n388) );
  XNOR2_X1 U461 ( .A(n389), .B(n388), .ZN(n397) );
  XOR2_X1 U462 ( .A(KEYINPUT14), .B(G64GAT), .Z(n391) );
  XNOR2_X1 U463 ( .A(G1GAT), .B(G8GAT), .ZN(n390) );
  XNOR2_X1 U464 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U465 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n393) );
  XNOR2_X1 U466 ( .A(KEYINPUT12), .B(KEYINPUT82), .ZN(n392) );
  XNOR2_X1 U467 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U468 ( .A(n395), .B(n394), .Z(n396) );
  XOR2_X1 U469 ( .A(n397), .B(n396), .Z(n584) );
  INV_X1 U470 ( .A(n584), .ZN(n604) );
  NOR2_X1 U471 ( .A1(n607), .A2(n604), .ZN(n398) );
  XNOR2_X1 U472 ( .A(n398), .B(KEYINPUT45), .ZN(n438) );
  NAND2_X1 U473 ( .A1(n399), .A2(n400), .ZN(n404) );
  INV_X1 U474 ( .A(n399), .ZN(n402) );
  INV_X1 U475 ( .A(n400), .ZN(n401) );
  NAND2_X1 U476 ( .A1(n402), .A2(n401), .ZN(n403) );
  NAND2_X1 U477 ( .A1(n404), .A2(n403), .ZN(n406) );
  AND2_X1 U478 ( .A1(G230GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U479 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U480 ( .A(KEYINPUT77), .B(n407), .Z(n413) );
  XOR2_X1 U481 ( .A(G176GAT), .B(G64GAT), .Z(n462) );
  XNOR2_X1 U482 ( .A(n462), .B(KEYINPUT74), .ZN(n411) );
  XOR2_X1 U483 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n409) );
  XNOR2_X1 U484 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n408) );
  XOR2_X1 U485 ( .A(n409), .B(n408), .Z(n410) );
  BUF_X1 U486 ( .A(n414), .Z(n415) );
  XNOR2_X1 U487 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U488 ( .A(n418), .B(n417), .ZN(n600) );
  XOR2_X1 U489 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n420) );
  XNOR2_X1 U490 ( .A(KEYINPUT70), .B(KEYINPUT30), .ZN(n419) );
  XNOR2_X1 U491 ( .A(n420), .B(n419), .ZN(n434) );
  XOR2_X1 U492 ( .A(G22GAT), .B(G141GAT), .Z(n422) );
  XNOR2_X1 U493 ( .A(G36GAT), .B(G50GAT), .ZN(n421) );
  XNOR2_X1 U494 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U495 ( .A(KEYINPUT29), .B(KEYINPUT72), .Z(n424) );
  XNOR2_X1 U496 ( .A(G197GAT), .B(G15GAT), .ZN(n423) );
  XNOR2_X1 U497 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U498 ( .A(n426), .B(n425), .Z(n432) );
  XOR2_X1 U499 ( .A(G169GAT), .B(G8GAT), .Z(n454) );
  XOR2_X1 U500 ( .A(n454), .B(KEYINPUT68), .Z(n428) );
  NAND2_X1 U501 ( .A1(G229GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U502 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U503 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U504 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U505 ( .A(n434), .B(n433), .Z(n435) );
  XOR2_X1 U506 ( .A(n436), .B(n435), .Z(n582) );
  INV_X1 U507 ( .A(n582), .ZN(n595) );
  AND2_X1 U508 ( .A1(n600), .A2(n595), .ZN(n437) );
  AND2_X1 U509 ( .A1(n438), .A2(n437), .ZN(n452) );
  XNOR2_X1 U510 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n441) );
  AND2_X1 U511 ( .A1(n582), .A2(n441), .ZN(n440) );
  XNOR2_X1 U512 ( .A(n600), .B(KEYINPUT64), .ZN(n439) );
  XNOR2_X1 U513 ( .A(KEYINPUT41), .B(n439), .ZN(n573) );
  NAND2_X1 U514 ( .A1(n440), .A2(n573), .ZN(n445) );
  NAND2_X1 U515 ( .A1(n582), .A2(n573), .ZN(n443) );
  INV_X1 U516 ( .A(n441), .ZN(n442) );
  NAND2_X1 U517 ( .A1(n443), .A2(n442), .ZN(n444) );
  NAND2_X1 U518 ( .A1(n445), .A2(n444), .ZN(n446) );
  NAND2_X1 U519 ( .A1(n446), .A2(n604), .ZN(n447) );
  NOR2_X1 U520 ( .A1(n577), .A2(n447), .ZN(n450) );
  INV_X1 U521 ( .A(KEYINPUT112), .ZN(n448) );
  NOR2_X1 U522 ( .A1(n452), .A2(n451), .ZN(n453) );
  XNOR2_X1 U523 ( .A(n453), .B(KEYINPUT48), .ZN(n475) );
  NOR2_X1 U524 ( .A1(n524), .A2(n475), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n455), .B(n454), .ZN(n458) );
  AND2_X1 U526 ( .A1(G226GAT), .A2(G233GAT), .ZN(n456) );
  XOR2_X1 U527 ( .A(n459), .B(KEYINPUT94), .Z(n460) );
  XNOR2_X1 U528 ( .A(n461), .B(n460), .ZN(n464) );
  XOR2_X1 U529 ( .A(n466), .B(n465), .Z(n467) );
  XNOR2_X1 U530 ( .A(n467), .B(KEYINPUT96), .ZN(n468) );
  XNOR2_X1 U531 ( .A(KEYINPUT27), .B(n468), .ZN(n493) );
  NAND2_X1 U532 ( .A1(n469), .A2(n493), .ZN(n470) );
  XOR2_X1 U533 ( .A(n470), .B(KEYINPUT113), .Z(n555) );
  NAND2_X1 U534 ( .A1(n578), .A2(n582), .ZN(n474) );
  XOR2_X1 U535 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n472) );
  XNOR2_X1 U536 ( .A(n474), .B(n473), .ZN(G1344GAT) );
  INV_X1 U537 ( .A(n467), .ZN(n527) );
  NOR2_X1 U538 ( .A1(n527), .A2(n475), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n476), .B(KEYINPUT54), .ZN(n477) );
  NAND2_X1 U540 ( .A1(n477), .A2(n524), .ZN(n591) );
  NOR2_X1 U541 ( .A1(n491), .A2(n591), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n478), .B(KEYINPUT55), .ZN(n479) );
  NAND2_X1 U543 ( .A1(n588), .A2(n573), .ZN(n483) );
  XOR2_X1 U544 ( .A(G176GAT), .B(KEYINPUT56), .Z(n481) );
  XNOR2_X1 U545 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n480) );
  INV_X1 U546 ( .A(KEYINPUT38), .ZN(n503) );
  NAND2_X1 U547 ( .A1(n484), .A2(n493), .ZN(n485) );
  NAND2_X1 U548 ( .A1(n524), .A2(n485), .ZN(n490) );
  NOR2_X1 U549 ( .A1(n556), .A2(n527), .ZN(n486) );
  NOR2_X1 U550 ( .A1(n491), .A2(n486), .ZN(n487) );
  XNOR2_X1 U551 ( .A(KEYINPUT25), .B(n487), .ZN(n488) );
  XNOR2_X1 U552 ( .A(KEYINPUT97), .B(n488), .ZN(n489) );
  NOR2_X1 U553 ( .A1(n490), .A2(n489), .ZN(n497) );
  XNOR2_X1 U554 ( .A(n491), .B(KEYINPUT66), .ZN(n492) );
  XOR2_X1 U555 ( .A(n492), .B(KEYINPUT28), .Z(n557) );
  INV_X1 U556 ( .A(n557), .ZN(n549) );
  NAND2_X1 U557 ( .A1(n556), .A2(n493), .ZN(n494) );
  NOR2_X1 U558 ( .A1(n549), .A2(n494), .ZN(n495) );
  NOR2_X1 U559 ( .A1(n495), .A2(n524), .ZN(n496) );
  NAND2_X1 U560 ( .A1(n509), .A2(n604), .ZN(n498) );
  XOR2_X1 U561 ( .A(KEYINPUT103), .B(n498), .Z(n499) );
  NOR2_X1 U562 ( .A1(n607), .A2(n499), .ZN(n501) );
  NAND2_X1 U563 ( .A1(n600), .A2(n582), .ZN(n511) );
  NOR2_X1 U564 ( .A1(n543), .A2(n511), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n530) );
  NOR2_X1 U566 ( .A1(n556), .A2(n530), .ZN(n507) );
  XNOR2_X1 U567 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n505) );
  INV_X1 U568 ( .A(n567), .ZN(n587) );
  NOR2_X1 U569 ( .A1(n587), .A2(n604), .ZN(n508) );
  XNOR2_X1 U570 ( .A(KEYINPUT16), .B(n508), .ZN(n510) );
  NAND2_X1 U571 ( .A1(n510), .A2(n509), .ZN(n534) );
  NOR2_X1 U572 ( .A1(n511), .A2(n534), .ZN(n521) );
  NAND2_X1 U573 ( .A1(n521), .A2(n544), .ZN(n512) );
  XNOR2_X1 U574 ( .A(n512), .B(KEYINPUT34), .ZN(n513) );
  XNOR2_X1 U575 ( .A(G1GAT), .B(n513), .ZN(G1324GAT) );
  NAND2_X1 U576 ( .A1(n467), .A2(n521), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(KEYINPUT98), .ZN(n515) );
  XNOR2_X1 U578 ( .A(G8GAT), .B(n515), .ZN(G1325GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n517) );
  XNOR2_X1 U580 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(n520) );
  NAND2_X1 U582 ( .A1(n547), .A2(n521), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n518), .B(KEYINPUT99), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1326GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n549), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n522), .B(KEYINPUT102), .ZN(n523) );
  XNOR2_X1 U587 ( .A(G22GAT), .B(n523), .ZN(G1327GAT) );
  NOR2_X1 U588 ( .A1(n530), .A2(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1328GAT) );
  XNOR2_X1 U591 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n529) );
  NOR2_X1 U592 ( .A1(n527), .A2(n530), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(G1329GAT) );
  NOR2_X1 U594 ( .A1(n530), .A2(n557), .ZN(n531) );
  XOR2_X1 U595 ( .A(G50GAT), .B(n531), .Z(G1331GAT) );
  XNOR2_X1 U596 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n532), .B(KEYINPUT108), .ZN(n533) );
  XOR2_X1 U598 ( .A(KEYINPUT107), .B(n533), .Z(n536) );
  NAND2_X1 U599 ( .A1(n595), .A2(n573), .ZN(n542) );
  NOR2_X1 U600 ( .A1(n542), .A2(n534), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n539), .A2(n544), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1332GAT) );
  NAND2_X1 U603 ( .A1(n467), .A2(n539), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U605 ( .A1(n547), .A2(n539), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n538), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U607 ( .A(G78GAT), .B(KEYINPUT43), .Z(n541) );
  NAND2_X1 U608 ( .A1(n539), .A2(n549), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(G1335GAT) );
  NOR2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n550), .A2(n544), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n545), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U613 ( .A1(n550), .A2(n467), .ZN(n546) );
  XNOR2_X1 U614 ( .A(G92GAT), .B(n546), .ZN(G1337GAT) );
  NAND2_X1 U615 ( .A1(n547), .A2(n550), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U617 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n554) );
  XOR2_X1 U618 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n552) );
  NAND2_X1 U619 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1339GAT) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n566) );
  NOR2_X1 U624 ( .A1(n595), .A2(n566), .ZN(n559) );
  XOR2_X1 U625 ( .A(G113GAT), .B(n559), .Z(G1340GAT) );
  INV_X1 U626 ( .A(n573), .ZN(n560) );
  NOR2_X1 U627 ( .A1(n560), .A2(n566), .ZN(n562) );
  XNOR2_X1 U628 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G120GAT), .B(n563), .ZN(G1341GAT) );
  NOR2_X1 U631 ( .A1(n604), .A2(n566), .ZN(n564) );
  XOR2_X1 U632 ( .A(KEYINPUT50), .B(n564), .Z(n565) );
  XNOR2_X1 U633 ( .A(G127GAT), .B(n565), .ZN(G1342GAT) );
  NOR2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1343GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n571) );
  XNOR2_X1 U638 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U640 ( .A(KEYINPUT118), .B(n572), .Z(n575) );
  NAND2_X1 U641 ( .A1(n578), .A2(n573), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(G1345GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n584), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n576), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n580) );
  XOR2_X1 U646 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n579) );
  XNOR2_X1 U647 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U649 ( .A1(n582), .A2(n588), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n583), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U651 ( .A(G183GAT), .B(KEYINPUT123), .Z(n586) );
  NAND2_X1 U652 ( .A1(n588), .A2(n584), .ZN(n585) );
  XNOR2_X1 U653 ( .A(n586), .B(n585), .ZN(G1350GAT) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n589), .B(KEYINPUT58), .ZN(n590) );
  XNOR2_X1 U656 ( .A(G190GAT), .B(n590), .ZN(G1351GAT) );
  INV_X1 U657 ( .A(KEYINPUT124), .ZN(n594) );
  NOR2_X1 U658 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n594), .B(n593), .ZN(n606) );
  NOR2_X1 U660 ( .A1(n606), .A2(n595), .ZN(n599) );
  XOR2_X1 U661 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n597) );
  XNOR2_X1 U662 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n596) );
  XNOR2_X1 U663 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X1 U664 ( .A(n599), .B(n598), .ZN(G1352GAT) );
  XNOR2_X1 U665 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n602) );
  NOR2_X1 U666 ( .A1(n600), .A2(n606), .ZN(n601) );
  XNOR2_X1 U667 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U668 ( .A(G204GAT), .B(n603), .ZN(G1353GAT) );
  NOR2_X1 U669 ( .A1(n606), .A2(n604), .ZN(n605) );
  XOR2_X1 U670 ( .A(n605), .B(G211GAT), .Z(G1354GAT) );
  NOR2_X1 U671 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U672 ( .A(KEYINPUT62), .B(n608), .Z(n609) );
  XNOR2_X1 U673 ( .A(G218GAT), .B(n609), .ZN(G1355GAT) );
endmodule

