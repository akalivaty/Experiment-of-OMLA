//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017, new_n1018;
  XOR2_X1   g000(.A(G57gat), .B(G85gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(G148gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G141gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT77), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(G141gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n218), .B1(G155gat), .B2(G162gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n213), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT78), .B(G141gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n214), .B1(new_n226), .B2(new_n211), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n223), .B1(new_n218), .B2(new_n224), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n221), .A2(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n231));
  INV_X1    g030(.A(G113gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G120gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n232), .A2(G120gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238));
  INV_X1    g037(.A(G127gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(G134gat), .ZN(new_n240));
  INV_X1    g039(.A(G134gat), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT67), .B1(new_n241), .B2(G127gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n239), .A2(G134gat), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n237), .B(new_n240), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(G134gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n241), .A2(G127gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT67), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n237), .B1(new_n248), .B2(new_n240), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n236), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n235), .B1(new_n251), .B2(new_n233), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n234), .A2(KEYINPUT69), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n246), .A2(new_n247), .A3(new_n231), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n230), .A2(new_n250), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n230), .B1(new_n250), .B2(new_n256), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n208), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n244), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n264), .A2(new_n236), .B1(new_n254), .B2(new_n255), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n230), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n265), .A2(KEYINPUT79), .A3(new_n266), .A4(new_n230), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n257), .A2(KEYINPUT4), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n273), .A2(new_n230), .B1(new_n250), .B2(new_n256), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n221), .A2(new_n225), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n229), .A2(new_n227), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n208), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n261), .B1(new_n272), .B2(new_n279), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n271), .A2(new_n267), .B1(new_n274), .B2(new_n278), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n282), .A3(new_n207), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n206), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n206), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n272), .A2(new_n279), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n286), .B(new_n283), .C1(new_n287), .C2(new_n261), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(KEYINPUT6), .B(new_n206), .C1(new_n280), .C2(new_n284), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT75), .ZN(new_n293));
  NAND2_X1  g092(.A1(G211gat), .A2(G218gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT22), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(G197gat), .A2(G204gat), .ZN(new_n297));
  AND2_X1   g096(.A1(G197gat), .A2(G204gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G211gat), .B(G218gat), .Z(new_n300));
  OAI21_X1  g099(.A(KEYINPUT74), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G197gat), .ZN(new_n302));
  INV_X1    g101(.A(G204gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G197gat), .A2(G204gat), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n304), .A2(new_n305), .B1(new_n295), .B2(new_n294), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n307));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n308), .B1(new_n306), .B2(KEYINPUT73), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n299), .A2(new_n311), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n301), .A2(new_n309), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(KEYINPUT23), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n315), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n321), .B1(KEYINPUT23), .B2(new_n314), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT64), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n320), .B(new_n322), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT24), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G183gat), .ZN(new_n329));
  INV_X1    g128(.A(G190gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(new_n319), .A3(new_n331), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n314), .A2(KEYINPUT23), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n322), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n323), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT25), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n325), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G226gat), .ZN(new_n338));
  INV_X1    g137(.A(G233gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n330), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n343), .A2(new_n345), .B1(G183gat), .B2(G190gat), .ZN(new_n346));
  OR2_X1    g145(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n348));
  AOI21_X1  g147(.A(G190gat), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OR2_X1    g148(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n344), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR3_X1   g153(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n346), .A2(new_n351), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n337), .A2(new_n340), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n326), .B1(new_n349), .B2(new_n344), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n350), .A2(new_n344), .ZN(new_n360));
  OAI22_X1  g159(.A1(new_n343), .A2(new_n360), .B1(new_n354), .B2(new_n355), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT66), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT66), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n346), .A2(new_n351), .A3(new_n363), .A4(new_n356), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n325), .A2(new_n336), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n340), .A2(KEYINPUT29), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n313), .B(new_n358), .C1(new_n367), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n362), .A2(new_n364), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n337), .A2(new_n371), .A3(new_n340), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n325), .A2(new_n357), .A3(new_n336), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n368), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT74), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n300), .B1(new_n299), .B2(new_n311), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n306), .A2(KEYINPUT73), .ZN(new_n379));
  OAI22_X1  g178(.A1(new_n376), .A2(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n293), .B1(new_n370), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n369), .B1(new_n337), .B2(new_n371), .ZN(new_n383));
  INV_X1    g182(.A(new_n340), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n373), .A2(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n383), .A2(new_n385), .A3(new_n380), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(KEYINPUT75), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT37), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(G64gat), .B(G92gat), .Z(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT76), .ZN(new_n390));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  AOI21_X1  g191(.A(new_n313), .B1(new_n372), .B2(new_n374), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT75), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT37), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n370), .A2(new_n293), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n388), .A2(KEYINPUT38), .A3(new_n392), .A4(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n395), .B1(new_n375), .B2(new_n313), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n358), .B1(new_n367), .B2(new_n369), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n399), .B1(new_n313), .B2(new_n400), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n397), .A2(new_n392), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n398), .B1(new_n402), .B2(KEYINPUT38), .ZN(new_n403));
  INV_X1    g202(.A(new_n392), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n394), .A2(new_n404), .A3(new_n396), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n292), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n392), .B1(new_n382), .B2(new_n387), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT30), .A3(new_n405), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n394), .A2(new_n409), .A3(new_n396), .A4(new_n404), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT86), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n274), .A2(new_n278), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n257), .A2(KEYINPUT4), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n266), .B1(new_n265), .B2(new_n230), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n418), .B2(new_n208), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n281), .A2(KEYINPUT86), .A3(new_n207), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n413), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n414), .A3(new_n208), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT86), .B1(new_n281), .B2(new_n207), .ZN(new_n423));
  OR3_X1    g222(.A1(new_n258), .A2(new_n259), .A3(new_n208), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT39), .A4(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n421), .A2(new_n425), .A3(KEYINPUT40), .A4(new_n286), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n426), .A2(new_n285), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n421), .A2(new_n286), .A3(new_n425), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT40), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G78gat), .B(G106gat), .Z(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(G22gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT81), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G228gat), .A2(G233gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n380), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n230), .B1(new_n439), .B2(new_n273), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n230), .A2(new_n273), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n380), .B1(new_n441), .B2(new_n438), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n437), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT29), .B1(new_n230), .B2(new_n273), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n380), .ZN(new_n446));
  INV_X1    g245(.A(new_n225), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n214), .A2(new_n215), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n219), .B1(new_n448), .B2(KEYINPUT77), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n449), .B2(new_n217), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n209), .A2(KEYINPUT78), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n209), .A2(KEYINPUT78), .ZN(new_n452));
  OAI21_X1  g251(.A(G148gat), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n228), .B1(new_n453), .B2(new_n214), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n450), .A2(new_n454), .A3(KEYINPUT3), .ZN(new_n455));
  OAI211_X1 g254(.A(KEYINPUT83), .B(new_n313), .C1(new_n455), .C2(KEYINPUT29), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n446), .A2(new_n436), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n301), .A2(new_n309), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n299), .A2(new_n300), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT29), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT3), .B1(new_n460), .B2(KEYINPUT82), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n301), .A2(new_n309), .B1(new_n300), .B2(new_n299), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(KEYINPUT29), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n230), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n443), .B1(new_n457), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT84), .B(G50gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT31), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n443), .B(new_n467), .C1(new_n457), .C2(new_n465), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n469), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n435), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(KEYINPUT82), .A3(new_n438), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(new_n464), .A3(new_n273), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n277), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n478), .A2(new_n436), .A3(new_n456), .A4(new_n446), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n467), .B1(new_n479), .B2(new_n443), .ZN(new_n480));
  INV_X1    g279(.A(new_n471), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT31), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n434), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n474), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n406), .A2(new_n431), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n472), .A2(new_n473), .A3(new_n435), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n434), .B1(new_n482), .B2(new_n483), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n290), .A2(new_n291), .B1(new_n408), .B2(new_n410), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n474), .A2(KEYINPUT85), .A3(new_n484), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n337), .A2(new_n265), .A3(new_n371), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n265), .B1(new_n337), .B2(new_n371), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G227gat), .A2(G233gat), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n497), .A2(KEYINPUT72), .A3(KEYINPUT34), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n250), .A2(new_n256), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n365), .B2(new_n366), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n337), .A2(new_n371), .A3(new_n265), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n498), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT71), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT32), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n503), .B2(new_n504), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G43gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(G71gat), .B(G99gat), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n511), .B(new_n512), .Z(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT33), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n508), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n504), .B1(new_n495), .B2(new_n496), .ZN(new_n516));
  AND4_X1   g315(.A1(new_n508), .A2(new_n516), .A3(KEYINPUT32), .A4(new_n514), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT70), .B1(new_n519), .B2(new_n509), .ZN(new_n520));
  INV_X1    g319(.A(new_n513), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT33), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n521), .B1(new_n516), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n524), .A3(KEYINPUT32), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n520), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n507), .B1(new_n518), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n516), .A2(KEYINPUT32), .A3(new_n514), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT71), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n508), .A3(new_n514), .ZN(new_n530));
  AND4_X1   g329(.A1(new_n526), .A2(new_n529), .A3(new_n530), .A4(new_n507), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT36), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT36), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n527), .B2(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n486), .A2(new_n494), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n485), .A2(new_n532), .A3(new_n491), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT35), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n485), .A2(new_n532), .A3(new_n491), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT16), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n545), .B2(G1gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(G1gat), .B2(new_n544), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G8gat), .ZN(new_n548));
  XOR2_X1   g347(.A(G71gat), .B(G78gat), .Z(new_n549));
  AOI21_X1  g348(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n549), .B1(new_n552), .B2(KEYINPUT92), .ZN(new_n553));
  XOR2_X1   g352(.A(G57gat), .B(G64gat), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n552), .B(new_n554), .C1(KEYINPUT92), .C2(new_n549), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n548), .B1(new_n558), .B2(KEYINPUT21), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n558), .B(KEYINPUT21), .Z(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(new_n548), .ZN(new_n561));
  XNOR2_X1  g360(.A(G127gat), .B(G155gat), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n561), .B(new_n562), .Z(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n561), .B(new_n562), .ZN(new_n566));
  INV_X1    g365(.A(new_n564), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(new_n329), .ZN(new_n571));
  INV_X1    g370(.A(G211gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n565), .A2(new_n568), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(new_n302), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT11), .B(G169gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT12), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G43gat), .B(G50gat), .Z(new_n586));
  INV_X1    g385(.A(KEYINPUT15), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT14), .ZN(new_n588));
  INV_X1    g387(.A(G29gat), .ZN(new_n589));
  INV_X1    g388(.A(G36gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n586), .A2(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G29gat), .A2(G36gat), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n593), .B(new_n594), .C1(new_n587), .C2(new_n586), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n591), .A2(KEYINPUT88), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n592), .B1(new_n591), .B2(KEYINPUT88), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n586), .A2(new_n587), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT17), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT89), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT89), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n595), .A2(new_n600), .A3(new_n604), .A4(KEYINPUT17), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n548), .B1(new_n602), .B2(new_n601), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n606), .A2(new_n607), .B1(new_n601), .B2(new_n548), .ZN(new_n608));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT90), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT18), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n548), .B(new_n601), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n609), .B(KEYINPUT13), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n610), .B2(new_n611), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n585), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n610), .A2(new_n611), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n619), .A2(new_n612), .A3(new_n616), .A4(new_n584), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n622));
  INV_X1    g421(.A(G230gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n623), .A2(new_n339), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT98), .B(G92gat), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT8), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(G99gat), .B2(G106gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n634));
  AOI21_X1  g433(.A(G85gat), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT99), .B1(new_n635), .B2(new_n630), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G99gat), .B(G106gat), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT7), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n640), .B2(KEYINPUT96), .ZN(new_n641));
  NAND2_X1  g440(.A1(G85gat), .A2(G92gat), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(G92gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n641), .B1(new_n626), .B2(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n643), .B(new_n645), .C1(new_n639), .C2(new_n640), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n637), .A2(new_n638), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n638), .B1(new_n637), .B2(new_n646), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n557), .B(new_n556), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n637), .A2(new_n646), .ZN(new_n651));
  INV_X1    g450(.A(new_n638), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n638), .A3(new_n646), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n558), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n649), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n647), .A2(new_n648), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(KEYINPUT10), .A3(new_n558), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n624), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n649), .A2(new_n655), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n660), .A2(new_n624), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n622), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR4_X1   g467(.A1(new_n659), .A2(new_n661), .A3(KEYINPUT100), .A4(new_n665), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n662), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n668), .A2(new_n670), .B1(new_n671), .B2(new_n665), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n621), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n657), .B1(new_n602), .B2(new_n601), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n606), .ZN(new_n675));
  NAND2_X1  g474(.A1(G232gat), .A2(G233gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT95), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AOI22_X1  g477(.A1(new_n657), .A2(new_n601), .B1(KEYINPUT41), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G134gat), .B(G162gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n678), .A2(KEYINPUT41), .ZN(new_n683));
  XNOR2_X1  g482(.A(G190gat), .B(G218gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n682), .B(new_n685), .Z(new_n686));
  NOR3_X1   g485(.A1(new_n579), .A2(new_n673), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n543), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n292), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g490(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n692));
  OR2_X1    g491(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n689), .A2(new_n412), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(KEYINPUT42), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n689), .A2(new_n412), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(G8gat), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n695), .B1(new_n694), .B2(new_n698), .ZN(G1325gat));
  INV_X1    g498(.A(G15gat), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n688), .A2(new_n700), .A3(new_n536), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n689), .A2(new_n532), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n700), .B2(new_n702), .ZN(G1326gat));
  NAND2_X1  g502(.A1(new_n490), .A2(new_n493), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT43), .B(G22gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  INV_X1    g506(.A(new_n579), .ZN(new_n708));
  INV_X1    g507(.A(new_n672), .ZN(new_n709));
  INV_X1    g508(.A(new_n621), .ZN(new_n710));
  INV_X1    g509(.A(new_n686), .ZN(new_n711));
  NOR4_X1   g510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n712), .A2(new_n543), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n589), .A3(new_n292), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT45), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n543), .B2(new_n686), .ZN(new_n717));
  AOI211_X1 g516(.A(KEYINPUT44), .B(new_n711), .C1(new_n537), .C2(new_n542), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n578), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT101), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n575), .B1(new_n565), .B2(new_n568), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT101), .B1(new_n577), .B2(new_n578), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n673), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n719), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n292), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n715), .B1(new_n731), .B2(new_n589), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT102), .Z(G1328gat));
  NAND3_X1  g532(.A1(new_n713), .A2(new_n590), .A3(new_n412), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT46), .Z(new_n735));
  NAND2_X1  g534(.A1(new_n729), .A2(new_n412), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n737), .B2(new_n590), .ZN(G1329gat));
  INV_X1    g537(.A(new_n536), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n729), .A2(G43gat), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n713), .ZN(new_n741));
  INV_X1    g540(.A(new_n532), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n740), .B1(G43gat), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g544(.A(G50gat), .ZN(new_n746));
  INV_X1    g545(.A(new_n704), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n713), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n543), .A2(new_n686), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT44), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n711), .B1(new_n537), .B2(new_n542), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n716), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(new_n747), .A3(new_n727), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n750), .B1(new_n756), .B2(G50gat), .ZN(new_n757));
  INV_X1    g556(.A(new_n485), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n758), .A3(new_n727), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G50gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n748), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n757), .B1(new_n761), .B2(KEYINPUT48), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT103), .ZN(G1331gat));
  NOR2_X1   g562(.A1(new_n686), .A2(new_n579), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(new_n709), .A3(new_n710), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT104), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n543), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n292), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g569(.A(new_n411), .B(new_n767), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n771));
  NOR2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1333gat));
  NAND3_X1  g572(.A1(new_n768), .A2(G71gat), .A3(new_n739), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n767), .A2(new_n742), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(G71gat), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g576(.A1(new_n768), .A2(new_n747), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g578(.A1(new_n708), .A2(new_n621), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n753), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT51), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n672), .ZN(new_n783));
  AOI21_X1  g582(.A(G85gat), .B1(new_n783), .B2(new_n292), .ZN(new_n784));
  INV_X1    g583(.A(new_n780), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(new_n672), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n717), .B2(new_n718), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT105), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT105), .B(new_n786), .C1(new_n717), .C2(new_n718), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n290), .A2(new_n291), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n626), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n784), .B1(new_n791), .B2(new_n793), .ZN(G1336gat));
  AOI21_X1  g593(.A(KEYINPUT105), .B1(new_n755), .B2(new_n786), .ZN(new_n795));
  INV_X1    g594(.A(new_n790), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n412), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n625), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(KEYINPUT106), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT106), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n411), .B1(new_n789), .B2(new_n790), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(new_n625), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n781), .A2(KEYINPUT107), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n782), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n781), .A2(KEYINPUT107), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n411), .A2(G92gat), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n804), .A2(new_n709), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n799), .A2(new_n802), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT52), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(new_n783), .B2(new_n807), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n755), .A2(new_n412), .A3(new_n786), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(new_n625), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n814), .ZN(G1337gat));
  INV_X1    g614(.A(G99gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n783), .A2(new_n816), .A3(new_n532), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n536), .B1(new_n789), .B2(new_n790), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n816), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT108), .ZN(G1338gat));
  NOR3_X1   g619(.A1(new_n485), .A2(new_n672), .A3(G106gat), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n804), .A2(new_n806), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(G106gat), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n791), .B2(new_n747), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT53), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G106gat), .B1(new_n787), .B2(new_n485), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  INV_X1    g626(.A(new_n821), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n826), .B(new_n827), .C1(new_n782), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n829), .ZN(G1339gat));
  NAND3_X1  g629(.A1(new_n656), .A2(new_n658), .A3(new_n624), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n659), .B2(KEYINPUT109), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT109), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n656), .A2(new_n833), .A3(new_n658), .A4(new_n624), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(KEYINPUT54), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n666), .B1(new_n659), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(KEYINPUT55), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT110), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n835), .A2(new_n840), .A3(KEYINPUT55), .A4(new_n837), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n667), .A2(new_n669), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT55), .B1(new_n835), .B2(new_n837), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n842), .A2(new_n844), .A3(new_n621), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n608), .A2(new_n609), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n614), .A2(new_n615), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n583), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n620), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n672), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n686), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n843), .B1(new_n839), .B2(new_n841), .ZN(new_n855));
  INV_X1    g654(.A(new_n851), .ZN(new_n856));
  AND4_X1   g655(.A1(new_n686), .A2(new_n855), .A3(new_n846), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n725), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NOR4_X1   g657(.A1(new_n579), .A2(new_n686), .A3(new_n709), .A4(new_n621), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n792), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n758), .A2(new_n742), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n411), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT111), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n232), .A3(new_n621), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n843), .B(new_n845), .C1(new_n839), .C2(new_n841), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n686), .A3(new_n856), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n852), .B1(new_n867), .B2(new_n621), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(new_n686), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n859), .B1(new_n870), .B2(new_n725), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n292), .A2(new_n411), .ZN(new_n872));
  OR4_X1    g671(.A1(new_n747), .A2(new_n871), .A3(new_n742), .A4(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G113gat), .B1(new_n873), .B2(new_n710), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n866), .A2(new_n874), .ZN(G1340gat));
  INV_X1    g674(.A(G120gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n865), .A2(new_n876), .A3(new_n709), .ZN(new_n877));
  OAI21_X1  g676(.A(G120gat), .B1(new_n873), .B2(new_n672), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(G1341gat));
  NOR3_X1   g681(.A1(new_n873), .A2(new_n239), .A3(new_n725), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n863), .A2(new_n411), .A3(new_n708), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n884), .A2(KEYINPUT113), .ZN(new_n885));
  AOI21_X1  g684(.A(G127gat), .B1(new_n884), .B2(KEYINPUT113), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(G1342gat));
  NAND4_X1  g686(.A1(new_n863), .A2(new_n241), .A3(new_n411), .A4(new_n686), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n889));
  OAI21_X1  g688(.A(G134gat), .B1(new_n873), .B2(new_n711), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT114), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n889), .A2(KEYINPUT114), .A3(new_n890), .A4(new_n891), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1343gat));
  INV_X1    g695(.A(new_n226), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n835), .A2(new_n837), .ZN(new_n898));
  XNOR2_X1  g697(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n618), .A2(new_n620), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n852), .B1(new_n855), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n868), .B1(new_n901), .B2(new_n686), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n859), .B1(new_n902), .B2(new_n579), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT57), .B1(new_n903), .B2(new_n704), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n858), .A2(new_n860), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT57), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n906), .A3(new_n758), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n739), .A2(new_n872), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT115), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n904), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT117), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n904), .A2(new_n907), .A3(new_n912), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n897), .B1(new_n914), .B2(new_n621), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n536), .A2(KEYINPUT118), .A3(new_n758), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT118), .B1(new_n536), .B2(new_n758), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n710), .A2(G141gat), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n861), .A2(new_n411), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT58), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n904), .A2(new_n907), .A3(new_n621), .A4(new_n909), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT58), .B1(new_n924), .B2(new_n226), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n905), .A2(new_n292), .A3(new_n919), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n926), .A2(KEYINPUT119), .A3(new_n411), .A4(new_n920), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT120), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n925), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n923), .A2(new_n935), .ZN(G1344gat));
  AND2_X1   g735(.A1(new_n926), .A2(new_n411), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n211), .A3(new_n709), .ZN(new_n938));
  AOI211_X1 g737(.A(KEYINPUT59), .B(new_n211), .C1(new_n914), .C2(new_n709), .ZN(new_n939));
  XOR2_X1   g738(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n940));
  OAI21_X1  g739(.A(KEYINPUT57), .B1(new_n871), .B2(new_n485), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n855), .A2(new_n900), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n686), .B1(new_n942), .B2(new_n853), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n579), .B1(new_n943), .B2(new_n857), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n860), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n906), .A3(new_n747), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n941), .A2(new_n709), .A3(new_n909), .A4(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n940), .B1(new_n947), .B2(G148gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n938), .B1(new_n939), .B2(new_n948), .ZN(G1345gat));
  AOI21_X1  g748(.A(G155gat), .B1(new_n937), .B2(new_n708), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n726), .A2(G155gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n914), .B2(new_n951), .ZN(G1346gat));
  NOR3_X1   g751(.A1(new_n711), .A2(G162gat), .A3(new_n412), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n926), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n914), .A2(new_n955), .A3(new_n686), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G162gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n955), .B1(new_n914), .B2(new_n686), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1347gat));
  NOR2_X1   g758(.A1(new_n871), .A2(new_n292), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(new_n412), .A3(new_n862), .ZN(new_n961));
  INV_X1    g760(.A(G169gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(new_n962), .A3(new_n621), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n412), .A2(new_n792), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n742), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT123), .Z(new_n966));
  NAND3_X1  g765(.A1(new_n905), .A2(new_n704), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n905), .A2(new_n969), .A3(new_n704), .A4(new_n966), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(new_n621), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n963), .B1(new_n972), .B2(new_n962), .ZN(G1348gat));
  AOI21_X1  g772(.A(G176gat), .B1(new_n961), .B2(new_n709), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n709), .A2(G176gat), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n974), .B1(new_n971), .B2(new_n975), .ZN(G1349gat));
  AOI21_X1  g775(.A(new_n329), .B1(new_n971), .B2(new_n726), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n579), .B1(new_n347), .B2(new_n348), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n961), .A2(new_n978), .ZN(new_n979));
  OR3_X1    g778(.A1(new_n977), .A2(new_n979), .A3(KEYINPUT60), .ZN(new_n980));
  OAI21_X1  g779(.A(KEYINPUT60), .B1(new_n977), .B2(new_n979), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1350gat));
  NAND3_X1  g781(.A1(new_n968), .A2(new_n686), .A3(new_n970), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n983), .A2(new_n984), .A3(G190gat), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT126), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n983), .A2(KEYINPUT126), .A3(new_n984), .A4(G190gat), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n983), .A2(G190gat), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n987), .B(new_n988), .C1(new_n984), .C2(new_n989), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n961), .A2(new_n330), .A3(new_n686), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT125), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1351gat));
  AND4_X1   g792(.A1(new_n758), .A2(new_n960), .A3(new_n412), .A4(new_n536), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n994), .A2(new_n302), .A3(new_n621), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n739), .A2(new_n964), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n941), .A2(new_n946), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g796(.A(G197gat), .B1(new_n997), .B2(new_n710), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n995), .A2(new_n998), .ZN(G1352gat));
  NAND3_X1  g798(.A1(new_n994), .A2(new_n303), .A3(new_n709), .ZN(new_n1000));
  OR2_X1    g799(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n941), .A2(new_n709), .A3(new_n946), .ZN(new_n1002));
  INV_X1    g801(.A(new_n996), .ZN(new_n1003));
  OAI21_X1  g802(.A(G204gat), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1001), .A2(new_n1004), .A3(new_n1005), .ZN(G1353gat));
  NAND3_X1  g805(.A1(new_n994), .A2(new_n572), .A3(new_n708), .ZN(new_n1007));
  NAND4_X1  g806(.A1(new_n941), .A2(new_n708), .A3(new_n946), .A4(new_n996), .ZN(new_n1008));
  AND3_X1   g807(.A1(new_n1008), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1009));
  AOI21_X1  g808(.A(KEYINPUT63), .B1(new_n1008), .B2(G211gat), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT127), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g812(.A(KEYINPUT127), .B(new_n1007), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(G1354gat));
  AOI21_X1  g814(.A(G218gat), .B1(new_n994), .B2(new_n686), .ZN(new_n1016));
  INV_X1    g815(.A(new_n997), .ZN(new_n1017));
  AND2_X1   g816(.A1(new_n686), .A2(G218gat), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(G1355gat));
endmodule


