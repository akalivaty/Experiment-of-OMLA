//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n556, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(G319));
  OR2_X1    g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n464), .A2(KEYINPUT67), .A3(G101), .A4(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n463), .A2(G137), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n470), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n469), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  AOI21_X1  g048(.A(new_n464), .B1(new_n461), .B2(new_n462), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT68), .Z(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n479), .B1(G136), .B2(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(new_n474), .A2(G126), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT70), .B1(new_n464), .B2(G114), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(new_n489), .A3(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n486), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AOI211_X1 g069(.A(KEYINPUT71), .B(new_n492), .C1(new_n487), .C2(new_n490), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n485), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n498), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n470), .B2(new_n498), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n496), .A2(new_n505), .ZN(G164));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT72), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n507), .A2(new_n508), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT5), .B(G543), .Z(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n520), .A2(new_n513), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n522), .A2(G651), .B1(new_n523), .B2(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n518), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n510), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n509), .A2(G89), .ZN(new_n531));
  NAND2_X1  g106(.A1(G63), .A2(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n520), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G168));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT5), .B(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n509), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n535), .A2(new_n510), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n536), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G651), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n539), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n520), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n523), .A2(G81), .B1(new_n515), .B2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g130(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n556));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n515), .A2(G53), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT9), .Z(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT75), .B(G65), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n536), .A2(new_n562), .B1(G78), .B2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G91), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n563), .A2(new_n541), .B1(new_n537), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  OR2_X1    g143(.A1(new_n536), .A2(G74), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(new_n515), .B2(G49), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n523), .A2(G87), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n523), .A2(G86), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n515), .A2(G48), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n536), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n541), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT76), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n573), .A2(new_n574), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  NOR3_X1   g156(.A1(new_n580), .A2(new_n581), .A3(new_n577), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n579), .A2(new_n582), .ZN(G305));
  INV_X1    g158(.A(G47), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n584), .A2(new_n510), .B1(new_n537), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n541), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n523), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT10), .Z(new_n593));
  NAND2_X1  g168(.A1(new_n536), .A2(G66), .ZN(new_n594));
  INV_X1    g169(.A(G79), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT77), .B1(new_n595), .B2(new_n514), .ZN(new_n596));
  OR3_X1    g171(.A1(new_n595), .A2(new_n514), .A3(KEYINPUT77), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n515), .B2(G54), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n566), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(new_n566), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n601), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n601), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(KEYINPUT78), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(KEYINPUT78), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n611), .B(new_n612), .C1(G868), .C2(new_n553), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g189(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n463), .A2(G135), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n474), .A2(G123), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n464), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT79), .B(G2096), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n618), .A2(new_n625), .ZN(G156));
  INV_X1    g201(.A(G14), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n627), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n641), .A2(KEYINPUT80), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT80), .ZN(new_n643));
  NOR3_X1   g218(.A1(new_n638), .A2(new_n643), .A3(new_n639), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n640), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n650), .B2(KEYINPUT18), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT81), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT18), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(KEYINPUT17), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n648), .A2(new_n649), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n653), .B(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n660));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n664), .A2(new_n665), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  MUX2_X1   g246(.A(new_n671), .B(new_n670), .S(new_n663), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT84), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(KEYINPUT83), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n660), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n679), .A3(new_n660), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n684), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n682), .B1(new_n686), .B2(new_n680), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n685), .A2(new_n687), .A3(new_n689), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G19), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n553), .B2(new_n694), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(G1341), .Z(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G27), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G164), .B2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G2078), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n694), .A2(G21), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G168), .B2(new_n694), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1966), .ZN(new_n705));
  AND2_X1   g280(.A1(KEYINPUT24), .A2(G34), .ZN(new_n706));
  NOR2_X1   g281(.A1(KEYINPUT24), .A2(G34), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n698), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT87), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G160), .B2(G29), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G2084), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n705), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G32), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n474), .A2(G129), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(KEYINPUT26), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(KEYINPUT26), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT88), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n463), .A2(G141), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(new_n713), .B(new_n723), .S(G29), .Z(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT89), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n697), .A2(new_n702), .A3(new_n712), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n698), .A2(G33), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(new_n464), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT25), .ZN(new_n732));
  NAND2_X1  g307(.A1(G103), .A2(G2104), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G2105), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n463), .A2(G139), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n729), .B1(new_n738), .B2(new_n698), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2072), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n694), .A2(G5), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G301), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1961), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n724), .B2(new_n725), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT31), .B(G11), .Z(new_n746));
  INV_X1    g321(.A(G28), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT90), .Z(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n747), .B2(KEYINPUT30), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n751), .B1(new_n698), .B2(new_n623), .C1(new_n742), .C2(new_n743), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n463), .A2(G140), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n474), .A2(G128), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n464), .A2(G116), .ZN(new_n755));
  OAI21_X1  g330(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n753), .B(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G29), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n698), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2067), .ZN(new_n762));
  OR4_X1    g337(.A1(new_n740), .A2(new_n745), .A3(new_n752), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n694), .A2(G4), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n601), .B2(new_n694), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1348), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n694), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(G1956), .Z(new_n770));
  NOR4_X1   g345(.A1(new_n728), .A2(new_n763), .A3(new_n766), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n483), .A2(G29), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n698), .A2(G35), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT91), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(KEYINPUT29), .ZN(new_n776));
  INV_X1    g351(.A(G2090), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n772), .A2(new_n778), .A3(new_n774), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT92), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n776), .A2(new_n779), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G2090), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n771), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT34), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT86), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n694), .B1(new_n570), .B2(new_n571), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n694), .A2(G23), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(KEYINPUT33), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n787), .A2(KEYINPUT33), .A3(new_n789), .ZN(new_n792));
  OAI21_X1  g367(.A(G1976), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n792), .ZN(new_n794));
  INV_X1    g369(.A(G1976), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n794), .A2(new_n790), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(G16), .A2(G22), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G303), .B2(new_n694), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1971), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT32), .B(G1981), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT85), .ZN(new_n803));
  NOR2_X1   g378(.A1(G6), .A2(G16), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n803), .B(new_n805), .C1(G305), .C2(new_n694), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n575), .A2(KEYINPUT76), .A3(new_n578), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n581), .B1(new_n580), .B2(new_n577), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n694), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT85), .B1(new_n809), .B2(new_n804), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n802), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n801), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n806), .A2(new_n802), .A3(new_n810), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n786), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n811), .ZN(new_n815));
  INV_X1    g390(.A(G1971), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n799), .B(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n793), .B2(new_n796), .ZN(new_n818));
  AND4_X1   g393(.A1(new_n786), .A2(new_n815), .A3(new_n818), .A4(new_n813), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n785), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n815), .A2(new_n818), .A3(new_n813), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT86), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n812), .A2(new_n786), .A3(new_n813), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT34), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n694), .A2(G24), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n589), .B2(new_n694), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1986), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n698), .A2(G25), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n474), .A2(G119), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n463), .A2(G131), .ZN(new_n830));
  OR2_X1    g405(.A1(G95), .A2(G2105), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n831), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n828), .B1(new_n834), .B2(new_n698), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT35), .B(G1991), .Z(new_n836));
  XOR2_X1   g411(.A(new_n835), .B(new_n836), .Z(new_n837));
  NOR2_X1   g412(.A1(new_n827), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n820), .A2(new_n824), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n820), .A2(new_n841), .A3(new_n824), .A4(new_n838), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n784), .B1(new_n840), .B2(new_n842), .ZN(G311));
  INV_X1    g418(.A(KEYINPUT93), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n842), .ZN(new_n845));
  INV_X1    g420(.A(new_n784), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g422(.A(KEYINPUT93), .B(new_n784), .C1(new_n840), .C2(new_n842), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(G150));
  NAND2_X1  g424(.A1(new_n601), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n523), .A2(G93), .B1(new_n515), .B2(G55), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n536), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n541), .B2(new_n853), .ZN(new_n854));
  OR3_X1    g429(.A1(new_n551), .A2(new_n854), .A3(new_n552), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n551), .B2(new_n552), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n851), .B(new_n857), .Z(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n860));
  XNOR2_X1  g435(.A(KEYINPUT94), .B(G860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n861), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n854), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(G145));
  INV_X1    g441(.A(G37), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT95), .B1(new_n503), .B2(new_n504), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n498), .B1(new_n501), .B2(new_n500), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT4), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT95), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n502), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n464), .A2(KEYINPUT70), .A3(G114), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n493), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT71), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n491), .A2(new_n486), .A3(new_n493), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n877), .A2(new_n878), .B1(G126), .B2(new_n474), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n723), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n833), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n463), .A2(G142), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n474), .A2(G130), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n464), .A2(G118), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n883), .B(new_n884), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n616), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n757), .B(KEYINPUT96), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n737), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n889), .A2(new_n737), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  INV_X1    g469(.A(new_n888), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n882), .B(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n472), .B(new_n623), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n483), .B(new_n899), .Z(new_n900));
  OAI21_X1  g475(.A(new_n867), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n898), .B2(new_n900), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT98), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n906), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n904), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT98), .A3(new_n902), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n909), .A2(new_n912), .A3(KEYINPUT40), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT40), .B1(new_n909), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(G395));
  NAND2_X1  g490(.A1(G166), .A2(G290), .ZN(new_n916));
  NAND2_X1  g491(.A1(G303), .A2(new_n589), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G288), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n579), .B2(new_n582), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n579), .A2(new_n582), .A3(new_n919), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(G305), .A2(G288), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n924), .A2(new_n920), .A3(new_n917), .A4(new_n916), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(new_n925), .A3(KEYINPUT102), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT102), .B1(new_n923), .B2(new_n925), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n927), .B1(new_n932), .B2(KEYINPUT42), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n609), .B(new_n857), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n600), .A2(new_n566), .A3(KEYINPUT99), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n600), .A2(new_n566), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n593), .B(new_n599), .C1(new_n561), .C2(new_n565), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(KEYINPUT99), .A3(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n935), .A2(new_n938), .A3(KEYINPUT100), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT100), .B1(new_n935), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT41), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n935), .B2(new_n938), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n936), .A2(new_n937), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(new_n942), .ZN(new_n946));
  AOI211_X1 g521(.A(KEYINPUT101), .B(KEYINPUT41), .C1(new_n936), .C2(new_n937), .ZN(new_n947));
  OR3_X1    g522(.A1(new_n943), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n941), .B1(new_n948), .B2(new_n934), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n933), .B(new_n949), .ZN(new_n950));
  MUX2_X1   g525(.A(new_n854), .B(new_n950), .S(G868), .Z(G295));
  MUX2_X1   g526(.A(new_n854), .B(new_n950), .S(G868), .Z(G331));
  XNOR2_X1  g527(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n855), .A2(G301), .A3(new_n856), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(G301), .B1(new_n855), .B2(new_n856), .ZN(new_n957));
  OAI21_X1  g532(.A(G286), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n957), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(G168), .A3(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n935), .A2(new_n938), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n943), .A2(new_n946), .A3(new_n947), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n964), .B(KEYINPUT104), .C1(new_n965), .C2(new_n961), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n961), .A2(new_n967), .A3(new_n963), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(G37), .B1(new_n969), .B2(new_n931), .ZN(new_n970));
  INV_X1    g545(.A(new_n968), .ZN(new_n971));
  INV_X1    g546(.A(new_n961), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n948), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n967), .B1(new_n961), .B2(new_n963), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT105), .B1(new_n929), .B2(new_n930), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT102), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n926), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n928), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n975), .A2(new_n976), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n954), .B1(new_n970), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n932), .B1(new_n966), .B2(new_n968), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n961), .B1(new_n939), .B2(new_n940), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n935), .A2(new_n938), .A3(new_n942), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n936), .A2(KEYINPUT41), .A3(new_n937), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n958), .A2(new_n960), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n976), .A2(new_n984), .A3(new_n980), .A4(new_n987), .ZN(new_n988));
  NOR4_X1   g563(.A1(new_n983), .A2(new_n988), .A3(KEYINPUT43), .A4(G37), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n953), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n867), .B1(new_n975), .B2(new_n932), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT43), .B1(new_n991), .B2(new_n988), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n970), .A2(new_n981), .A3(new_n954), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n993), .A3(KEYINPUT44), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n990), .A2(new_n994), .ZN(G397));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n880), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n469), .B(G40), .C1(new_n464), .C2(new_n471), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1986), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n589), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT107), .Z(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n1002), .B2(new_n589), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n723), .B(G1996), .ZN(new_n1007));
  INV_X1    g582(.A(G2067), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n757), .B(new_n1008), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n834), .A2(new_n836), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n834), .A2(new_n836), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1001), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT60), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n601), .B2(KEYINPUT120), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n870), .A2(new_n871), .A3(new_n502), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n871), .B1(new_n870), .B2(new_n502), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1016), .B(new_n996), .C1(new_n1019), .C2(new_n496), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n996), .B1(new_n496), .B2(new_n505), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT50), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1000), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT116), .ZN(new_n1025));
  INV_X1    g600(.A(G1348), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1020), .A2(new_n1022), .A3(new_n1027), .A4(new_n1023), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n873), .B2(new_n879), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(new_n1008), .A3(new_n1023), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1029), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1030), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1015), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n600), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT117), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1029), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1014), .A3(new_n1042), .ZN(new_n1043));
  OAI221_X1 g618(.A(new_n1015), .B1(KEYINPUT120), .B2(new_n601), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1000), .B1(new_n1021), .B2(new_n998), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT45), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT108), .B1(new_n997), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT108), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1031), .A2(new_n1050), .A3(KEYINPUT45), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1047), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT56), .B(G2072), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1023), .B1(new_n1021), .B2(KEYINPUT50), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(KEYINPUT50), .B2(new_n997), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1056), .A2(G1956), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n566), .B(KEYINPUT57), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1058), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT61), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1058), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT61), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n1059), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1031), .A2(new_n1050), .A3(KEYINPUT45), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1050), .B1(new_n1031), .B2(KEYINPUT45), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1046), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI211_X1 g645(.A(G1384), .B(new_n1000), .C1(new_n879), .C2(new_n873), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT58), .B(G1341), .ZN(new_n1072));
  OAI22_X1  g647(.A1(new_n1070), .A2(G1996), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n553), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1075));
  OR2_X1    g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1062), .A2(new_n1067), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1041), .A2(new_n601), .A3(new_n1042), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT118), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1041), .A2(new_n1081), .A3(new_n601), .A4(new_n1042), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(new_n1082), .A3(new_n1065), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1045), .A2(new_n1078), .B1(new_n1083), .B2(new_n1059), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1070), .B2(G2078), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1025), .A2(new_n743), .A3(new_n1028), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n471), .A2(KEYINPUT124), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n471), .A2(KEYINPUT124), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(G2105), .ZN(new_n1091));
  AND4_X1   g666(.A1(KEYINPUT53), .A2(new_n469), .A3(G40), .A4(new_n701), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1088), .A2(new_n999), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1086), .A2(new_n1087), .A3(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1086), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1031), .A2(KEYINPUT45), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1023), .B1(new_n1021), .B2(new_n998), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(KEYINPUT53), .A3(new_n701), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1087), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1087), .A2(new_n1100), .A3(KEYINPUT123), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1096), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1095), .B1(new_n1105), .B2(G301), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1087), .A2(new_n1100), .A3(KEYINPUT123), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT123), .B1(new_n1087), .B2(new_n1100), .ZN(new_n1110));
  OAI211_X1 g685(.A(G301), .B(new_n1086), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(KEYINPUT125), .A3(G301), .A4(new_n1086), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1107), .B1(new_n1094), .B2(G171), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(G1981), .B1(new_n580), .B2(new_n577), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT111), .B(G1981), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n578), .A2(new_n573), .A3(new_n574), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT49), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT110), .ZN(new_n1123));
  INV_X1    g698(.A(G8), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1123), .B(new_n1124), .C1(new_n1031), .C2(new_n1023), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n880), .A2(new_n996), .A3(new_n1023), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT110), .B1(new_n1126), .B2(G8), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1122), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n919), .A2(G1976), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT52), .B1(G288), .B2(new_n795), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1129), .B(new_n1130), .C1(new_n1125), .C2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT52), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1123), .B1(new_n1071), .B2(new_n1124), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1126), .A2(KEYINPUT110), .A3(G8), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1136), .B2(new_n1129), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1132), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(G303), .A2(G8), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT55), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT109), .B(G1971), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1070), .A2(new_n1142), .B1(new_n777), .B2(new_n1056), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1140), .B1(new_n1143), .B2(new_n1124), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1140), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1141), .B1(new_n1088), .B2(new_n1046), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1024), .A2(G2090), .ZN(new_n1147));
  OAI211_X1 g722(.A(G8), .B(new_n1145), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1138), .A2(new_n1144), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(G1966), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n1152));
  INV_X1    g727(.A(G2084), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1020), .A2(new_n1022), .A3(new_n1153), .A4(new_n1023), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1152), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(G168), .A2(new_n1124), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT122), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT121), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1162));
  AND4_X1   g737(.A1(KEYINPUT122), .A2(new_n1161), .A3(new_n1162), .A4(new_n1158), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(G168), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT51), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n1124), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1160), .A2(G8), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1158), .A2(KEYINPUT51), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1149), .B1(new_n1164), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1108), .A2(new_n1117), .A3(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1084), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1169), .A2(G286), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1138), .A2(new_n1144), .A3(new_n1148), .A4(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(KEYINPUT112), .B(KEYINPUT63), .Z(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT113), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT113), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1177), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1138), .A2(new_n1148), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1176), .A2(KEYINPUT63), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1147), .B1(new_n1070), .B2(new_n1142), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1185), .A2(new_n1124), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1186), .A2(KEYINPUT114), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1140), .B1(new_n1186), .B2(KEYINPUT114), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1183), .B(new_n1184), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1180), .A2(new_n1182), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1164), .A2(new_n1191), .A3(new_n1172), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1149), .A2(new_n1105), .A3(G301), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1157), .A2(KEYINPUT122), .A3(new_n1158), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1161), .A2(new_n1162), .A3(new_n1158), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT122), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1165), .A2(new_n1167), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT62), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1192), .A2(new_n1193), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1148), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1128), .A2(new_n795), .A3(new_n919), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n1120), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n1202), .A2(new_n1138), .B1(new_n1204), .B2(new_n1136), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1190), .A2(new_n1201), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1013), .B1(new_n1175), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1208));
  OAI22_X1  g783(.A1(new_n1208), .A2(new_n1011), .B1(G2067), .B2(new_n757), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n1209), .A2(new_n1001), .ZN(new_n1210));
  OR3_X1    g785(.A1(new_n999), .A2(G1996), .A3(new_n1000), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT46), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1009), .A2(new_n723), .ZN(new_n1213));
  AOI22_X1  g788(.A1(new_n1211), .A2(new_n1212), .B1(new_n1001), .B2(new_n1213), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1215));
  AND2_X1   g790(.A1(new_n1215), .A2(KEYINPUT126), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1215), .A2(KEYINPUT126), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1214), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(KEYINPUT47), .ZN(new_n1219));
  OR2_X1    g794(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1004), .A2(new_n1001), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n1221), .B(KEYINPUT127), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT48), .ZN(new_n1223));
  OR2_X1    g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1001), .A2(new_n1012), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1220), .A2(new_n1227), .ZN(new_n1228));
  AOI211_X1 g803(.A(new_n1210), .B(new_n1228), .C1(new_n1219), .C2(new_n1218), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1207), .A2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g805(.A1(new_n982), .A2(new_n989), .ZN(new_n1232));
  INV_X1    g806(.A(G319), .ZN(new_n1233));
  NOR2_X1   g807(.A1(G227), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g808(.A1(new_n645), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g809(.A(new_n1235), .B1(new_n691), .B2(new_n692), .ZN(new_n1236));
  NOR2_X1   g810(.A1(new_n907), .A2(new_n908), .ZN(new_n1237));
  AOI21_X1  g811(.A(KEYINPUT98), .B1(new_n911), .B2(new_n902), .ZN(new_n1238));
  OAI21_X1  g812(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g813(.A1(new_n1232), .A2(new_n1239), .ZN(G308));
  OAI221_X1 g814(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .C1(new_n982), .C2(new_n989), .ZN(G225));
endmodule


