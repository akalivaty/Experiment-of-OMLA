//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n589,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT68), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT70), .Z(G217));
  NOR4_X1   g027(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT71), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT72), .A2(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT72), .A2(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT73), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n469), .A2(new_n470), .B1(G113), .B2(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT73), .A4(G125), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n465), .A2(KEYINPUT74), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT74), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(G101), .A3(new_n478), .ZN(new_n479));
  OR2_X1    g054(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(G2104), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n474), .A2(new_n476), .A3(KEYINPUT3), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G137), .ZN(new_n485));
  NOR3_X1   g060(.A1(new_n462), .A2(new_n463), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n479), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n473), .A2(new_n488), .ZN(G160));
  NOR2_X1   g064(.A1(new_n484), .A2(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n464), .C2(G112), .ZN(new_n492));
  INV_X1    g067(.A(G136), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT74), .B(G2104), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(KEYINPUT75), .B2(KEYINPUT3), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n494), .A2(KEYINPUT3), .B1(new_n496), .B2(new_n481), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n478), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n491), .B(new_n492), .C1(new_n493), .C2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G162));
  NOR2_X1   g075(.A1(new_n478), .A2(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n503), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  NOR3_X1   g083(.A1(new_n462), .A2(new_n463), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n497), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n466), .A2(new_n468), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n513), .A2(new_n509), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n506), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n517), .A2(G62), .ZN(new_n518));
  AND2_X1   g093(.A1(G75), .A2(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(G651), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT77), .B1(new_n521), .B2(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT77), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT6), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT78), .B1(new_n524), .B2(KEYINPUT6), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(new_n521), .A3(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n526), .A2(new_n530), .A3(G88), .A4(new_n517), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n520), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n526), .A2(new_n530), .A3(G50), .A4(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(KEYINPUT79), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(KEYINPUT79), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(G166));
  AND2_X1   g111(.A1(new_n526), .A2(new_n530), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n526), .A2(new_n530), .A3(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  AND2_X1   g116(.A1(KEYINPUT5), .A2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(KEYINPUT5), .A2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(G651), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n545), .A2(G63), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n539), .A2(new_n541), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT80), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT80), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n539), .A2(new_n552), .A3(new_n541), .A4(new_n549), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(G168));
  NAND2_X1  g129(.A1(new_n538), .A2(G90), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n540), .A2(G52), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n524), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(G301));
  INV_X1    g134(.A(G301), .ZN(G171));
  NAND2_X1  g135(.A1(new_n540), .A2(G43), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n537), .A2(G81), .A3(new_n517), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(new_n524), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n561), .A2(new_n562), .A3(new_n564), .A4(KEYINPUT81), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G860), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT82), .ZN(G153));
  NAND4_X1  g147(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  AND4_X1   g151(.A1(G91), .A2(new_n526), .A3(new_n530), .A4(new_n517), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n517), .A2(G65), .ZN(new_n578));
  AND2_X1   g153(.A1(G78), .A2(G543), .ZN(new_n579));
  OAI211_X1 g154(.A(KEYINPUT83), .B(G651), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n579), .B1(new_n517), .B2(G65), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(new_n524), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n577), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n526), .A2(new_n530), .A3(G53), .A4(G543), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT9), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G299));
  AND2_X1   g162(.A1(new_n551), .A2(new_n553), .ZN(G286));
  NAND2_X1  g163(.A1(new_n534), .A2(new_n535), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n589), .A2(new_n531), .A3(new_n520), .ZN(G303));
  NAND4_X1  g165(.A1(new_n526), .A2(new_n530), .A3(G87), .A4(new_n517), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n526), .A2(new_n530), .A3(G49), .A4(G543), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n593), .B(G651), .C1(new_n517), .C2(G74), .ZN(new_n594));
  NAND2_X1  g169(.A1(G74), .A2(G651), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n544), .A2(KEYINPUT84), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n591), .A2(new_n592), .A3(new_n594), .A4(new_n596), .ZN(G288));
  NAND4_X1  g172(.A1(new_n526), .A2(new_n530), .A3(G86), .A4(new_n517), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n526), .A2(new_n530), .A3(G48), .A4(G543), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  OR2_X1    g175(.A1(KEYINPUT5), .A2(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(KEYINPUT5), .A2(G543), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g178(.A1(G73), .A2(G543), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n598), .A2(new_n599), .A3(new_n605), .ZN(G305));
  NAND2_X1  g181(.A1(new_n540), .A2(G47), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n537), .A2(new_n517), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  OAI221_X1 g185(.A(new_n607), .B1(new_n524), .B2(new_n608), .C1(new_n609), .C2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n538), .A2(KEYINPUT10), .A3(G92), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n540), .A2(G54), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n524), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n612), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n612), .B1(new_n621), .B2(G868), .ZN(G321));
  NOR2_X1   g198(.A1(G299), .A2(G868), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g200(.A(new_n624), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n621), .B1(new_n627), .B2(G860), .ZN(G148));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n569), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n621), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n631), .A2(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n630), .B1(new_n632), .B2(new_n629), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT85), .Z(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g210(.A1(new_n494), .A2(G2105), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n636), .A2(new_n466), .A3(new_n468), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2100), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n490), .A2(G123), .ZN(new_n642));
  OAI221_X1 g217(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n643));
  INV_X1    g218(.A(G135), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n498), .ZN(new_n645));
  INV_X1    g220(.A(G2096), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n641), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT87), .Z(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n657), .B(new_n658), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(new_n663), .A3(G14), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT88), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(new_n646), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  INV_X1    g261(.A(new_n681), .ZN(new_n687));
  INV_X1    g262(.A(new_n684), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(new_n683), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n686), .B(new_n690), .C1(new_n687), .C2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G25), .ZN(new_n699));
  INV_X1    g274(.A(new_n498), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G131), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n490), .A2(G119), .ZN(new_n702));
  OAI221_X1 g277(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(new_n698), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(G24), .B(G290), .S(G16), .Z(new_n709));
  XOR2_X1   g284(.A(KEYINPUT90), .B(G1986), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT91), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n709), .B(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(G16), .A2(G23), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT92), .Z(new_n714));
  NAND2_X1  g289(.A1(G288), .A2(KEYINPUT93), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n594), .A2(new_n596), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n716), .A2(new_n717), .A3(new_n591), .A4(new_n592), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT33), .B(G1976), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(G22), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G166), .B2(new_n720), .ZN(new_n725));
  INV_X1    g300(.A(G1971), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  MUX2_X1   g302(.A(G6), .B(G305), .S(G16), .Z(new_n728));
  XOR2_X1   g303(.A(KEYINPUT32), .B(G1981), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n723), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n708), .B(new_n712), .C1(new_n731), .C2(KEYINPUT34), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT94), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT95), .A2(KEYINPUT36), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(G160), .A2(G29), .ZN(new_n738));
  INV_X1    g313(.A(G34), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(KEYINPUT24), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n739), .B2(KEYINPUT24), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(KEYINPUT96), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(KEYINPUT96), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2084), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n720), .A2(G5), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G171), .B2(new_n720), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n490), .A2(G129), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT26), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n636), .A2(G105), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G141), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n748), .B(new_n753), .C1(new_n754), .C2(new_n498), .ZN(new_n755));
  MUX2_X1   g330(.A(G32), .B(new_n755), .S(G29), .Z(new_n756));
  XOR2_X1   g331(.A(KEYINPUT27), .B(G1996), .Z(new_n757));
  OAI221_X1 g332(.A(new_n745), .B1(G1961), .B2(new_n747), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n698), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n698), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2090), .ZN(new_n762));
  INV_X1    g337(.A(G1341), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n720), .A2(G19), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n569), .B2(G16), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n758), .B(new_n762), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n747), .A2(G1961), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT99), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n720), .A2(G21), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G168), .B2(new_n720), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n770), .A2(G1966), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(G1966), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n765), .A2(new_n763), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n768), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G4), .A2(G16), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n621), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1348), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n720), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT23), .ZN(new_n779));
  INV_X1    g354(.A(G299), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n720), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1956), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n645), .A2(new_n698), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT97), .ZN(new_n785));
  INV_X1    g360(.A(G2078), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n698), .A2(G27), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT100), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n515), .B2(G29), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n785), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G11), .ZN(new_n791));
  INV_X1    g366(.A(G28), .ZN(new_n792));
  AOI21_X1  g367(.A(G29), .B1(new_n792), .B2(KEYINPUT30), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(KEYINPUT30), .B2(new_n792), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n793), .A2(KEYINPUT98), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n698), .A2(G33), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT25), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n700), .A2(G139), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n466), .A2(new_n468), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n802), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n800), .B(new_n801), .C1(new_n464), .C2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n798), .B1(new_n804), .B2(G29), .ZN(new_n805));
  INV_X1    g380(.A(G2072), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n797), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n806), .B2(new_n805), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n756), .A2(new_n757), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n789), .A2(new_n786), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n698), .A2(G26), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT28), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n490), .A2(G128), .ZN(new_n814));
  OAI221_X1 g389(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n815));
  INV_X1    g390(.A(G140), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n814), .B(new_n815), .C1(new_n816), .C2(new_n498), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n813), .B1(new_n817), .B2(G29), .ZN(new_n818));
  INV_X1    g393(.A(G2067), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n790), .A2(new_n808), .A3(new_n811), .A4(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n766), .A2(new_n774), .A3(new_n783), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n737), .A2(new_n822), .ZN(G311));
  INV_X1    g398(.A(G311), .ZN(G150));
  NAND2_X1  g399(.A1(new_n540), .A2(G55), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  OAI221_X1 g402(.A(new_n825), .B1(new_n524), .B2(new_n826), .C1(new_n609), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n569), .A2(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(new_n565), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT38), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n621), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n570), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n828), .A2(G860), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT101), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n837), .A2(new_n840), .ZN(G145));
  INV_X1    g416(.A(G37), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n645), .B(G160), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G162), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n704), .B(KEYINPUT102), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n490), .A2(G130), .ZN(new_n846));
  OAI221_X1 g421(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n464), .C2(G118), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G142), .B2(new_n700), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n845), .B(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n639), .Z(new_n851));
  XNOR2_X1  g426(.A(G164), .B(new_n817), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n755), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n804), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n851), .A2(new_n854), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n844), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n844), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n859), .B2(new_n856), .ZN(new_n860));
  INV_X1    g435(.A(new_n856), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(KEYINPUT103), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n842), .B(new_n857), .C1(new_n860), .C2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g439(.A1(new_n828), .A2(new_n629), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n632), .B(new_n831), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n631), .A2(new_n780), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT104), .B1(new_n621), .B2(G299), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n621), .A2(G299), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n869), .A2(new_n874), .A3(new_n870), .A4(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  OR3_X1    g451(.A1(new_n867), .A2(new_n876), .A3(KEYINPUT105), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT105), .B1(new_n867), .B2(new_n876), .ZN(new_n878));
  INV_X1    g453(.A(new_n872), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n877), .B(new_n878), .C1(new_n866), .C2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G303), .B(new_n719), .ZN(new_n881));
  XNOR2_X1  g456(.A(G290), .B(G305), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n880), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n865), .B1(new_n885), .B2(new_n629), .ZN(G295));
  OAI21_X1  g461(.A(new_n865), .B1(new_n885), .B2(new_n629), .ZN(G331));
  NOR2_X1   g462(.A1(G168), .A2(G301), .ZN(new_n888));
  AOI21_X1  g463(.A(G171), .B1(new_n551), .B2(new_n553), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n829), .B(new_n830), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(G286), .A2(G171), .ZN(new_n891));
  INV_X1    g466(.A(new_n889), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n831), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n893), .A3(KEYINPUT106), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n891), .A2(new_n895), .A3(new_n831), .A4(new_n892), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n894), .A2(new_n873), .A3(new_n875), .A4(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n872), .A2(new_n890), .A3(new_n893), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n883), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n842), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n883), .B1(new_n897), .B2(new_n898), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n899), .A2(new_n842), .ZN(new_n903));
  INV_X1    g478(.A(new_n883), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n890), .A2(new_n893), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n905), .A2(new_n873), .A3(new_n875), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n879), .B1(new_n894), .B2(new_n896), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT107), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n910), .B(new_n904), .C1(new_n906), .C2(new_n907), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n903), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n902), .B1(new_n912), .B2(KEYINPUT43), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(KEYINPUT44), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n912), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n918));
  OR3_X1    g493(.A1(new_n900), .A2(KEYINPUT43), .A3(new_n901), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n914), .B1(new_n920), .B2(KEYINPUT44), .ZN(G397));
  NAND3_X1  g496(.A1(new_n509), .A2(new_n483), .A3(new_n482), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT4), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n513), .A2(new_n509), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G1384), .B1(new_n925), .B2(new_n506), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n469), .A2(new_n470), .ZN(new_n927));
  NAND2_X1  g502(.A1(G113), .A2(G2104), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n472), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n464), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n497), .A2(new_n486), .B1(new_n636), .B2(G101), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(G40), .A3(new_n932), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n926), .A2(KEYINPUT45), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n817), .B(new_n819), .ZN(new_n935));
  INV_X1    g510(.A(G1996), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n755), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n704), .B(new_n707), .Z(new_n939));
  OAI21_X1  g514(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(G290), .A2(G1986), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n934), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n943), .A2(KEYINPUT48), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(KEYINPUT48), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n941), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n935), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n934), .B1(new_n947), .B2(new_n755), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n934), .A2(new_n936), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(KEYINPUT46), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n949), .A2(KEYINPUT46), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n952), .B(KEYINPUT47), .Z(new_n953));
  NAND2_X1  g528(.A1(new_n705), .A2(new_n707), .ZN(new_n954));
  OAI22_X1  g529(.A1(new_n938), .A2(new_n954), .B1(G2067), .B2(new_n817), .ZN(new_n955));
  AOI211_X1 g530(.A(new_n946), .B(new_n953), .C1(new_n934), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n922), .A2(KEYINPUT4), .B1(new_n513), .B2(new_n509), .ZN(new_n958));
  OAI22_X1  g533(.A1(new_n484), .A2(new_n504), .B1(new_n501), .B2(new_n502), .ZN(new_n959));
  OAI211_X1 g534(.A(KEYINPUT45), .B(new_n957), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n933), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT117), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT45), .B1(new_n515), .B2(new_n957), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT117), .B1(new_n967), .B2(new_n933), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1966), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n515), .A2(new_n973), .A3(new_n957), .ZN(new_n974));
  INV_X1    g549(.A(G40), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n473), .A2(new_n488), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(G2084), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n971), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT110), .B(G8), .Z(new_n981));
  NOR2_X1   g556(.A1(G168), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n984));
  INV_X1    g559(.A(new_n982), .ZN(new_n985));
  AOI21_X1  g560(.A(G1966), .B1(new_n966), .B2(new_n968), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(new_n978), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n984), .B(new_n985), .C1(new_n987), .C2(new_n981), .ZN(new_n988));
  OAI21_X1  g563(.A(G8), .B1(new_n986), .B2(new_n978), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n984), .B1(new_n989), .B2(new_n985), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT125), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI211_X1 g567(.A(KEYINPUT125), .B(new_n984), .C1(new_n989), .C2(new_n985), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n983), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n964), .A2(new_n786), .A3(new_n960), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n998));
  INV_X1    g573(.A(G1961), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n997), .A2(new_n998), .B1(new_n977), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n998), .A2(G2078), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n966), .A2(new_n968), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G171), .ZN(new_n1004));
  INV_X1    g579(.A(new_n981), .ZN(new_n1005));
  INV_X1    g580(.A(G2090), .ZN(new_n1006));
  AND4_X1   g581(.A1(new_n1006), .A2(new_n972), .A3(new_n974), .A4(new_n976), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1971), .B1(new_n964), .B2(new_n960), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(G166), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(KEYINPUT113), .A2(G86), .ZN(new_n1017));
  NOR2_X1   g592(.A1(KEYINPUT113), .A2(G86), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n526), .A2(new_n530), .A3(new_n517), .A4(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n599), .A2(new_n1020), .A3(new_n605), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(G1981), .ZN(new_n1022));
  INV_X1    g597(.A(G1981), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n598), .A2(new_n599), .A3(new_n605), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(KEYINPUT49), .A3(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1025), .B(new_n1005), .C1(new_n933), .C2(new_n962), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT49), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT114), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n981), .B1(new_n926), .B2(new_n976), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1027), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1025), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n715), .A2(new_n718), .A3(G1976), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1028), .A2(new_n1032), .B1(KEYINPUT52), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n926), .A2(new_n976), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT111), .B(G1976), .Z(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1036), .A2(new_n1033), .A3(new_n1005), .A4(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT112), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1029), .A2(new_n1041), .A3(new_n1033), .A4(new_n1038), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1014), .B(G8), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1016), .A2(new_n1035), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NOR4_X1   g620(.A1(new_n995), .A2(new_n996), .A3(new_n1004), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT127), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n997), .A2(new_n998), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n977), .A2(new_n999), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n964), .A2(new_n960), .A3(new_n1001), .ZN(new_n1050));
  AND4_X1   g625(.A1(G301), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT126), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1051), .A2(new_n1052), .B1(G171), .B2(new_n1003), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT126), .B1(new_n1054), .B2(G171), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT54), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(G171), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1000), .A2(new_n1002), .A3(G301), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(KEYINPUT54), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1043), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1059), .A2(new_n1063), .A3(new_n1016), .A4(new_n1044), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1056), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n994), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1036), .A2(G2067), .ZN(new_n1067));
  INV_X1    g642(.A(G1348), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n977), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1069), .A2(KEYINPUT60), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n621), .A2(KEYINPUT124), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n621), .A2(KEYINPUT124), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1069), .A2(KEYINPUT60), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n964), .A2(new_n936), .A3(new_n960), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n1036), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n567), .A2(KEYINPUT122), .A3(new_n568), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1078), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  AOI211_X1 g660(.A(KEYINPUT59), .B(new_n1083), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n584), .A2(new_n586), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n584), .B2(new_n586), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1956), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n977), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT120), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n977), .A2(new_n1095), .A3(new_n1092), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n964), .A2(new_n960), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1091), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1091), .A2(new_n1099), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n977), .A2(new_n1095), .A3(new_n1092), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1095), .B1(new_n977), .B2(new_n1092), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT61), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1087), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1099), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1091), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT61), .B1(new_n1109), .B2(new_n1104), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1106), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n1115), .B2(new_n1109), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1104), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1114), .B1(new_n1100), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT123), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1077), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1069), .A2(new_n631), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1104), .B1(new_n1100), .B2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(KEYINPUT121), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1066), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n972), .A2(new_n974), .A3(new_n1006), .A4(new_n976), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n967), .A2(new_n961), .A3(new_n933), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(G1971), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1014), .B1(new_n1127), .B2(G8), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT118), .B1(new_n1062), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(G168), .B(new_n1005), .C1(new_n986), .C2(new_n978), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1044), .A2(KEYINPUT63), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1015), .B1(new_n1133), .B2(new_n1012), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1134), .A2(new_n1135), .A3(new_n1043), .A4(new_n1035), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1129), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1045), .B2(new_n1130), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1062), .A2(new_n1044), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1005), .B1(new_n962), .B2(new_n933), .ZN(new_n1142));
  NOR2_X1   g717(.A1(G288), .A2(G1976), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1022), .A2(KEYINPUT49), .A3(new_n1024), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1031), .B1(new_n1145), .B2(new_n1030), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1026), .A2(KEYINPUT114), .A3(new_n1027), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1143), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1024), .B(KEYINPUT115), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1142), .B1(new_n1150), .B2(KEYINPUT116), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT116), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1148), .A2(new_n1152), .A3(new_n1149), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1141), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1140), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n1140), .B2(new_n1154), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1047), .B1(new_n1124), .B2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1000), .A2(new_n1052), .A3(G301), .A4(new_n1050), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1055), .A2(new_n1004), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT54), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1045), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n1059), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n982), .B1(new_n980), .B2(G8), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT125), .B1(new_n1166), .B2(new_n984), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n990), .A2(new_n991), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(new_n988), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1165), .B1(new_n1169), .B2(new_n983), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1111), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1116), .A2(new_n1118), .A3(KEYINPUT123), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1076), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1122), .B(KEYINPUT121), .Z(new_n1174));
  OAI21_X1  g749(.A(new_n1170), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1140), .A2(new_n1154), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT119), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1140), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1175), .A2(new_n1179), .A3(KEYINPUT127), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1046), .B1(new_n1159), .B2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(G290), .B(G1986), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n941), .B1(new_n934), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT109), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n956), .B1(new_n1181), .B2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g760(.A(G319), .ZN(new_n1187));
  NOR4_X1   g761(.A1(G229), .A2(G401), .A3(new_n1187), .A4(G227), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n863), .A2(new_n913), .A3(new_n1188), .ZN(G225));
  INV_X1    g763(.A(G225), .ZN(G308));
endmodule


