//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950;
  XOR2_X1   g000(.A(G183gat), .B(G211gat), .Z(new_n202));
  NAND2_X1  g001(.A1(G231gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G15gat), .B(G22gat), .Z(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(KEYINPUT99), .A2(G8gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(KEYINPUT97), .A2(G1gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(KEYINPUT97), .A2(G1gat), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n213), .A2(KEYINPUT16), .A3(new_n214), .ZN(new_n215));
  OR3_X1    g014(.A1(new_n215), .A2(new_n208), .A3(KEYINPUT98), .ZN(new_n216));
  NAND2_X1  g015(.A1(KEYINPUT99), .A2(G8gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT98), .B1(new_n215), .B2(new_n208), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n212), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n215), .A2(new_n208), .ZN(new_n220));
  OAI21_X1  g019(.A(G8gat), .B1(new_n220), .B2(new_n210), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G57gat), .B(G64gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G71gat), .B(G78gat), .Z(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n222), .B1(KEYINPUT21), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT104), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT103), .B(KEYINPUT19), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n227), .A2(KEYINPUT21), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n232), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(G127gat), .B(G155gat), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n235), .A2(new_n236), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n207), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n239), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n237), .A3(new_n206), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(G43gat), .B(G50gat), .Z(new_n244));
  INV_X1    g043(.A(KEYINPUT15), .ZN(new_n245));
  INV_X1    g044(.A(G29gat), .ZN(new_n246));
  INV_X1    g045(.A(G36gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n244), .A2(new_n245), .B1(KEYINPUT96), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n247), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT14), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n249), .B(new_n251), .C1(KEYINPUT96), .C2(new_n248), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n244), .A2(new_n245), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT17), .ZN(new_n255));
  INV_X1    g054(.A(G85gat), .ZN(new_n256));
  INV_X1    g055(.A(G92gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT7), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT7), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(G85gat), .A3(G92gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(G99gat), .A2(G106gat), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n258), .A2(new_n260), .B1(KEYINPUT8), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(G85gat), .B2(G92gat), .ZN(new_n263));
  XOR2_X1   g062(.A(G99gat), .B(G106gat), .Z(new_n264));
  XOR2_X1   g063(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n255), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n254), .A2(new_n265), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT41), .ZN(new_n269));
  NAND2_X1  g068(.A1(G232gat), .A2(G233gat), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n267), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G190gat), .B(G218gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G134gat), .B(G162gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n269), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n273), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n243), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT89), .ZN(new_n280));
  XNOR2_X1  g079(.A(G155gat), .B(G162gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G141gat), .B(G148gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(KEYINPUT2), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT81), .ZN(new_n286));
  AND2_X1   g085(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n288));
  INV_X1    g087(.A(G155gat), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT2), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n282), .A2(new_n283), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT80), .B(G162gat), .ZN(new_n294));
  OAI211_X1 g093(.A(KEYINPUT81), .B(KEYINPUT2), .C1(new_n294), .C2(new_n289), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT82), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT82), .A4(new_n295), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n285), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT3), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT29), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT76), .ZN(new_n303));
  INV_X1    g102(.A(G197gat), .ZN(new_n304));
  INV_X1    g103(.A(G204gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G197gat), .A2(G204gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G211gat), .A2(G218gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT22), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G211gat), .B(G218gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n303), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n306), .A2(new_n307), .B1(new_n310), .B2(new_n309), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(KEYINPUT76), .A3(new_n313), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n312), .A2(KEYINPUT75), .A3(new_n314), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n316), .B2(new_n313), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n280), .B1(new_n302), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n323), .B(KEYINPUT77), .ZN(new_n327));
  AOI211_X1 g126(.A(KEYINPUT3), .B(new_n285), .C1(new_n298), .C2(new_n299), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n327), .B(KEYINPUT89), .C1(new_n328), .C2(KEYINPUT29), .ZN(new_n329));
  INV_X1    g128(.A(G228gat), .ZN(new_n330));
  INV_X1    g129(.A(G233gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n326), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n298), .A2(new_n299), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n284), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT29), .B1(new_n318), .B2(new_n322), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(KEYINPUT3), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT88), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT87), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n302), .B2(new_n323), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n315), .A2(new_n317), .B1(new_n314), .B2(new_n312), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n301), .B1(new_n341), .B2(KEYINPUT29), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n323), .ZN(new_n344));
  OAI211_X1 g143(.A(KEYINPUT87), .B(new_n344), .C1(new_n328), .C2(KEYINPUT29), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n332), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n333), .A2(new_n338), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G22gat), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT91), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G78gat), .B(G106gat), .ZN(new_n351));
  INV_X1    g150(.A(G50gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  XOR2_X1   g154(.A(KEYINPUT90), .B(G22gat), .Z(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n348), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT91), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n346), .A2(new_n347), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT88), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n337), .B(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n326), .A2(new_n329), .A3(new_n332), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n359), .B(G22gat), .C1(new_n361), .C2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n358), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n333), .A2(new_n338), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n368), .A2(new_n357), .A3(new_n360), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n357), .B1(new_n368), .B2(new_n360), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n355), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n300), .A2(new_n301), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT72), .ZN(new_n374));
  INV_X1    g173(.A(G113gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(G120gat), .ZN(new_n376));
  INV_X1    g175(.A(G120gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(G113gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n374), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(G113gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(G120gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(KEYINPUT72), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT70), .B(G134gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G127gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT71), .ZN(new_n387));
  INV_X1    g186(.A(G127gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(G134gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(new_n387), .A3(G127gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n384), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G134gat), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT1), .B1(new_n393), .B2(G127gat), .ZN(new_n394));
  OAI221_X1 g193(.A(new_n394), .B1(G127gat), .B2(new_n393), .C1(new_n376), .C2(new_n378), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n373), .A2(new_n328), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n400), .B1(new_n300), .B2(new_n396), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n334), .A2(new_n403), .A3(new_n284), .A4(new_n396), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n398), .A2(new_n405), .A3(KEYINPUT5), .ZN(new_n406));
  INV_X1    g205(.A(new_n396), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n335), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n334), .A2(new_n284), .A3(new_n396), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT5), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n400), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412));
  AOI211_X1 g211(.A(new_n412), .B(new_n403), .C1(new_n300), .C2(new_n396), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT85), .B1(new_n409), .B2(KEYINPUT4), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n404), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n300), .A2(KEYINPUT84), .A3(new_n403), .A4(new_n396), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n397), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n406), .B(new_n411), .C1(new_n420), .C2(KEYINPUT5), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n422));
  XNOR2_X1  g221(.A(G57gat), .B(G85gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425));
  XOR2_X1   g224(.A(new_n424), .B(new_n425), .Z(new_n426));
  NAND2_X1  g225(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n409), .A2(KEYINPUT4), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n412), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n409), .A2(KEYINPUT85), .A3(KEYINPUT4), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n430), .A2(new_n431), .A3(new_n417), .A4(new_n418), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n398), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT5), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n426), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n406), .A4(new_n411), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n427), .A2(new_n428), .A3(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n433), .A2(new_n434), .B1(new_n400), .B2(new_n410), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n436), .A4(new_n406), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G8gat), .B(G36gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(new_n257), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT79), .B(G64gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT25), .ZN(new_n447));
  NOR2_X1   g246(.A1(G169gat), .A2(G176gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT23), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT23), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n450), .B1(G169gat), .B2(G176gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G183gat), .A2(G190gat), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT24), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n459));
  NAND3_X1  g258(.A1(KEYINPUT67), .A2(G183gat), .A3(G190gat), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n455), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n454), .A2(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT69), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n459), .A4(new_n460), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n453), .A2(new_n457), .ZN(new_n467));
  NOR2_X1   g266(.A1(G183gat), .A2(G190gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n452), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G169gat), .A2(G176gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n471), .B(KEYINPUT66), .Z(new_n472));
  AOI21_X1  g271(.A(new_n447), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT26), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n448), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT27), .B(G183gat), .ZN(new_n478));
  INV_X1    g277(.A(G190gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT28), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT28), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n482), .A3(new_n479), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n477), .A2(new_n481), .A3(new_n453), .A4(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT65), .B(G176gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(new_n450), .ZN(new_n486));
  INV_X1    g285(.A(G169gat), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT25), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT64), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n453), .B2(new_n457), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n453), .A2(new_n489), .A3(new_n457), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n469), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n488), .A2(new_n472), .A3(new_n451), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n484), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n473), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G226gat), .A2(G233gat), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n496), .B(KEYINPUT78), .Z(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n497), .A2(KEYINPUT29), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n498), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(new_n325), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n495), .A2(new_n499), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n344), .B1(new_n502), .B2(new_n498), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n446), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n500), .A2(new_n323), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n498), .A3(new_n327), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n445), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(KEYINPUT30), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n501), .A2(new_n503), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n445), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n484), .A2(new_n493), .ZN(new_n514));
  INV_X1    g313(.A(new_n472), .ZN(new_n515));
  AOI211_X1 g314(.A(new_n452), .B(new_n515), .C1(new_n466), .C2(new_n469), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n514), .B(new_n396), .C1(new_n447), .C2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G227gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(new_n331), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n407), .B1(new_n473), .B2(new_n494), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT34), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G43gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G71gat), .ZN(new_n527));
  XOR2_X1   g326(.A(KEYINPUT73), .B(G99gat), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n520), .B1(new_n517), .B2(new_n521), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(KEYINPUT33), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT32), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n521), .ZN(new_n535));
  AOI221_X4 g334(.A(new_n532), .B1(KEYINPUT33), .B2(new_n529), .C1(new_n535), .C2(new_n519), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n525), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n519), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT32), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT33), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n541), .A3(new_n529), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n531), .A2(new_n533), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n524), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n537), .A2(new_n544), .A3(KEYINPUT74), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT74), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n525), .B(new_n546), .C1(new_n536), .C2(new_n534), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n372), .A2(new_n441), .A3(new_n513), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT35), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT94), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n438), .A2(KEYINPUT93), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT93), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n427), .A2(new_n437), .A3(new_n553), .A4(new_n428), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n440), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT35), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n537), .A2(new_n544), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(new_n367), .B2(new_n371), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n556), .A2(new_n557), .A3(new_n559), .A4(new_n513), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT94), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n549), .A2(new_n561), .A3(KEYINPUT35), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n551), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n512), .B1(new_n438), .B2(new_n440), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(new_n372), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n558), .A2(KEYINPUT36), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n545), .A2(KEYINPUT36), .A3(new_n547), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n445), .B1(new_n509), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n570), .B2(new_n509), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n572), .A2(KEYINPUT38), .B1(new_n509), .B2(new_n445), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT38), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n500), .A2(new_n327), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n575), .B(KEYINPUT37), .C1(new_n344), .C2(new_n500), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  AND4_X1   g376(.A1(new_n440), .A2(new_n555), .A3(new_n573), .A4(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT39), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT92), .B1(new_n433), .B2(new_n400), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n581));
  AOI211_X1 g380(.A(new_n581), .B(new_n399), .C1(new_n432), .C2(new_n398), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n579), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n420), .B2(new_n399), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n433), .A2(KEYINPUT92), .A3(new_n400), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n579), .B1(new_n408), .B2(new_n401), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n583), .A2(new_n426), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT40), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n583), .A2(KEYINPUT40), .A3(new_n426), .A4(new_n587), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n590), .A2(new_n437), .A3(new_n591), .A4(new_n512), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n372), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n569), .B1(new_n578), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n279), .B1(new_n563), .B2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n222), .B(KEYINPUT100), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n255), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n254), .A2(new_n222), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G229gat), .A2(G233gat), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n602), .A2(KEYINPUT18), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n600), .B1(new_n222), .B2(new_n254), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n601), .B(KEYINPUT13), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(KEYINPUT18), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n603), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G169gat), .B(G197gat), .Z(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT95), .B(KEYINPUT11), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT12), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n603), .A2(new_n616), .A3(new_n606), .A4(new_n607), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n265), .A2(KEYINPUT10), .A3(new_n227), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n263), .A2(KEYINPUT105), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n227), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n265), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(G230gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(new_n331), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  OR3_X1    g427(.A1(new_n623), .A2(new_n626), .A3(new_n331), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n619), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n595), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n441), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT106), .B(G1gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1324gat));
  NOR2_X1   g440(.A1(new_n638), .A2(new_n513), .ZN(new_n642));
  NAND2_X1  g441(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n643));
  OR2_X1    g442(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(KEYINPUT42), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(KEYINPUT42), .ZN(new_n648));
  INV_X1    g447(.A(G8gat), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n642), .ZN(G1325gat));
  INV_X1    g449(.A(G15gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n568), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n638), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n558), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n595), .A2(new_n637), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n653), .B1(new_n651), .B2(new_n655), .ZN(G1326gat));
  NOR2_X1   g455(.A1(new_n638), .A2(new_n372), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT43), .B(G22gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  NOR3_X1   g458(.A1(new_n243), .A2(new_n619), .A3(new_n636), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n440), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(new_n552), .B2(new_n554), .ZN(new_n663));
  INV_X1    g462(.A(new_n559), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n513), .A2(new_n557), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n561), .B1(new_n549), .B2(KEYINPUT35), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n367), .A2(new_n371), .B1(new_n547), .B2(new_n545), .ZN(new_n668));
  AOI211_X1 g467(.A(KEYINPUT94), .B(new_n557), .C1(new_n668), .C2(new_n564), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n652), .B1(new_n372), .B2(new_n564), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n592), .A2(new_n372), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n663), .A2(new_n573), .A3(new_n577), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n277), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT44), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n278), .B1(new_n563), .B2(new_n594), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT108), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n278), .A2(KEYINPUT44), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n670), .A2(new_n674), .A3(KEYINPUT109), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n563), .B2(new_n594), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n682), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n661), .B1(new_n681), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n441), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT110), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n687), .A2(KEYINPUT110), .A3(new_n688), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(G29gat), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n675), .A2(new_n661), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n246), .A3(new_n688), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n693), .A2(new_n697), .ZN(G1328gat));
  NAND3_X1  g497(.A1(new_n694), .A2(new_n247), .A3(new_n512), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT111), .B(KEYINPUT46), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AOI211_X1 g500(.A(new_n513), .B(new_n661), .C1(new_n681), .C2(new_n686), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n247), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT112), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT112), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n701), .B(new_n705), .C1(new_n702), .C2(new_n247), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(G1329gat));
  AOI21_X1  g506(.A(new_n676), .B1(new_n675), .B2(KEYINPUT44), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n678), .A2(KEYINPUT108), .A3(new_n679), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n686), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n568), .A3(new_n660), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT113), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n687), .A2(KEYINPUT113), .A3(new_n568), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(G43gat), .A3(new_n714), .ZN(new_n715));
  NOR4_X1   g514(.A1(new_n675), .A2(new_n661), .A3(G43gat), .A4(new_n558), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n711), .A2(G43gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n717), .B1(new_n720), .B2(new_n716), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1330gat));
  INV_X1    g521(.A(new_n372), .ZN(new_n723));
  AOI21_X1  g522(.A(G50gat), .B1(new_n694), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n372), .A2(new_n352), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n687), .B2(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT48), .Z(G1331gat));
  NOR2_X1   g526(.A1(new_n683), .A2(new_n685), .ZN(new_n728));
  INV_X1    g527(.A(new_n636), .ZN(new_n729));
  NOR4_X1   g528(.A1(new_n728), .A2(new_n618), .A3(new_n729), .A4(new_n279), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n688), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g531(.A1(new_n728), .A2(new_n729), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n279), .A2(new_n618), .ZN(new_n734));
  NAND2_X1  g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n733), .A2(new_n512), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT114), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n730), .A2(new_n738), .A3(new_n512), .A4(new_n735), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n737), .B2(new_n739), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(G1333gat));
  NAND2_X1  g542(.A1(new_n733), .A2(new_n734), .ZN(new_n744));
  OAI21_X1  g543(.A(G71gat), .B1(new_n744), .B2(new_n652), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n746));
  INV_X1    g545(.A(G71gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n747), .A3(new_n654), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n746), .B1(new_n745), .B2(new_n748), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n730), .A2(new_n723), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n243), .A2(new_n618), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(KEYINPUT115), .B(KEYINPUT51), .C1(new_n675), .C2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n758), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n678), .A2(new_n760), .A3(new_n754), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n756), .A2(new_n636), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(G85gat), .B1(new_n764), .B2(new_n688), .ZN(new_n765));
  AOI211_X1 g564(.A(new_n729), .B(new_n755), .C1(new_n681), .C2(new_n686), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n441), .A2(new_n256), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(G1336gat));
  NOR2_X1   g567(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n513), .A2(G92gat), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n756), .A2(new_n636), .A3(new_n762), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n710), .A2(new_n636), .A3(new_n512), .A4(new_n754), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n769), .B(new_n773), .C1(new_n774), .C2(G92gat), .ZN(new_n775));
  INV_X1    g574(.A(new_n769), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(G92gat), .ZN(new_n777));
  INV_X1    g576(.A(new_n773), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n775), .A2(new_n779), .ZN(G1337gat));
  NAND3_X1  g579(.A1(new_n766), .A2(KEYINPUT117), .A3(new_n568), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n710), .A2(new_n636), .A3(new_n568), .A4(new_n754), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n781), .A2(new_n784), .A3(G99gat), .ZN(new_n785));
  OR3_X1    g584(.A1(new_n763), .A2(G99gat), .A3(new_n558), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(G1338gat));
  INV_X1    g586(.A(G106gat), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n372), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n710), .A2(new_n636), .A3(new_n754), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n763), .B2(new_n372), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(G1339gat));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n628), .A2(KEYINPUT54), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n625), .A2(new_n627), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n628), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n633), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n796), .A2(KEYINPUT55), .A3(new_n633), .A4(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n634), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n615), .B2(new_n617), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n604), .A2(new_n605), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n601), .B1(new_n597), .B2(new_n600), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n613), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n617), .A3(new_n636), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT118), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n809), .B(new_n812), .C1(new_n619), .C2(new_n803), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n278), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n808), .A2(new_n617), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n278), .A2(new_n803), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n243), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n243), .A2(new_n619), .A3(new_n729), .A4(new_n278), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n795), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n813), .A2(new_n278), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n816), .B1(new_n822), .B2(new_n811), .ZN(new_n823));
  OAI211_X1 g622(.A(KEYINPUT119), .B(new_n819), .C1(new_n823), .C2(new_n243), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n441), .A2(new_n512), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n821), .A2(new_n824), .A3(new_n559), .A4(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n619), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n821), .A2(new_n824), .A3(new_n668), .A4(new_n825), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n375), .A3(new_n618), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(G1340gat));
  OAI21_X1  g632(.A(G120gat), .B1(new_n826), .B2(new_n729), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n636), .A2(new_n377), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n834), .B1(new_n830), .B2(new_n835), .ZN(G1341gat));
  INV_X1    g635(.A(new_n243), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n826), .A2(new_n388), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n831), .A2(new_n243), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n388), .ZN(G1342gat));
  INV_X1    g639(.A(new_n385), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n830), .A2(new_n841), .A3(new_n278), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n826), .B2(new_n278), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n842), .A2(KEYINPUT121), .A3(new_n843), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT121), .B1(new_n842), .B2(new_n843), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(G1343gat));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n821), .A2(new_n824), .A3(new_n849), .A4(new_n723), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n278), .B1(new_n804), .B2(new_n810), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n243), .B1(new_n851), .B2(new_n817), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n819), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI211_X1 g653(.A(KEYINPUT122), .B(new_n243), .C1(new_n851), .C2(new_n817), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n723), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT57), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n568), .A2(new_n441), .A3(new_n512), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n850), .A2(new_n857), .A3(new_n618), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(G141gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n821), .A2(new_n824), .A3(new_n723), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n619), .A2(G141gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT58), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n860), .A2(new_n867), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n729), .A2(G148gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n862), .A2(new_n858), .A3(new_n870), .ZN(new_n871));
  XOR2_X1   g670(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n872));
  OAI21_X1  g671(.A(new_n849), .B1(new_n820), .B2(new_n852), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n372), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n874), .B1(new_n861), .B2(KEYINPUT57), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n636), .A3(new_n858), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n872), .B1(new_n876), .B2(G148gat), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n850), .A2(new_n857), .A3(new_n636), .A4(new_n858), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n878), .A2(new_n879), .A3(G148gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n871), .B1(new_n877), .B2(new_n880), .ZN(G1345gat));
  NAND3_X1  g680(.A1(new_n850), .A2(new_n857), .A3(new_n858), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(new_n289), .A3(new_n837), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n862), .A2(new_n243), .A3(new_n858), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n289), .B2(new_n884), .ZN(G1346gat));
  NOR3_X1   g684(.A1(new_n882), .A2(new_n294), .A3(new_n278), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n862), .A2(new_n277), .A3(new_n858), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n294), .B2(new_n887), .ZN(G1347gat));
  AND2_X1   g687(.A1(new_n821), .A2(new_n824), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n688), .A2(new_n513), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n559), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G169gat), .B1(new_n891), .B2(new_n619), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n821), .A2(new_n824), .ZN(new_n893));
  INV_X1    g692(.A(new_n668), .ZN(new_n894));
  INV_X1    g693(.A(new_n890), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n487), .A3(new_n618), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n892), .A2(new_n897), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n896), .B2(new_n636), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n893), .A2(new_n664), .A3(new_n895), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n636), .A2(new_n485), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(G1349gat));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n889), .A2(new_n668), .A3(new_n890), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n243), .A2(new_n478), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(G183gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n900), .B2(new_n243), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT60), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G183gat), .B1(new_n891), .B2(new_n837), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n243), .A3(new_n478), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n910), .A2(new_n903), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n909), .A2(new_n913), .ZN(G1350gat));
  NAND2_X1  g713(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n915));
  OAI211_X1 g714(.A(G190gat), .B(new_n915), .C1(new_n891), .C2(new_n278), .ZN(new_n916));
  NOR2_X1   g715(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n479), .B1(new_n900), .B2(new_n277), .ZN(new_n919));
  INV_X1    g718(.A(new_n917), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n896), .A2(new_n479), .A3(new_n277), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(G1351gat));
  NAND2_X1  g722(.A1(new_n861), .A2(KEYINPUT57), .ZN(new_n924));
  INV_X1    g723(.A(new_n874), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n895), .A2(new_n568), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n924), .A2(new_n618), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT126), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n875), .A2(new_n929), .A3(new_n618), .A4(new_n926), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(G197gat), .A3(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n861), .A2(new_n568), .A3(new_n895), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n304), .A3(new_n618), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1352gat));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n305), .A3(new_n636), .ZN(new_n935));
  XOR2_X1   g734(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n932), .A2(new_n305), .A3(new_n636), .A4(new_n936), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n875), .A2(new_n636), .A3(new_n926), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n938), .B(new_n939), .C1(new_n305), .C2(new_n940), .ZN(G1353gat));
  NAND2_X1  g740(.A1(new_n862), .A2(new_n926), .ZN(new_n942));
  OR3_X1    g741(.A1(new_n942), .A2(G211gat), .A3(new_n837), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n924), .A2(new_n243), .A3(new_n925), .A4(new_n926), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n944), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT63), .B1(new_n944), .B2(G211gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G1354gat));
  NAND3_X1  g746(.A1(new_n875), .A2(new_n277), .A3(new_n926), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G218gat), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n278), .A2(G218gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n942), .B2(new_n950), .ZN(G1355gat));
endmodule


