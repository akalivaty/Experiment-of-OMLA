//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G119), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT68), .A3(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT2), .B(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G113), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT2), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G113), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n205), .A2(new_n194), .A3(new_n196), .A4(new_n197), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n200), .A2(new_n206), .A3(KEYINPUT69), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT69), .B1(new_n200), .B2(new_n206), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G134), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G137), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT11), .ZN(new_n218));
  OAI22_X1  g032(.A1(new_n217), .A2(new_n218), .B1(new_n212), .B2(G134), .ZN(new_n219));
  OAI22_X1  g033(.A1(new_n214), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n217), .A2(new_n218), .A3(new_n212), .A4(G134), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n216), .B1(new_n222), .B2(new_n211), .ZN(new_n223));
  XNOR2_X1  g037(.A(G143), .B(G146), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G128), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT67), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n227), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n236));
  INV_X1    g050(.A(G143), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(G146), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(KEYINPUT65), .A3(G143), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(G146), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n226), .B1(new_n235), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n223), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n244), .A2(new_n247), .B1(new_n245), .B2(new_n224), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n221), .A2(new_n220), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n214), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n249), .A2(new_n211), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n211), .B1(new_n249), .B2(new_n250), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n243), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT30), .B1(new_n254), .B2(KEYINPUT64), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT64), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT30), .ZN(new_n257));
  AOI211_X1 g071(.A(new_n256), .B(new_n257), .C1(new_n243), .C2(new_n253), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n210), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n200), .A2(new_n206), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n207), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n253), .A3(new_n243), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n191), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n254), .A2(new_n210), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(new_n264), .ZN(new_n268));
  INV_X1    g082(.A(new_n191), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n249), .A2(new_n250), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G131), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n222), .A2(new_n211), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n273), .A2(new_n248), .B1(new_n242), .B2(new_n223), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT28), .B1(new_n274), .B2(new_n263), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n268), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n265), .A2(new_n276), .A3(KEYINPUT29), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(KEYINPUT29), .ZN(new_n278));
  INV_X1    g092(.A(G902), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(G472), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n257), .B1(new_n274), .B2(new_n256), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n254), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n263), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n264), .A2(new_n191), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT31), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT31), .ZN(new_n287));
  INV_X1    g101(.A(new_n285), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n259), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n269), .B1(new_n268), .B2(new_n275), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n286), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  NOR2_X1   g106(.A1(G472), .A2(G902), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n281), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n281), .B(KEYINPUT70), .C1(new_n294), .C2(new_n295), .ZN(new_n299));
  XNOR2_X1  g113(.A(G125), .B(G140), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT16), .ZN(new_n301));
  INV_X1    g115(.A(G125), .ZN(new_n302));
  OR3_X1    g116(.A1(new_n302), .A2(KEYINPUT16), .A3(G140), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(G146), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n300), .A2(new_n233), .ZN(new_n305));
  XOR2_X1   g119(.A(KEYINPUT24), .B(G110), .Z(new_n306));
  NAND2_X1  g120(.A1(new_n195), .A2(G128), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n227), .A2(G119), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT71), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n307), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n306), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n195), .B2(G128), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n227), .A2(KEYINPUT23), .A3(G119), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(new_n307), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(G110), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n304), .B(new_n305), .C1(new_n313), .C2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n310), .A2(new_n312), .A3(new_n306), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n301), .A2(G146), .A3(new_n303), .ZN(new_n321));
  AOI21_X1  g135(.A(G146), .B1(new_n301), .B2(new_n303), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n317), .A2(new_n324), .ZN(new_n326));
  INV_X1    g140(.A(G110), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n319), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g145(.A(KEYINPUT73), .B(new_n319), .C1(new_n323), .C2(new_n328), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G137), .ZN(new_n333));
  INV_X1    g147(.A(G953), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(G221), .A3(G234), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(KEYINPUT74), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n331), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n319), .B(new_n336), .C1(new_n323), .C2(new_n328), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n340));
  AOI21_X1  g154(.A(G902), .B1(new_n340), .B2(KEYINPUT75), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n340), .A2(KEYINPUT75), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G217), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(G234), .B2(new_n279), .ZN(new_n346));
  INV_X1    g160(.A(new_n343), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n338), .A2(new_n339), .A3(new_n347), .A4(new_n341), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n338), .A2(new_n339), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n346), .A2(G902), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT76), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n346), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n342), .B2(new_n343), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n359), .A2(new_n348), .B1(new_n351), .B2(new_n353), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT77), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n298), .A2(new_n299), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT90), .ZN(new_n364));
  XNOR2_X1  g178(.A(G110), .B(G140), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n334), .A2(G227), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n273), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n242), .A2(KEYINPUT10), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n370));
  INV_X1    g184(.A(G107), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G104), .ZN(new_n372));
  AND2_X1   g186(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n373));
  NOR2_X1   g187(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G101), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(G104), .A3(new_n371), .ZN(new_n378));
  INV_X1    g192(.A(G104), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G107), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n375), .A2(new_n376), .A3(new_n378), .A4(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT79), .B1(new_n371), .B2(G104), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n379), .A3(G107), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n384), .A3(new_n372), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G101), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n369), .A2(new_n370), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  INV_X1    g203(.A(new_n234), .ZN(new_n390));
  OAI21_X1  g204(.A(G128), .B1(new_n225), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n244), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n389), .B1(new_n392), .B2(new_n226), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n381), .A2(new_n386), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT81), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  INV_X1    g211(.A(new_n375), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n378), .A2(new_n380), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n397), .B(G101), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n381), .A2(KEYINPUT4), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n371), .A2(G104), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n379), .A2(G107), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n377), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n376), .B1(new_n404), .B2(new_n375), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n248), .B(new_n400), .C1(new_n401), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n234), .A2(new_n240), .A3(G128), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT80), .B1(new_n408), .B2(new_n232), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n234), .A2(new_n240), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n233), .A2(G143), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n410), .A2(new_n227), .B1(KEYINPUT1), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n224), .A2(new_n225), .A3(new_n413), .A4(G128), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT10), .B1(new_n394), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n407), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n368), .B1(new_n396), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n370), .B1(new_n369), .B2(new_n387), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n393), .A2(KEYINPUT81), .A3(new_n394), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n409), .A2(new_n412), .A3(new_n414), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n389), .B1(new_n422), .B2(new_n387), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n406), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n421), .A2(new_n424), .A3(new_n273), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n367), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n417), .A2(new_n368), .A3(new_n419), .A4(new_n420), .ZN(new_n427));
  INV_X1    g241(.A(new_n367), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n394), .B2(new_n242), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n394), .A2(new_n415), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n234), .A2(new_n240), .A3(G128), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n391), .A2(new_n244), .B1(new_n225), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT82), .A3(new_n387), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n430), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n435), .A2(KEYINPUT12), .A3(new_n273), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT12), .B1(new_n435), .B2(new_n273), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n427), .B(new_n428), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n426), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G469), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n279), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(new_n279), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n273), .B1(new_n421), .B2(new_n424), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n427), .A2(new_n444), .A3(new_n428), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n435), .A2(new_n273), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT12), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n435), .A2(KEYINPUT12), .A3(new_n273), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n421), .A2(new_n424), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n448), .A2(new_n449), .B1(new_n450), .B2(new_n368), .ZN(new_n451));
  OAI211_X1 g265(.A(G469), .B(new_n445), .C1(new_n451), .C2(new_n428), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n441), .A2(new_n443), .A3(new_n452), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n454));
  AOI21_X1  g268(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n455));
  OAI21_X1  g269(.A(G131), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n187), .A2(G214), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n237), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(KEYINPUT86), .A3(G131), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT17), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n301), .A2(new_n303), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n233), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n304), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT17), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n454), .A2(new_n455), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n211), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n458), .A2(new_n463), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n465), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(G113), .B(G122), .Z(new_n475));
  XOR2_X1   g289(.A(KEYINPUT87), .B(G104), .Z(new_n476));
  XOR2_X1   g290(.A(new_n475), .B(new_n476), .Z(new_n477));
  INV_X1    g291(.A(KEYINPUT18), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n471), .B1(new_n478), .B2(new_n211), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n462), .A2(KEYINPUT18), .A3(G131), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n300), .B(new_n233), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n474), .A2(new_n477), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n477), .B1(new_n474), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n279), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT88), .B(G475), .Z(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G478), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT9), .B(G234), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n491), .A2(new_n345), .A3(G953), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n237), .A2(G128), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n227), .A2(G143), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n214), .ZN(new_n496));
  XNOR2_X1  g310(.A(G116), .B(G122), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n371), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n193), .A2(KEYINPUT14), .A3(G122), .ZN(new_n499));
  INV_X1    g313(.A(new_n497), .ZN(new_n500));
  OAI211_X1 g314(.A(G107), .B(new_n499), .C1(new_n500), .C2(KEYINPUT14), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n493), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n503), .A2(KEYINPUT13), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n494), .B1(new_n503), .B2(KEYINPUT13), .ZN(new_n505));
  OAI21_X1  g319(.A(G134), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n495), .A2(new_n214), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n497), .B(new_n371), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n492), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n502), .A2(new_n509), .A3(new_n492), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n490), .B1(new_n513), .B2(new_n279), .ZN(new_n514));
  INV_X1    g328(.A(new_n512), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n279), .B(new_n490), .C1(new_n515), .C2(new_n510), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT20), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n458), .A2(new_n463), .A3(new_n472), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n300), .B(KEYINPUT19), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n233), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n304), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n477), .B1(new_n523), .B2(new_n482), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n474), .A2(new_n477), .A3(new_n482), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(G475), .A2(G902), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n519), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n528), .ZN(new_n530));
  AOI211_X1 g344(.A(KEYINPUT20), .B(new_n530), .C1(new_n525), .C2(new_n526), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n487), .B(new_n518), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n334), .A2(G952), .ZN(new_n533));
  INV_X1    g347(.A(G234), .ZN(new_n534));
  INV_X1    g348(.A(G237), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(G902), .B(G953), .C1(new_n534), .C2(new_n535), .ZN(new_n538));
  XOR2_X1   g352(.A(new_n538), .B(KEYINPUT89), .Z(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT21), .B(G898), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G221), .B1(new_n491), .B2(G902), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n453), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G210), .B1(G237), .B2(G902), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n193), .A2(G119), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT5), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n201), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n198), .B2(new_n548), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n394), .A2(new_n206), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n400), .B1(new_n401), .B2(new_n405), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n263), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT6), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G122), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT83), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n433), .A2(new_n302), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n248), .A2(new_n302), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G224), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(G953), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n564), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n561), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n551), .B(new_n555), .C1(new_n263), .C2(new_n552), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT6), .ZN(new_n570));
  OAI21_X1  g384(.A(G101), .B1(new_n398), .B2(new_n399), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(KEYINPUT4), .A3(new_n381), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n572), .A2(new_n262), .A3(new_n207), .A4(new_n400), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n557), .B1(new_n573), .B2(new_n551), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n559), .B(new_n568), .C1(new_n570), .C2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n555), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n550), .A2(new_n206), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n578), .A2(new_n387), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n387), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT84), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n564), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n562), .A2(new_n584), .B1(KEYINPUT7), .B2(new_n566), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n566), .A2(KEYINPUT7), .ZN(new_n586));
  AOI211_X1 g400(.A(new_n583), .B(new_n586), .C1(new_n560), .C2(new_n561), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n569), .B(new_n581), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n279), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n546), .B1(new_n576), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT85), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n562), .A2(new_n584), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n586), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n562), .A2(new_n582), .A3(KEYINPUT7), .A4(new_n566), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n569), .A2(new_n581), .ZN(new_n596));
  AOI21_X1  g410(.A(G902), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n575), .A3(new_n545), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n590), .A2(new_n591), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(G214), .B1(G237), .B2(G902), .ZN(new_n600));
  OAI211_X1 g414(.A(KEYINPUT85), .B(new_n546), .C1(new_n576), .C2(new_n589), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n364), .B1(new_n544), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n543), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n452), .A2(new_n443), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n604), .B1(new_n606), .B2(new_n441), .ZN(new_n607));
  INV_X1    g421(.A(new_n602), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT90), .A4(new_n542), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n363), .A2(new_n603), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT91), .B(G101), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G3));
  INV_X1    g426(.A(new_n541), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n590), .A2(KEYINPUT92), .A3(new_n598), .ZN(new_n614));
  INV_X1    g428(.A(new_n600), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n545), .B1(new_n597), .B2(new_n575), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT92), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT93), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n614), .A2(new_n618), .A3(KEYINPUT93), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n513), .A2(new_n488), .A3(new_n279), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n488), .B2(new_n279), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n513), .B(KEYINPUT33), .Z(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(G478), .ZN(new_n626));
  INV_X1    g440(.A(new_n482), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n468), .B1(KEYINPUT17), .B2(new_n464), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n627), .B1(new_n628), .B2(new_n473), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n524), .B1(new_n629), .B2(new_n477), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT20), .B1(new_n630), .B2(new_n530), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n527), .A2(new_n519), .A3(new_n528), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n487), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  AND4_X1   g449(.A1(new_n613), .A2(new_n621), .A3(new_n622), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n291), .A2(new_n279), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n637), .A2(G472), .B1(new_n291), .B2(new_n293), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n357), .A3(new_n361), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n453), .A2(new_n543), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  AND3_X1   g458(.A1(new_n614), .A2(new_n618), .A3(KEYINPUT93), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT93), .B1(new_n614), .B2(new_n618), .ZN(new_n646));
  INV_X1    g460(.A(new_n518), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n633), .A2(new_n647), .A3(new_n487), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n648), .A2(new_n541), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n645), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n641), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT94), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NAND2_X1  g468(.A1(new_n637), .A2(G472), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n291), .A2(new_n293), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n337), .A2(KEYINPUT36), .ZN(new_n658));
  INV_X1    g472(.A(new_n331), .ZN(new_n659));
  INV_X1    g473(.A(new_n332), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n331), .B(new_n332), .C1(KEYINPUT36), .C2(new_n337), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n353), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n349), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n657), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n609), .A2(new_n603), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT37), .B(G110), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G12));
  AND3_X1   g484(.A1(new_n298), .A2(new_n299), .A3(new_n665), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n645), .A2(new_n640), .A3(new_n646), .ZN(new_n672));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n539), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n536), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n648), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n671), .A2(new_n672), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  NAND2_X1  g493(.A1(new_n599), .A2(new_n601), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT96), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n675), .B(KEYINPUT39), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n607), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n683), .B1(KEYINPUT40), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n259), .A2(new_n264), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n191), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n267), .A2(new_n264), .A3(new_n269), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT97), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n689), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n687), .B2(new_n191), .ZN(new_n694));
  AOI21_X1  g508(.A(G902), .B1(new_n694), .B2(KEYINPUT97), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G472), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n656), .A2(KEYINPUT32), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n665), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n634), .A2(new_n647), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n701), .A2(new_n600), .A3(new_n703), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n686), .B(new_n704), .C1(KEYINPUT40), .C2(new_n685), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT98), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n237), .ZN(G45));
  AND3_X1   g521(.A1(new_n626), .A2(new_n634), .A3(new_n675), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n298), .A2(new_n299), .A3(new_n665), .A4(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n645), .A2(new_n646), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n607), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT99), .B(G146), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G48));
  NOR2_X1   g528(.A1(new_n425), .A2(new_n367), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n448), .A2(new_n449), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n427), .A2(new_n444), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n715), .A2(new_n716), .B1(new_n717), .B2(new_n367), .ZN(new_n718));
  OAI21_X1  g532(.A(G469), .B1(new_n718), .B2(G902), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n543), .A3(new_n441), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT100), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n719), .A2(KEYINPUT100), .A3(new_n543), .A4(new_n441), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n363), .A2(new_n636), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT41), .B(G113), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G15));
  AOI21_X1  g541(.A(KEYINPUT70), .B1(new_n700), .B2(new_n281), .ZN(new_n728));
  INV_X1    g542(.A(new_n299), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n362), .A3(new_n650), .A4(new_n724), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT101), .B(G116), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G18));
  AND4_X1   g547(.A1(new_n298), .A2(new_n299), .A3(new_n542), .A4(new_n665), .ZN(new_n734));
  AND4_X1   g548(.A1(new_n621), .A2(new_n722), .A3(new_n622), .A4(new_n723), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  OAI21_X1  g551(.A(KEYINPUT102), .B1(new_n657), .B2(new_n355), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT102), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n638), .A2(new_n739), .A3(new_n360), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n645), .A2(new_n646), .A3(new_n702), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n724), .A3(new_n613), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  NAND4_X1  g558(.A1(new_n724), .A2(new_n710), .A3(new_n667), .A4(new_n708), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  NOR2_X1   g560(.A1(new_n604), .A2(new_n615), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n599), .B2(new_n601), .ZN(new_n749));
  AOI211_X1 g563(.A(G469), .B(G902), .C1(new_n426), .C2(new_n438), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT103), .B1(new_n605), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT103), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n441), .A2(new_n752), .A3(new_n443), .A4(new_n452), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n749), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n298), .A2(new_n299), .A3(new_n362), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n708), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(KEYINPUT42), .ZN(new_n759));
  AND4_X1   g573(.A1(new_n708), .A2(new_n749), .A3(new_n751), .A4(new_n753), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT104), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n296), .A2(new_n761), .A3(new_n360), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n761), .B1(new_n296), .B2(new_n360), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n757), .A2(new_n759), .B1(new_n764), .B2(KEYINPUT42), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n754), .A2(new_n298), .A3(new_n299), .A4(new_n362), .ZN(new_n768));
  INV_X1    g582(.A(new_n677), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n363), .A2(KEYINPUT105), .A3(new_n677), .A4(new_n754), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NAND2_X1  g587(.A1(new_n680), .A2(new_n600), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT107), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n634), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n626), .A2(new_n633), .A3(new_n487), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n777), .B(new_n778), .Z(new_n779));
  OAI21_X1  g593(.A(KEYINPUT108), .B1(new_n638), .B2(new_n666), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n638), .A2(new_n666), .A3(KEYINPUT108), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n774), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n445), .B1(new_n451), .B2(new_n428), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n440), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT106), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n787), .B2(new_n786), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n788), .A2(KEYINPUT106), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n443), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT46), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n750), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n604), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n684), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n785), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  XNOR2_X1  g613(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT47), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n796), .B1(KEYINPUT109), .B2(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n730), .A2(new_n362), .A3(new_n758), .A4(new_n774), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n676), .A2(new_n604), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n294), .A2(new_n295), .ZN(new_n809));
  INV_X1    g623(.A(G472), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n692), .B2(new_n695), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n666), .B(new_n808), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n751), .A2(new_n753), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n807), .B1(new_n814), .B2(new_n742), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n621), .A2(new_n622), .A3(new_n703), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n816), .A2(new_n812), .A3(KEYINPUT114), .A4(new_n813), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n730), .A2(new_n665), .A3(new_n672), .A4(new_n708), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n678), .A2(new_n819), .A3(new_n745), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT52), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n710), .A2(new_n722), .A3(new_n723), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n667), .A2(new_n708), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n298), .A2(new_n677), .A3(new_n299), .A4(new_n665), .ZN(new_n824));
  OAI22_X1  g638(.A1(new_n822), .A2(new_n823), .B1(new_n824), .B2(new_n711), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n712), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n751), .A2(new_n753), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n701), .A2(new_n827), .A3(new_n808), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT114), .B1(new_n828), .B2(new_n816), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n814), .A2(new_n807), .A3(new_n742), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n826), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n821), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n755), .A2(new_n823), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n532), .A2(new_n676), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT112), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n838), .A2(new_n640), .A3(new_n774), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n836), .B1(new_n671), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n772), .A2(new_n765), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n641), .A2(new_n608), .A3(new_n613), .A4(new_n635), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n648), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n633), .A2(new_n647), .A3(KEYINPUT110), .A4(new_n487), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT111), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n608), .A3(new_n847), .A4(new_n613), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n845), .A3(new_n613), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT111), .B1(new_n849), .B2(new_n602), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n641), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n610), .A2(new_n668), .A3(new_n842), .A4(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n725), .A2(new_n736), .A3(new_n731), .A4(new_n743), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n841), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT53), .B1(new_n835), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(KEYINPUT115), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n722), .A2(new_n723), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n756), .A2(new_n857), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n858), .A2(new_n650), .B1(new_n734), .B2(new_n735), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n725), .A4(new_n743), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n609), .A2(new_n603), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n842), .B1(new_n862), .B2(new_n756), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n851), .A2(new_n668), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n856), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n834), .A2(new_n867), .A3(new_n841), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n855), .A2(new_n868), .A3(KEYINPUT116), .A4(KEYINPUT54), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n835), .B(new_n854), .C1(KEYINPUT113), .C2(KEYINPUT53), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n772), .A2(new_n765), .A3(new_n840), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n853), .A2(new_n852), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n821), .A3(new_n833), .A4(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT113), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n873), .B(new_n865), .C1(new_n874), .C2(new_n834), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT54), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n867), .A2(new_n841), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n879), .A2(new_n835), .B1(new_n873), .B2(new_n865), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n869), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n857), .A2(new_n774), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n697), .A2(new_n700), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AND4_X1   g700(.A1(new_n362), .A2(new_n884), .A3(new_n537), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n635), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n779), .A2(new_n537), .A3(new_n741), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n735), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n533), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT119), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT48), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n884), .A2(new_n537), .A3(new_n779), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n762), .A2(new_n763), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n897), .B2(new_n896), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n888), .A2(new_n900), .A3(new_n533), .A4(new_n890), .ZN(new_n901));
  OAI211_X1 g715(.A(KEYINPUT120), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n892), .A2(new_n899), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT121), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n894), .A2(new_n657), .A3(new_n666), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT118), .Z(new_n906));
  NAND4_X1  g720(.A1(new_n889), .A2(new_n615), .A3(new_n683), .A4(new_n724), .ZN(new_n907));
  OR3_X1    g721(.A1(new_n907), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n908));
  XOR2_X1   g722(.A(KEYINPUT117), .B(KEYINPUT50), .Z(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n626), .A2(new_n634), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n887), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n906), .A2(new_n908), .A3(new_n910), .A4(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n719), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n750), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n801), .A2(new_n803), .B1(new_n604), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n889), .A2(new_n600), .A3(new_n680), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT51), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n914), .A2(new_n919), .A3(KEYINPUT51), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n904), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI22_X1  g738(.A1(new_n883), .A2(new_n924), .B1(G952), .B2(G953), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n916), .B(KEYINPUT49), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n778), .A2(new_n355), .A3(new_n748), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n926), .A2(new_n683), .A3(new_n886), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n925), .A2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n334), .A2(G952), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n559), .B1(new_n570), .B2(new_n574), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(new_n568), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n879), .A2(new_n835), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n873), .A2(new_n865), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(G210), .A3(G902), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT122), .B1(new_n880), .B2(new_n279), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n942), .B(G902), .C1(new_n855), .C2(new_n868), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n546), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n933), .A2(KEYINPUT56), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n930), .B(new_n940), .C1(new_n944), .C2(new_n945), .ZN(G51));
  XNOR2_X1  g760(.A(new_n880), .B(KEYINPUT54), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n442), .B(KEYINPUT57), .Z(new_n948));
  OAI21_X1  g762(.A(new_n439), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n790), .A2(new_n791), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n941), .A2(new_n950), .A3(new_n943), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n930), .B1(new_n949), .B2(new_n951), .ZN(G54));
  AND2_X1   g766(.A1(KEYINPUT58), .A2(G475), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n941), .A2(new_n943), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(new_n630), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n954), .B2(new_n630), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n941), .A2(new_n943), .A3(new_n527), .A4(new_n953), .ZN(new_n958));
  INV_X1    g772(.A(new_n930), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n956), .A2(new_n957), .A3(new_n960), .ZN(G60));
  XOR2_X1   g775(.A(new_n625), .B(KEYINPUT124), .Z(new_n962));
  NOR2_X1   g776(.A1(new_n488), .A2(new_n279), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT59), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n959), .B1(new_n947), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n964), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n883), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n966), .B1(new_n968), .B2(new_n962), .ZN(G63));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT60), .Z(new_n971));
  NAND2_X1  g785(.A1(new_n937), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n350), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n937), .A2(new_n663), .A3(new_n971), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n959), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G66));
  OAI21_X1  g791(.A(G953), .B1(new_n540), .B2(new_n563), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n872), .B2(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n931), .B1(G898), .B2(new_n334), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT125), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n979), .B(new_n981), .ZN(G69));
  AOI21_X1  g796(.A(new_n334), .B1(G227), .B2(G900), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n282), .A2(new_n283), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(new_n521), .ZN(new_n985));
  OR3_X1    g799(.A1(new_n797), .A2(new_n816), .A3(new_n895), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n986), .A2(new_n765), .A3(new_n772), .A4(new_n826), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n805), .A2(new_n798), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n334), .B(new_n985), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n846), .A2(new_n635), .ZN(new_n990));
  NOR4_X1   g804(.A1(new_n756), .A2(new_n990), .A3(new_n685), .A4(new_n774), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n992));
  OR3_X1    g806(.A1(new_n706), .A2(new_n992), .A3(new_n820), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n706), .B2(new_n820), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n988), .ZN(new_n996));
  AOI21_X1  g810(.A(G953), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n989), .B1(new_n997), .B2(new_n985), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n983), .B1(new_n998), .B2(new_n673), .ZN(new_n999));
  INV_X1    g813(.A(new_n983), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n989), .B(new_n1000), .C1(new_n997), .C2(new_n985), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(G72));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT63), .Z(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT126), .Z(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n987), .A2(new_n988), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1006), .B1(new_n1007), .B2(new_n872), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n259), .A2(new_n264), .A3(new_n269), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT127), .Z(new_n1010));
  OAI21_X1  g824(.A(new_n959), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n995), .A2(new_n872), .A3(new_n996), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n688), .B1(new_n1012), .B2(new_n1005), .ZN(new_n1013));
  AND4_X1   g827(.A1(new_n688), .A2(new_n876), .A3(new_n1009), .A4(new_n1004), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(G57));
endmodule


