

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792;

  NOR2_X1 U386 ( .A1(n608), .A2(n450), .ZN(n616) );
  NAND2_X2 U387 ( .A1(n416), .A2(n412), .ZN(n592) );
  AND2_X1 U388 ( .A1(n661), .A2(n472), .ZN(n364) );
  INV_X2 U389 ( .A(G143), .ZN(n476) );
  XNOR2_X1 U390 ( .A(n453), .B(KEYINPUT76), .ZN(n636) );
  NOR2_X1 U391 ( .A1(n708), .A2(n709), .ZN(n453) );
  XNOR2_X2 U392 ( .A(n509), .B(n475), .ZN(n524) );
  XNOR2_X2 U393 ( .A(n476), .B(G128), .ZN(n509) );
  INV_X1 U394 ( .A(n696), .ZN(n693) );
  INV_X1 U395 ( .A(G116), .ZN(n459) );
  AND2_X1 U396 ( .A1(n391), .A2(n389), .ZN(n388) );
  BUF_X1 U397 ( .A(n751), .Z(n365) );
  OR2_X1 U398 ( .A1(n704), .A2(n429), .ZN(n432) );
  XNOR2_X1 U399 ( .A(n588), .B(n587), .ZN(n620) );
  NAND2_X1 U400 ( .A1(n409), .A2(n408), .ZN(n609) );
  XNOR2_X1 U401 ( .A(n527), .B(n528), .ZN(n614) );
  XNOR2_X1 U402 ( .A(n551), .B(n550), .ZN(n645) );
  XNOR2_X1 U403 ( .A(n513), .B(n512), .ZN(n670) );
  XNOR2_X1 U404 ( .A(n764), .B(n421), .ZN(n513) );
  XNOR2_X1 U405 ( .A(n461), .B(KEYINPUT3), .ZN(n460) );
  XNOR2_X1 U406 ( .A(n486), .B(n435), .ZN(n539) );
  XNOR2_X1 U407 ( .A(n459), .B(G113), .ZN(n458) );
  XNOR2_X1 U408 ( .A(G146), .B(G125), .ZN(n503) );
  BUF_X1 U409 ( .A(n630), .Z(n366) );
  XNOR2_X2 U410 ( .A(n452), .B(G110), .ZN(n763) );
  XNOR2_X2 U411 ( .A(G107), .B(G104), .ZN(n452) );
  XNOR2_X2 U412 ( .A(n451), .B(n557), .ZN(n421) );
  XNOR2_X1 U413 ( .A(n503), .B(KEYINPUT10), .ZN(n537) );
  NAND2_X1 U414 ( .A1(G214), .A2(n564), .ZN(n722) );
  AND2_X1 U415 ( .A1(n657), .A2(n404), .ZN(n403) );
  OR2_X1 U416 ( .A1(n746), .A2(n413), .ZN(n412) );
  NAND2_X1 U417 ( .A1(n415), .A2(n414), .ZN(n413) );
  INV_X1 U418 ( .A(G902), .ZN(n414) );
  NOR2_X1 U419 ( .A1(G902), .A2(n748), .ZN(n488) );
  NOR2_X1 U420 ( .A1(n744), .A2(G902), .ZN(n527) );
  NAND2_X1 U421 ( .A1(G221), .A2(n539), .ZN(n547) );
  INV_X1 U422 ( .A(KEYINPUT64), .ZN(n431) );
  NAND2_X1 U423 ( .A1(n751), .A2(G475), .ZN(n425) );
  INV_X1 U424 ( .A(KEYINPUT94), .ZN(n500) );
  INV_X1 U425 ( .A(KEYINPUT67), .ZN(n472) );
  INV_X1 U426 ( .A(KEYINPUT38), .ZN(n380) );
  INV_X1 U427 ( .A(n572), .ZN(n440) );
  INV_X1 U428 ( .A(n722), .ZN(n428) );
  OR2_X1 U429 ( .A1(n645), .A2(n648), .ZN(n709) );
  XNOR2_X1 U430 ( .A(G140), .B(KEYINPUT98), .ZN(n542) );
  XNOR2_X1 U431 ( .A(G137), .B(G119), .ZN(n540) );
  XNOR2_X1 U432 ( .A(G110), .B(KEYINPUT99), .ZN(n536) );
  XNOR2_X1 U433 ( .A(n420), .B(KEYINPUT7), .ZN(n484) );
  XNOR2_X1 U434 ( .A(G122), .B(KEYINPUT9), .ZN(n420) );
  XNOR2_X1 U435 ( .A(G116), .B(G107), .ZN(n487) );
  INV_X1 U436 ( .A(G134), .ZN(n475) );
  INV_X1 U437 ( .A(KEYINPUT8), .ZN(n435) );
  XNOR2_X1 U438 ( .A(G143), .B(G104), .ZN(n494) );
  INV_X1 U439 ( .A(KEYINPUT86), .ZN(n445) );
  AND2_X1 U440 ( .A1(n401), .A2(n398), .ZN(n397) );
  NAND2_X1 U441 ( .A1(n400), .A2(n399), .ZN(n398) );
  OR2_X1 U442 ( .A1(n403), .A2(KEYINPUT36), .ZN(n401) );
  NAND2_X1 U443 ( .A1(n395), .A2(n403), .ZN(n394) );
  NOR2_X1 U444 ( .A1(n402), .A2(n399), .ZN(n396) );
  INV_X1 U445 ( .A(n481), .ZN(n402) );
  NAND2_X1 U446 ( .A1(n442), .A2(n441), .ZN(n634) );
  OR2_X1 U447 ( .A1(n437), .A2(n711), .ZN(n646) );
  XNOR2_X1 U448 ( .A(n427), .B(n426), .ZN(n575) );
  INV_X1 U449 ( .A(KEYINPUT28), .ZN(n426) );
  AND2_X1 U450 ( .A1(n411), .A2(n410), .ZN(n409) );
  XNOR2_X1 U451 ( .A(n611), .B(KEYINPUT6), .ZN(n657) );
  AND2_X2 U452 ( .A1(n383), .A2(n669), .ZN(n751) );
  XNOR2_X1 U453 ( .A(n526), .B(n525), .ZN(n744) );
  XNOR2_X1 U454 ( .A(n522), .B(n369), .ZN(n523) );
  INV_X1 U455 ( .A(KEYINPUT17), .ZN(n505) );
  NAND2_X1 U456 ( .A1(n463), .A2(n462), .ZN(n461) );
  INV_X1 U457 ( .A(G119), .ZN(n499) );
  XNOR2_X1 U458 ( .A(n614), .B(KEYINPUT1), .ZN(n708) );
  NOR2_X1 U459 ( .A1(G953), .A2(G237), .ZN(n558) );
  XNOR2_X1 U460 ( .A(KEYINPUT4), .B(KEYINPUT66), .ZN(n775) );
  XNOR2_X1 U461 ( .A(G113), .B(G122), .ZN(n489) );
  XOR2_X1 U462 ( .A(KEYINPUT103), .B(KEYINPUT105), .Z(n490) );
  XNOR2_X1 U463 ( .A(n448), .B(n493), .ZN(n495) );
  XOR2_X1 U464 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n493) );
  XNOR2_X1 U465 ( .A(n492), .B(n449), .ZN(n448) );
  INV_X1 U466 ( .A(KEYINPUT104), .ZN(n449) );
  NAND2_X1 U467 ( .A1(n471), .A2(n470), .ZN(n467) );
  NOR2_X1 U468 ( .A1(n660), .A2(n472), .ZN(n470) );
  XNOR2_X1 U469 ( .A(n524), .B(G137), .ZN(n772) );
  XNOR2_X1 U470 ( .A(n775), .B(G101), .ZN(n557) );
  INV_X1 U471 ( .A(KEYINPUT36), .ZN(n399) );
  INV_X1 U472 ( .A(KEYINPUT33), .ZN(n473) );
  NAND2_X1 U473 ( .A1(n657), .A2(n636), .ZN(n474) );
  NOR2_X1 U474 ( .A1(G902), .A2(G237), .ZN(n514) );
  NOR2_X1 U475 ( .A1(n407), .A2(n406), .ZN(n405) );
  AND2_X1 U476 ( .A1(n418), .A2(n417), .ZN(n416) );
  XNOR2_X1 U477 ( .A(n501), .B(G122), .ZN(n502) );
  XOR2_X1 U478 ( .A(KEYINPUT75), .B(KEYINPUT16), .Z(n501) );
  XNOR2_X1 U479 ( .A(KEYINPUT15), .B(G902), .ZN(n668) );
  NOR2_X1 U480 ( .A1(n664), .A2(KEYINPUT2), .ZN(n665) );
  XNOR2_X1 U481 ( .A(n772), .B(G146), .ZN(n555) );
  XNOR2_X1 U482 ( .A(n763), .B(KEYINPUT72), .ZN(n451) );
  NAND2_X1 U483 ( .A1(KEYINPUT2), .A2(KEYINPUT86), .ZN(n429) );
  NOR2_X1 U484 ( .A1(n726), .A2(n725), .ZN(n594) );
  AND2_X1 U485 ( .A1(n640), .A2(n440), .ZN(n439) );
  INV_X1 U486 ( .A(KEYINPUT30), .ZN(n565) );
  NAND2_X1 U487 ( .A1(n751), .A2(G472), .ZN(n678) );
  XNOR2_X1 U488 ( .A(n548), .B(n549), .ZN(n750) );
  XNOR2_X1 U489 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U490 ( .A(n483), .B(n482), .ZN(n748) );
  XNOR2_X1 U491 ( .A(n524), .B(n433), .ZN(n483) );
  XNOR2_X1 U492 ( .A(n484), .B(n487), .ZN(n433) );
  NAND2_X1 U493 ( .A1(n751), .A2(G210), .ZN(n478) );
  INV_X1 U494 ( .A(n381), .ZN(n702) );
  XNOR2_X1 U495 ( .A(n590), .B(n589), .ZN(n791) );
  INV_X1 U496 ( .A(KEYINPUT40), .ZN(n589) );
  XNOR2_X1 U497 ( .A(n447), .B(n446), .ZN(n789) );
  INV_X1 U498 ( .A(KEYINPUT112), .ZN(n446) );
  NAND2_X1 U499 ( .A1(n397), .A2(n394), .ZN(n480) );
  NAND2_X1 U500 ( .A1(n455), .A2(n635), .ZN(n454) );
  XNOR2_X1 U501 ( .A(n634), .B(n633), .ZN(n455) );
  XNOR2_X1 U502 ( .A(n465), .B(KEYINPUT32), .ZN(n464) );
  INV_X1 U503 ( .A(KEYINPUT68), .ZN(n465) );
  XNOR2_X1 U504 ( .A(n576), .B(KEYINPUT83), .ZN(n694) );
  INV_X1 U505 ( .A(n694), .ZN(n688) );
  XNOR2_X1 U506 ( .A(n609), .B(n610), .ZN(n696) );
  NOR2_X1 U507 ( .A1(n657), .A2(n656), .ZN(n658) );
  INV_X1 U508 ( .A(KEYINPUT60), .ZN(n422) );
  XNOR2_X1 U509 ( .A(n742), .B(n386), .ZN(n745) );
  XNOR2_X1 U510 ( .A(n744), .B(n743), .ZN(n386) );
  XNOR2_X1 U511 ( .A(n385), .B(n384), .ZN(G75) );
  INV_X1 U512 ( .A(KEYINPUT53), .ZN(n384) );
  XOR2_X1 U513 ( .A(n740), .B(KEYINPUT119), .Z(n367) );
  AND2_X1 U514 ( .A1(n367), .A2(KEYINPUT120), .ZN(n368) );
  XNOR2_X1 U515 ( .A(G131), .B(G140), .ZN(n369) );
  INV_X1 U516 ( .A(n611), .ZN(n715) );
  XNOR2_X1 U517 ( .A(n488), .B(G478), .ZN(n593) );
  NAND2_X1 U518 ( .A1(n644), .A2(n643), .ZN(n370) );
  NAND2_X1 U519 ( .A1(n607), .A2(KEYINPUT47), .ZN(n371) );
  AND2_X1 U520 ( .A1(n432), .A2(n368), .ZN(n372) );
  AND2_X1 U521 ( .A1(n403), .A2(n693), .ZN(n373) );
  OR2_X1 U522 ( .A1(n715), .A2(n653), .ZN(n374) );
  OR2_X1 U523 ( .A1(n648), .A2(n725), .ZN(n375) );
  BUF_X1 U524 ( .A(n708), .Z(n437) );
  INV_X1 U525 ( .A(n437), .ZN(n479) );
  INV_X1 U526 ( .A(KEYINPUT106), .ZN(n419) );
  INV_X1 U527 ( .A(n755), .ZN(n444) );
  XOR2_X1 U528 ( .A(n677), .B(n676), .Z(n376) );
  XNOR2_X1 U529 ( .A(n746), .B(KEYINPUT59), .ZN(n377) );
  AND2_X1 U530 ( .A1(n660), .A2(n472), .ZN(n378) );
  XOR2_X1 U531 ( .A(n674), .B(KEYINPUT87), .Z(n379) );
  INV_X1 U532 ( .A(G953), .ZN(n759) );
  NAND2_X1 U533 ( .A1(n382), .A2(n722), .ZN(n456) );
  XNOR2_X1 U534 ( .A(n382), .B(n380), .ZN(n723) );
  NAND2_X1 U535 ( .A1(n586), .A2(n382), .ZN(n568) );
  OR2_X1 U536 ( .A1(n619), .A2(n382), .ZN(n381) );
  XNOR2_X2 U537 ( .A(n515), .B(n485), .ZN(n382) );
  NOR2_X1 U538 ( .A1(n364), .A2(n378), .ZN(n468) );
  NAND2_X1 U539 ( .A1(n667), .A2(n666), .ZN(n383) );
  XNOR2_X1 U540 ( .A(n478), .B(n673), .ZN(n477) );
  XNOR2_X1 U541 ( .A(n425), .B(n377), .ZN(n424) );
  NAND2_X1 U542 ( .A1(n393), .A2(n759), .ZN(n385) );
  NAND2_X1 U543 ( .A1(n652), .A2(n650), .ZN(n651) );
  XNOR2_X1 U544 ( .A(n457), .B(n649), .ZN(n652) );
  NAND2_X1 U545 ( .A1(n432), .A2(n367), .ZN(n390) );
  NAND2_X1 U546 ( .A1(n388), .A2(n387), .ZN(n393) );
  NAND2_X1 U547 ( .A1(n707), .A2(n372), .ZN(n387) );
  NAND2_X1 U548 ( .A1(n390), .A2(n741), .ZN(n389) );
  NAND2_X1 U549 ( .A1(n392), .A2(n741), .ZN(n391) );
  INV_X1 U550 ( .A(n707), .ZN(n392) );
  NAND2_X1 U551 ( .A1(n693), .A2(n481), .ZN(n400) );
  AND2_X1 U552 ( .A1(n396), .A2(n693), .ZN(n395) );
  INV_X1 U553 ( .A(n612), .ZN(n404) );
  NAND2_X1 U554 ( .A1(n405), .A2(n416), .ZN(n408) );
  NAND2_X1 U555 ( .A1(n412), .A2(KEYINPUT106), .ZN(n406) );
  INV_X1 U556 ( .A(n593), .ZN(n407) );
  OR2_X1 U557 ( .A1(n593), .A2(KEYINPUT106), .ZN(n410) );
  NAND2_X1 U558 ( .A1(n592), .A2(n419), .ZN(n411) );
  INV_X1 U559 ( .A(n498), .ZN(n415) );
  NAND2_X1 U560 ( .A1(n498), .A2(G902), .ZN(n417) );
  NAND2_X1 U561 ( .A1(n746), .A2(n498), .ZN(n418) );
  XNOR2_X1 U562 ( .A(n421), .B(n523), .ZN(n526) );
  XNOR2_X1 U563 ( .A(n423), .B(n422), .ZN(G60) );
  NAND2_X1 U564 ( .A1(n424), .A2(n444), .ZN(n423) );
  NOR2_X1 U565 ( .A1(G902), .A2(n675), .ZN(n563) );
  NOR2_X1 U566 ( .A1(n611), .A2(n612), .ZN(n427) );
  OR2_X2 U567 ( .A1(n611), .A2(n428), .ZN(n566) );
  AND2_X2 U568 ( .A1(n439), .A2(n567), .ZN(n586) );
  NAND2_X1 U569 ( .A1(n539), .A2(G217), .ZN(n482) );
  NAND2_X1 U570 ( .A1(n723), .A2(n722), .ZN(n726) );
  XNOR2_X1 U571 ( .A(n430), .B(n379), .ZN(G51) );
  NAND2_X1 U572 ( .A1(n477), .A2(n444), .ZN(n430) );
  NOR2_X1 U573 ( .A1(n370), .A2(n469), .ZN(n434) );
  NOR2_X2 U574 ( .A1(n788), .A2(n687), .ZN(n661) );
  NAND2_X1 U575 ( .A1(n777), .A2(G234), .ZN(n486) );
  XNOR2_X2 U576 ( .A(n431), .B(G953), .ZN(n777) );
  INV_X1 U577 ( .A(n638), .ZN(n442) );
  XNOR2_X2 U578 ( .A(n632), .B(KEYINPUT0), .ZN(n638) );
  NAND2_X1 U579 ( .A1(n434), .A2(n466), .ZN(n436) );
  XNOR2_X2 U580 ( .A(n436), .B(KEYINPUT45), .ZN(n760) );
  NOR2_X1 U581 ( .A1(n787), .A2(KEYINPUT44), .ZN(n654) );
  NAND2_X1 U582 ( .A1(n438), .A2(n444), .ZN(n443) );
  XNOR2_X1 U583 ( .A(n678), .B(n376), .ZN(n438) );
  NAND2_X1 U584 ( .A1(n480), .A2(n479), .ZN(n447) );
  XNOR2_X1 U585 ( .A(n776), .B(n445), .ZN(n705) );
  NAND2_X1 U586 ( .A1(n654), .A2(n661), .ZN(n655) );
  INV_X1 U587 ( .A(n736), .ZN(n441) );
  NAND2_X1 U588 ( .A1(n499), .A2(KEYINPUT94), .ZN(n463) );
  NAND2_X1 U589 ( .A1(n760), .A2(n776), .ZN(n662) );
  NAND2_X1 U590 ( .A1(n500), .A2(G119), .ZN(n462) );
  XNOR2_X1 U591 ( .A(n443), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X2 U592 ( .A1(n656), .A2(n374), .ZN(n687) );
  NOR2_X2 U593 ( .A1(n638), .A2(n375), .ZN(n457) );
  NOR2_X1 U594 ( .A1(n750), .A2(G902), .ZN(n550) );
  NAND2_X1 U595 ( .A1(n615), .A2(n371), .ZN(n450) );
  NOR2_X2 U596 ( .A1(n791), .A2(n786), .ZN(n599) );
  INV_X1 U597 ( .A(n645), .ZN(n653) );
  XNOR2_X2 U598 ( .A(n454), .B(KEYINPUT35), .ZN(n787) );
  NAND2_X1 U599 ( .A1(n630), .A2(n631), .ZN(n632) );
  XNOR2_X1 U600 ( .A(n613), .B(KEYINPUT19), .ZN(n630) );
  XNOR2_X2 U601 ( .A(n456), .B(n571), .ZN(n613) );
  XNOR2_X2 U602 ( .A(n460), .B(n458), .ZN(n556) );
  XNOR2_X2 U603 ( .A(n651), .B(n464), .ZN(n788) );
  XNOR2_X2 U604 ( .A(n556), .B(n502), .ZN(n764) );
  NAND2_X1 U605 ( .A1(n468), .A2(n467), .ZN(n466) );
  NAND2_X1 U606 ( .A1(n655), .A2(n679), .ZN(n469) );
  INV_X1 U607 ( .A(n661), .ZN(n471) );
  XNOR2_X2 U608 ( .A(n474), .B(n473), .ZN(n736) );
  INV_X1 U609 ( .A(n613), .ZN(n481) );
  NOR2_X1 U610 ( .A1(n614), .A2(n709), .ZN(n640) );
  AND2_X2 U611 ( .A1(n624), .A2(n623), .ZN(n663) );
  NOR2_X1 U612 ( .A1(n777), .A2(G952), .ZN(n755) );
  AND2_X1 U613 ( .A1(G210), .A2(n564), .ZN(n485) );
  XNOR2_X1 U614 ( .A(n506), .B(n505), .ZN(n507) );
  INV_X1 U615 ( .A(n701), .ZN(n622) );
  XNOR2_X1 U616 ( .A(n508), .B(n507), .ZN(n511) );
  NOR2_X1 U617 ( .A1(n702), .A2(n622), .ZN(n623) );
  XNOR2_X1 U618 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n649) );
  XNOR2_X1 U619 ( .A(n537), .B(n536), .ZN(n538) );
  INV_X1 U620 ( .A(n668), .ZN(n669) );
  INV_X1 U621 ( .A(KEYINPUT120), .ZN(n741) );
  XNOR2_X1 U622 ( .A(KEYINPUT13), .B(G475), .ZN(n498) );
  XNOR2_X1 U623 ( .A(n537), .B(n369), .ZN(n773) );
  XNOR2_X1 U624 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U625 ( .A(n773), .B(n491), .ZN(n497) );
  NAND2_X1 U626 ( .A1(G214), .A2(n558), .ZN(n492) );
  XNOR2_X1 U627 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U628 ( .A(n497), .B(n496), .ZN(n746) );
  NOR2_X1 U629 ( .A1(n593), .A2(n592), .ZN(n635) );
  INV_X1 U630 ( .A(n635), .ZN(n569) );
  INV_X1 U631 ( .A(n503), .ZN(n504) );
  XOR2_X1 U632 ( .A(n504), .B(KEYINPUT18), .Z(n508) );
  NAND2_X1 U633 ( .A1(G224), .A2(n777), .ZN(n506) );
  XNOR2_X1 U634 ( .A(n509), .B(KEYINPUT95), .ZN(n510) );
  XNOR2_X1 U635 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U636 ( .A1(n670), .A2(n668), .ZN(n515) );
  XNOR2_X1 U637 ( .A(n514), .B(KEYINPUT77), .ZN(n564) );
  NAND2_X1 U638 ( .A1(G234), .A2(G237), .ZN(n516) );
  XNOR2_X1 U639 ( .A(n516), .B(KEYINPUT14), .ZN(n518) );
  NAND2_X1 U640 ( .A1(n518), .A2(G952), .ZN(n517) );
  XNOR2_X1 U641 ( .A(n517), .B(KEYINPUT96), .ZN(n735) );
  NOR2_X1 U642 ( .A1(G953), .A2(n735), .ZN(n627) );
  NAND2_X1 U643 ( .A1(G902), .A2(n518), .ZN(n625) );
  NOR2_X1 U644 ( .A1(n777), .A2(n625), .ZN(n519) );
  XNOR2_X1 U645 ( .A(n519), .B(KEYINPUT109), .ZN(n520) );
  NOR2_X1 U646 ( .A1(G900), .A2(n520), .ZN(n521) );
  NOR2_X1 U647 ( .A1(n627), .A2(n521), .ZN(n572) );
  XNOR2_X1 U648 ( .A(KEYINPUT70), .B(G469), .ZN(n528) );
  NAND2_X1 U649 ( .A1(G227), .A2(n777), .ZN(n522) );
  INV_X1 U650 ( .A(n555), .ZN(n525) );
  XOR2_X1 U651 ( .A(KEYINPUT101), .B(KEYINPUT21), .Z(n531) );
  NAND2_X1 U652 ( .A1(G234), .A2(n668), .ZN(n529) );
  XNOR2_X1 U653 ( .A(KEYINPUT20), .B(n529), .ZN(n532) );
  NAND2_X1 U654 ( .A1(G221), .A2(n532), .ZN(n530) );
  XNOR2_X1 U655 ( .A(n531), .B(n530), .ZN(n648) );
  INV_X1 U656 ( .A(n648), .ZN(n712) );
  XOR2_X1 U657 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n534) );
  NAND2_X1 U658 ( .A1(n532), .A2(G217), .ZN(n533) );
  XNOR2_X1 U659 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U660 ( .A(KEYINPUT100), .B(n535), .ZN(n551) );
  XOR2_X1 U661 ( .A(G128), .B(n538), .Z(n549) );
  XOR2_X1 U662 ( .A(KEYINPUT23), .B(KEYINPUT97), .Z(n541) );
  XNOR2_X1 U663 ( .A(n541), .B(n540), .ZN(n545) );
  XOR2_X1 U664 ( .A(KEYINPUT71), .B(KEYINPUT24), .Z(n543) );
  XNOR2_X1 U665 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U666 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U667 ( .A(KEYINPUT5), .B(KEYINPUT78), .Z(n553) );
  XNOR2_X1 U668 ( .A(G131), .B(KEYINPUT102), .ZN(n552) );
  XNOR2_X1 U669 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U670 ( .A(n555), .B(n554), .ZN(n562) );
  XOR2_X1 U671 ( .A(n556), .B(n557), .Z(n560) );
  NAND2_X1 U672 ( .A1(n558), .A2(G210), .ZN(n559) );
  XNOR2_X1 U673 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U674 ( .A(n562), .B(n561), .ZN(n675) );
  XNOR2_X2 U675 ( .A(n563), .B(G472), .ZN(n611) );
  XNOR2_X1 U676 ( .A(n566), .B(n565), .ZN(n567) );
  NOR2_X1 U677 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U678 ( .A(KEYINPUT110), .B(n570), .ZN(n792) );
  INV_X1 U679 ( .A(KEYINPUT91), .ZN(n571) );
  NOR2_X1 U680 ( .A1(n648), .A2(n572), .ZN(n573) );
  NAND2_X1 U681 ( .A1(n645), .A2(n573), .ZN(n612) );
  XOR2_X1 U682 ( .A(n614), .B(KEYINPUT111), .Z(n574) );
  NOR2_X1 U683 ( .A1(n575), .A2(n574), .ZN(n591) );
  NAND2_X1 U684 ( .A1(n366), .A2(n591), .ZN(n576) );
  NOR2_X1 U685 ( .A1(KEYINPUT84), .A2(n688), .ZN(n577) );
  NOR2_X1 U686 ( .A1(n792), .A2(n577), .ZN(n579) );
  NAND2_X1 U687 ( .A1(n407), .A2(n592), .ZN(n699) );
  INV_X1 U688 ( .A(n699), .ZN(n621) );
  NOR2_X1 U689 ( .A1(n609), .A2(n621), .ZN(n727) );
  INV_X1 U690 ( .A(n727), .ZN(n642) );
  NAND2_X1 U691 ( .A1(KEYINPUT85), .A2(n642), .ZN(n578) );
  NAND2_X1 U692 ( .A1(n579), .A2(n578), .ZN(n585) );
  NOR2_X1 U693 ( .A1(n727), .A2(KEYINPUT69), .ZN(n580) );
  NAND2_X1 U694 ( .A1(n694), .A2(n580), .ZN(n581) );
  NAND2_X1 U695 ( .A1(KEYINPUT84), .A2(n581), .ZN(n582) );
  NOR2_X1 U696 ( .A1(KEYINPUT85), .A2(n582), .ZN(n583) );
  NOR2_X1 U697 ( .A1(KEYINPUT47), .A2(n583), .ZN(n584) );
  NOR2_X1 U698 ( .A1(n585), .A2(n584), .ZN(n601) );
  NAND2_X1 U699 ( .A1(n723), .A2(n586), .ZN(n588) );
  XOR2_X1 U700 ( .A(KEYINPUT73), .B(KEYINPUT39), .Z(n587) );
  NAND2_X1 U701 ( .A1(n620), .A2(n609), .ZN(n590) );
  INV_X1 U702 ( .A(n591), .ZN(n595) );
  NAND2_X1 U703 ( .A1(n593), .A2(n592), .ZN(n725) );
  XNOR2_X1 U704 ( .A(KEYINPUT41), .B(n594), .ZN(n737) );
  NOR2_X1 U705 ( .A1(n595), .A2(n737), .ZN(n596) );
  XNOR2_X1 U706 ( .A(n596), .B(KEYINPUT42), .ZN(n786) );
  XOR2_X1 U707 ( .A(KEYINPUT46), .B(KEYINPUT88), .Z(n597) );
  XNOR2_X1 U708 ( .A(KEYINPUT65), .B(n597), .ZN(n598) );
  XNOR2_X1 U709 ( .A(n599), .B(n598), .ZN(n600) );
  NAND2_X1 U710 ( .A1(n601), .A2(n600), .ZN(n608) );
  NAND2_X1 U711 ( .A1(n694), .A2(KEYINPUT69), .ZN(n602) );
  NAND2_X1 U712 ( .A1(n642), .A2(n602), .ZN(n604) );
  INV_X1 U713 ( .A(KEYINPUT85), .ZN(n603) );
  NAND2_X1 U714 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U715 ( .A1(KEYINPUT84), .A2(n688), .ZN(n605) );
  NAND2_X1 U716 ( .A1(n606), .A2(n605), .ZN(n607) );
  INV_X1 U717 ( .A(KEYINPUT108), .ZN(n610) );
  XNOR2_X1 U718 ( .A(n789), .B(KEYINPUT89), .ZN(n615) );
  XNOR2_X1 U719 ( .A(n616), .B(KEYINPUT48), .ZN(n624) );
  NAND2_X1 U720 ( .A1(n373), .A2(n722), .ZN(n617) );
  NOR2_X1 U721 ( .A1(n479), .A2(n617), .ZN(n618) );
  XNOR2_X1 U722 ( .A(n618), .B(KEYINPUT43), .ZN(n619) );
  NAND2_X1 U723 ( .A1(n621), .A2(n620), .ZN(n701) );
  BUF_X2 U724 ( .A(n663), .Z(n776) );
  NOR2_X1 U725 ( .A1(G898), .A2(n759), .ZN(n767) );
  INV_X1 U726 ( .A(n625), .ZN(n626) );
  NAND2_X1 U727 ( .A1(n767), .A2(n626), .ZN(n629) );
  INV_X1 U728 ( .A(n627), .ZN(n628) );
  NAND2_X1 U729 ( .A1(n629), .A2(n628), .ZN(n631) );
  XNOR2_X1 U730 ( .A(KEYINPUT34), .B(KEYINPUT81), .ZN(n633) );
  NAND2_X1 U731 ( .A1(n787), .A2(KEYINPUT44), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n715), .A2(n636), .ZN(n718) );
  NOR2_X1 U733 ( .A1(n718), .A2(n638), .ZN(n637) );
  XNOR2_X1 U734 ( .A(n637), .B(KEYINPUT31), .ZN(n698) );
  NOR2_X1 U735 ( .A1(n638), .A2(n715), .ZN(n639) );
  NAND2_X1 U736 ( .A1(n640), .A2(n639), .ZN(n681) );
  NAND2_X1 U737 ( .A1(n698), .A2(n681), .ZN(n641) );
  NAND2_X1 U738 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U739 ( .A(n645), .B(KEYINPUT107), .ZN(n711) );
  NOR2_X1 U740 ( .A1(n657), .A2(n646), .ZN(n647) );
  XNOR2_X1 U741 ( .A(KEYINPUT82), .B(n647), .ZN(n650) );
  NAND2_X1 U742 ( .A1(n437), .A2(n652), .ZN(n656) );
  XNOR2_X1 U743 ( .A(n658), .B(KEYINPUT90), .ZN(n659) );
  NAND2_X1 U744 ( .A1(n659), .A2(n711), .ZN(n679) );
  INV_X1 U745 ( .A(KEYINPUT44), .ZN(n660) );
  NAND2_X1 U746 ( .A1(n662), .A2(KEYINPUT2), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n663), .B(KEYINPUT79), .ZN(n664) );
  NAND2_X1 U748 ( .A1(n665), .A2(n760), .ZN(n666) );
  XOR2_X1 U749 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n672) );
  XNOR2_X1 U750 ( .A(n670), .B(KEYINPUT92), .ZN(n671) );
  XNOR2_X1 U751 ( .A(n672), .B(n671), .ZN(n673) );
  INV_X1 U752 ( .A(KEYINPUT56), .ZN(n674) );
  XOR2_X1 U753 ( .A(n675), .B(KEYINPUT93), .Z(n677) );
  XOR2_X1 U754 ( .A(KEYINPUT62), .B(KEYINPUT113), .Z(n676) );
  XNOR2_X1 U755 ( .A(G101), .B(n679), .ZN(G3) );
  NOR2_X1 U756 ( .A1(n681), .A2(n696), .ZN(n680) );
  XOR2_X1 U757 ( .A(G104), .B(n680), .Z(G6) );
  NOR2_X1 U758 ( .A1(n699), .A2(n681), .ZN(n686) );
  XOR2_X1 U759 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n683) );
  XNOR2_X1 U760 ( .A(G107), .B(KEYINPUT26), .ZN(n682) );
  XNOR2_X1 U761 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U762 ( .A(KEYINPUT114), .B(n684), .ZN(n685) );
  XNOR2_X1 U763 ( .A(n686), .B(n685), .ZN(G9) );
  XOR2_X1 U764 ( .A(n687), .B(G110), .Z(G12) );
  NOR2_X1 U765 ( .A1(n688), .A2(n699), .ZN(n692) );
  XOR2_X1 U766 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n690) );
  XNOR2_X1 U767 ( .A(G128), .B(KEYINPUT117), .ZN(n689) );
  XNOR2_X1 U768 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U769 ( .A(n692), .B(n691), .ZN(G30) );
  NAND2_X1 U770 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U771 ( .A(n695), .B(G146), .ZN(G48) );
  NOR2_X1 U772 ( .A1(n698), .A2(n696), .ZN(n697) );
  XOR2_X1 U773 ( .A(G113), .B(n697), .Z(G15) );
  NOR2_X1 U774 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U775 ( .A(G116), .B(n700), .Z(G18) );
  XNOR2_X1 U776 ( .A(G134), .B(n701), .ZN(G36) );
  XOR2_X1 U777 ( .A(G140), .B(n702), .Z(n703) );
  XNOR2_X1 U778 ( .A(KEYINPUT118), .B(n703), .ZN(G42) );
  AND2_X1 U779 ( .A1(n760), .A2(n776), .ZN(n704) );
  NOR2_X1 U780 ( .A1(KEYINPUT2), .A2(n705), .ZN(n706) );
  NAND2_X1 U781 ( .A1(n706), .A2(n760), .ZN(n707) );
  NAND2_X1 U782 ( .A1(n709), .A2(n437), .ZN(n710) );
  XNOR2_X1 U783 ( .A(n710), .B(KEYINPUT50), .ZN(n717) );
  NOR2_X1 U784 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U785 ( .A(KEYINPUT49), .B(n713), .Z(n714) );
  NOR2_X1 U786 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U787 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U788 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U789 ( .A(KEYINPUT51), .B(n720), .ZN(n721) );
  NOR2_X1 U790 ( .A1(n737), .A2(n721), .ZN(n732) );
  NOR2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U792 ( .A1(n725), .A2(n724), .ZN(n729) );
  NOR2_X1 U793 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U794 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U795 ( .A1(n730), .A2(n736), .ZN(n731) );
  NOR2_X1 U796 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U797 ( .A(n733), .B(KEYINPUT52), .ZN(n734) );
  NOR2_X1 U798 ( .A1(n735), .A2(n734), .ZN(n739) );
  NOR2_X1 U799 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U800 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U801 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n743) );
  NAND2_X1 U802 ( .A1(n365), .A2(G469), .ZN(n742) );
  NOR2_X1 U803 ( .A1(n755), .A2(n745), .ZN(G54) );
  NAND2_X1 U804 ( .A1(G478), .A2(n751), .ZN(n747) );
  XNOR2_X1 U805 ( .A(n748), .B(n747), .ZN(n749) );
  NOR2_X1 U806 ( .A1(n755), .A2(n749), .ZN(G63) );
  XOR2_X1 U807 ( .A(n750), .B(KEYINPUT121), .Z(n753) );
  NAND2_X1 U808 ( .A1(n365), .A2(G217), .ZN(n752) );
  XNOR2_X1 U809 ( .A(n753), .B(n752), .ZN(n754) );
  NOR2_X1 U810 ( .A1(n755), .A2(n754), .ZN(G66) );
  XNOR2_X1 U811 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n771) );
  NAND2_X1 U812 ( .A1(G224), .A2(G953), .ZN(n756) );
  XNOR2_X1 U813 ( .A(n756), .B(KEYINPUT122), .ZN(n757) );
  XNOR2_X1 U814 ( .A(KEYINPUT61), .B(n757), .ZN(n758) );
  NAND2_X1 U815 ( .A1(G898), .A2(n758), .ZN(n762) );
  NAND2_X1 U816 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U817 ( .A1(n762), .A2(n761), .ZN(n769) );
  XNOR2_X1 U818 ( .A(n763), .B(G101), .ZN(n765) );
  XNOR2_X1 U819 ( .A(n765), .B(n764), .ZN(n766) );
  NOR2_X1 U820 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U821 ( .A(n769), .B(n768), .Z(n770) );
  XNOR2_X1 U822 ( .A(n771), .B(n770), .ZN(G69) );
  XNOR2_X1 U823 ( .A(n772), .B(n773), .ZN(n774) );
  XOR2_X1 U824 ( .A(n775), .B(n774), .Z(n780) );
  XOR2_X1 U825 ( .A(n776), .B(n780), .Z(n778) );
  NAND2_X1 U826 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U827 ( .A(KEYINPUT125), .B(n779), .Z(n784) );
  XNOR2_X1 U828 ( .A(G227), .B(n780), .ZN(n781) );
  NAND2_X1 U829 ( .A1(n781), .A2(G900), .ZN(n782) );
  NAND2_X1 U830 ( .A1(G953), .A2(n782), .ZN(n783) );
  NAND2_X1 U831 ( .A1(n784), .A2(n783), .ZN(G72) );
  XOR2_X1 U832 ( .A(G137), .B(KEYINPUT126), .Z(n785) );
  XNOR2_X1 U833 ( .A(n786), .B(n785), .ZN(G39) );
  XOR2_X1 U834 ( .A(n787), .B(G122), .Z(G24) );
  XOR2_X1 U835 ( .A(n788), .B(G119), .Z(G21) );
  XNOR2_X1 U836 ( .A(G125), .B(KEYINPUT37), .ZN(n790) );
  XNOR2_X1 U837 ( .A(n790), .B(n789), .ZN(G27) );
  XOR2_X1 U838 ( .A(n791), .B(G131), .Z(G33) );
  XOR2_X1 U839 ( .A(G143), .B(n792), .Z(G45) );
endmodule

