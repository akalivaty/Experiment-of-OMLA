

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595;

  XNOR2_X1 U327 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U328 ( .A(n416), .B(n415), .ZN(n574) );
  XNOR2_X1 U329 ( .A(n403), .B(n312), .ZN(n313) );
  XOR2_X1 U330 ( .A(n443), .B(KEYINPUT20), .Z(n295) );
  AND2_X1 U331 ( .A1(G229GAT), .A2(G233GAT), .ZN(n296) );
  XOR2_X1 U332 ( .A(n441), .B(n440), .Z(n297) );
  NOR2_X1 U333 ( .A1(n578), .A2(n562), .ZN(n387) );
  NOR2_X1 U334 ( .A1(n406), .A2(n570), .ZN(n407) );
  XNOR2_X1 U335 ( .A(n302), .B(n296), .ZN(n303) );
  XNOR2_X1 U336 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n415) );
  NOR2_X1 U337 ( .A1(n464), .A2(n528), .ZN(n460) );
  NOR2_X1 U338 ( .A1(n587), .A2(n486), .ZN(n487) );
  XNOR2_X1 U339 ( .A(n314), .B(n313), .ZN(n315) );
  INV_X1 U340 ( .A(G169GAT), .ZN(n453) );
  XOR2_X1 U341 ( .A(n451), .B(n450), .Z(n519) );
  XOR2_X1 U342 ( .A(KEYINPUT38), .B(n489), .Z(n499) );
  XNOR2_X1 U343 ( .A(n453), .B(KEYINPUT122), .ZN(n454) );
  XNOR2_X1 U344 ( .A(n455), .B(n454), .ZN(G1348GAT) );
  XOR2_X1 U345 ( .A(G141GAT), .B(G22GAT), .Z(n431) );
  XOR2_X1 U346 ( .A(G1GAT), .B(KEYINPUT69), .Z(n366) );
  XNOR2_X1 U347 ( .A(n431), .B(n366), .ZN(n299) );
  XOR2_X1 U348 ( .A(G15GAT), .B(G197GAT), .Z(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n304) );
  XOR2_X1 U350 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n301) );
  XNOR2_X1 U351 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U353 ( .A(n305), .B(KEYINPUT71), .Z(n314) );
  XOR2_X1 U354 ( .A(G50GAT), .B(G29GAT), .Z(n307) );
  XNOR2_X1 U355 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U357 ( .A(n308), .B(KEYINPUT68), .Z(n310) );
  XNOR2_X1 U358 ( .A(G36GAT), .B(KEYINPUT67), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n403) );
  XNOR2_X1 U360 ( .A(G169GAT), .B(G43GAT), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n311), .B(G113GAT), .ZN(n440) );
  XNOR2_X1 U362 ( .A(n440), .B(KEYINPUT66), .ZN(n312) );
  INV_X1 U363 ( .A(n315), .ZN(n578) );
  XOR2_X1 U364 ( .A(n315), .B(KEYINPUT72), .Z(n531) );
  XOR2_X1 U365 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n439) );
  XOR2_X1 U366 ( .A(KEYINPUT86), .B(KEYINPUT88), .Z(n317) );
  XNOR2_X1 U367 ( .A(KEYINPUT1), .B(KEYINPUT87), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n336) );
  XOR2_X1 U369 ( .A(G148GAT), .B(G155GAT), .Z(n319) );
  XNOR2_X1 U370 ( .A(G141GAT), .B(G120GAT), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U372 ( .A(KEYINPUT6), .B(G57GAT), .Z(n321) );
  XNOR2_X1 U373 ( .A(G113GAT), .B(G127GAT), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U375 ( .A(n323), .B(n322), .Z(n328) );
  XOR2_X1 U376 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n325) );
  NAND2_X1 U377 ( .A1(G225GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U379 ( .A(G1GAT), .B(n326), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U381 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n430) );
  XOR2_X1 U382 ( .A(G85GAT), .B(n430), .Z(n330) );
  XOR2_X1 U383 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n444) );
  XNOR2_X1 U384 ( .A(n444), .B(G134GAT), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U386 ( .A(n332), .B(n331), .Z(n334) );
  XNOR2_X1 U387 ( .A(G29GAT), .B(G162GAT), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U389 ( .A(n336), .B(n335), .Z(n514) );
  XOR2_X1 U390 ( .A(G92GAT), .B(G204GAT), .Z(n338) );
  XNOR2_X1 U391 ( .A(G36GAT), .B(G190GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n348) );
  XOR2_X1 U393 ( .A(KEYINPUT90), .B(G64GAT), .Z(n340) );
  XNOR2_X1 U394 ( .A(G169GAT), .B(KEYINPUT89), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U396 ( .A(G8GAT), .B(G211GAT), .Z(n355) );
  XOR2_X1 U397 ( .A(KEYINPUT78), .B(n355), .Z(n342) );
  XOR2_X1 U398 ( .A(G197GAT), .B(KEYINPUT21), .Z(n419) );
  XNOR2_X1 U399 ( .A(G218GAT), .B(n419), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U401 ( .A(n344), .B(n343), .Z(n346) );
  NAND2_X1 U402 ( .A1(G226GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n354) );
  XNOR2_X1 U405 ( .A(G183GAT), .B(KEYINPUT83), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n349), .B(G176GAT), .ZN(n350) );
  XOR2_X1 U407 ( .A(n350), .B(KEYINPUT17), .Z(n352) );
  XNOR2_X1 U408 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n351) );
  XOR2_X1 U409 ( .A(n352), .B(n351), .Z(n449) );
  INV_X1 U410 ( .A(n449), .ZN(n353) );
  XOR2_X1 U411 ( .A(n354), .B(n353), .Z(n493) );
  XOR2_X1 U412 ( .A(G155GAT), .B(G78GAT), .Z(n421) );
  XOR2_X1 U413 ( .A(n355), .B(n421), .Z(n357) );
  NAND2_X1 U414 ( .A1(G231GAT), .A2(G233GAT), .ZN(n356) );
  XOR2_X1 U415 ( .A(n357), .B(n356), .Z(n370) );
  XOR2_X1 U416 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n363) );
  XNOR2_X1 U417 ( .A(G57GAT), .B(G64GAT), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n358), .B(KEYINPUT13), .ZN(n378) );
  XOR2_X1 U419 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n360) );
  XNOR2_X1 U420 ( .A(G183GAT), .B(KEYINPUT14), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n378), .B(n361), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n365) );
  INV_X1 U424 ( .A(G71GAT), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n368) );
  XNOR2_X1 U426 ( .A(G22GAT), .B(n366), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n372) );
  XNOR2_X1 U429 ( .A(G15GAT), .B(G127GAT), .ZN(n446) );
  INV_X1 U430 ( .A(n446), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n587) );
  INV_X1 U432 ( .A(n587), .ZN(n556) );
  XOR2_X1 U433 ( .A(KEYINPUT108), .B(n556), .Z(n568) );
  XOR2_X1 U434 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n374) );
  NAND2_X1 U435 ( .A1(G230GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U437 ( .A(n375), .B(KEYINPUT33), .Z(n380) );
  XOR2_X1 U438 ( .A(G92GAT), .B(G85GAT), .Z(n377) );
  XNOR2_X1 U439 ( .A(G99GAT), .B(G106GAT), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n395) );
  XNOR2_X1 U441 ( .A(n395), .B(n378), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U443 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n382) );
  XNOR2_X1 U444 ( .A(G176GAT), .B(G78GAT), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U446 ( .A(n384), .B(n383), .Z(n386) );
  XOR2_X1 U447 ( .A(G120GAT), .B(G71GAT), .Z(n448) );
  XOR2_X1 U448 ( .A(G204GAT), .B(G148GAT), .Z(n420) );
  XNOR2_X1 U449 ( .A(n448), .B(n420), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n583) );
  XNOR2_X1 U451 ( .A(n583), .B(KEYINPUT41), .ZN(n562) );
  XNOR2_X1 U452 ( .A(n387), .B(KEYINPUT46), .ZN(n388) );
  NOR2_X1 U453 ( .A1(n568), .A2(n388), .ZN(n389) );
  XNOR2_X1 U454 ( .A(n389), .B(KEYINPUT109), .ZN(n406) );
  XOR2_X1 U455 ( .A(KEYINPUT79), .B(KEYINPUT77), .Z(n391) );
  XNOR2_X1 U456 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U458 ( .A(n392), .B(KEYINPUT78), .Z(n394) );
  XOR2_X1 U459 ( .A(G190GAT), .B(G134GAT), .Z(n441) );
  XNOR2_X1 U460 ( .A(G43GAT), .B(n441), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n394), .B(n393), .ZN(n399) );
  XOR2_X1 U462 ( .A(G218GAT), .B(G162GAT), .Z(n422) );
  XOR2_X1 U463 ( .A(n395), .B(n422), .Z(n397) );
  NAND2_X1 U464 ( .A1(G232GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U466 ( .A(n399), .B(n398), .Z(n405) );
  XOR2_X1 U467 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n401) );
  XNOR2_X1 U468 ( .A(KEYINPUT76), .B(KEYINPUT64), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U471 ( .A(n405), .B(n404), .Z(n560) );
  INV_X1 U472 ( .A(n560), .ZN(n570) );
  XNOR2_X1 U473 ( .A(n407), .B(KEYINPUT47), .ZN(n413) );
  XOR2_X1 U474 ( .A(KEYINPUT36), .B(n560), .Z(n591) );
  NAND2_X1 U475 ( .A1(n587), .A2(n591), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n408), .B(KEYINPUT110), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n409), .B(KEYINPUT45), .ZN(n410) );
  NOR2_X1 U478 ( .A1(n583), .A2(n410), .ZN(n411) );
  NAND2_X1 U479 ( .A1(n411), .A2(n531), .ZN(n412) );
  NAND2_X1 U480 ( .A1(n413), .A2(n412), .ZN(n414) );
  XNOR2_X1 U481 ( .A(KEYINPUT48), .B(n414), .ZN(n545) );
  NAND2_X1 U482 ( .A1(n493), .A2(n545), .ZN(n416) );
  XOR2_X1 U483 ( .A(G211GAT), .B(KEYINPUT23), .Z(n418) );
  XNOR2_X1 U484 ( .A(G50GAT), .B(G106GAT), .ZN(n417) );
  XNOR2_X1 U485 ( .A(n418), .B(n417), .ZN(n426) );
  XOR2_X1 U486 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U487 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n435) );
  XOR2_X1 U490 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n428) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U493 ( .A(n429), .B(KEYINPUT85), .Z(n433) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n464) );
  INV_X1 U497 ( .A(n464), .ZN(n436) );
  NOR2_X1 U498 ( .A1(n574), .A2(n436), .ZN(n437) );
  NAND2_X1 U499 ( .A1(n514), .A2(n437), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n452) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n297), .B(n442), .ZN(n443) );
  XNOR2_X1 U503 ( .A(G99GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n295), .B(n445), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U506 ( .A(n449), .B(n448), .Z(n450) );
  INV_X1 U507 ( .A(n519), .ZN(n528) );
  NAND2_X1 U508 ( .A1(n452), .A2(n528), .ZN(n567) );
  NOR2_X1 U509 ( .A1(n531), .A2(n567), .ZN(n455) );
  XOR2_X1 U510 ( .A(KEYINPUT34), .B(KEYINPUT95), .Z(n475) );
  NOR2_X1 U511 ( .A1(n570), .A2(n556), .ZN(n456) );
  XNOR2_X1 U512 ( .A(KEYINPUT16), .B(n456), .ZN(n470) );
  NAND2_X1 U513 ( .A1(n528), .A2(n493), .ZN(n457) );
  NAND2_X1 U514 ( .A1(n464), .A2(n457), .ZN(n458) );
  XOR2_X1 U515 ( .A(KEYINPUT25), .B(n458), .Z(n461) );
  INV_X1 U516 ( .A(n493), .ZN(n517) );
  XOR2_X1 U517 ( .A(KEYINPUT27), .B(KEYINPUT91), .Z(n459) );
  XOR2_X1 U518 ( .A(n517), .B(n459), .Z(n465) );
  XNOR2_X1 U519 ( .A(n460), .B(KEYINPUT26), .ZN(n576) );
  NAND2_X1 U520 ( .A1(n465), .A2(n576), .ZN(n546) );
  NAND2_X1 U521 ( .A1(n461), .A2(n546), .ZN(n462) );
  NAND2_X1 U522 ( .A1(n462), .A2(n514), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n463), .B(KEYINPUT92), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n464), .B(KEYINPUT28), .ZN(n525) );
  INV_X1 U525 ( .A(n525), .ZN(n498) );
  INV_X1 U526 ( .A(n514), .ZN(n575) );
  NAND2_X1 U527 ( .A1(n465), .A2(n575), .ZN(n466) );
  NOR2_X1 U528 ( .A1(n498), .A2(n466), .ZN(n530) );
  XNOR2_X1 U529 ( .A(n519), .B(KEYINPUT84), .ZN(n467) );
  NAND2_X1 U530 ( .A1(n530), .A2(n467), .ZN(n468) );
  NAND2_X1 U531 ( .A1(n469), .A2(n468), .ZN(n485) );
  NAND2_X1 U532 ( .A1(n470), .A2(n485), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n471), .B(KEYINPUT93), .ZN(n501) );
  NOR2_X1 U534 ( .A1(n583), .A2(n531), .ZN(n472) );
  XOR2_X1 U535 ( .A(KEYINPUT75), .B(n472), .Z(n488) );
  NAND2_X1 U536 ( .A1(n501), .A2(n488), .ZN(n473) );
  XOR2_X1 U537 ( .A(KEYINPUT94), .B(n473), .Z(n482) );
  NAND2_X1 U538 ( .A1(n482), .A2(n575), .ZN(n474) );
  XNOR2_X1 U539 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  NAND2_X1 U541 ( .A1(n482), .A2(n493), .ZN(n477) );
  XNOR2_X1 U542 ( .A(n477), .B(KEYINPUT96), .ZN(n478) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n478), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U545 ( .A1(n528), .A2(n482), .ZN(n479) );
  XNOR2_X1 U546 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U547 ( .A(G15GAT), .B(n481), .Z(G1326GAT) );
  NAND2_X1 U548 ( .A1(n482), .A2(n498), .ZN(n483) );
  XNOR2_X1 U549 ( .A(n483), .B(KEYINPUT98), .ZN(n484) );
  XNOR2_X1 U550 ( .A(G22GAT), .B(n484), .ZN(G1327GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT39), .B(KEYINPUT99), .Z(n491) );
  NAND2_X1 U552 ( .A1(n591), .A2(n485), .ZN(n486) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(n487), .Z(n513) );
  NAND2_X1 U554 ( .A1(n513), .A2(n488), .ZN(n489) );
  NAND2_X1 U555 ( .A1(n499), .A2(n575), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U557 ( .A(G29GAT), .B(n492), .Z(G1328GAT) );
  NAND2_X1 U558 ( .A1(n499), .A2(n493), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT100), .Z(n496) );
  NAND2_X1 U561 ( .A1(n528), .A2(n499), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U563 ( .A(n497), .B(G43GAT), .Z(G1330GAT) );
  NAND2_X1 U564 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U566 ( .A1(n315), .A2(n562), .ZN(n512) );
  NAND2_X1 U567 ( .A1(n501), .A2(n512), .ZN(n509) );
  NOR2_X1 U568 ( .A1(n514), .A2(n509), .ZN(n502) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n502), .Z(n503) );
  XNOR2_X1 U570 ( .A(KEYINPUT42), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n517), .A2(n509), .ZN(n505) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(KEYINPUT101), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n519), .A2(n509), .ZN(n507) );
  XNOR2_X1 U575 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n506) );
  XNOR2_X1 U576 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(n508), .ZN(G1334GAT) );
  NOR2_X1 U578 ( .A1(n525), .A2(n509), .ZN(n511) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n510) );
  XNOR2_X1 U580 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U581 ( .A1(n513), .A2(n512), .ZN(n524) );
  NOR2_X1 U582 ( .A1(n514), .A2(n524), .ZN(n515) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n515), .Z(n516) );
  XNOR2_X1 U584 ( .A(KEYINPUT104), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U585 ( .A1(n517), .A2(n524), .ZN(n518) );
  XOR2_X1 U586 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  NOR2_X1 U587 ( .A1(n519), .A2(n524), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(KEYINPUT105), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT106), .B(KEYINPUT44), .Z(n523) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(KEYINPUT107), .ZN(n522) );
  XNOR2_X1 U592 ( .A(n523), .B(n522), .ZN(n527) );
  NOR2_X1 U593 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U594 ( .A(n527), .B(n526), .Z(G1339GAT) );
  AND2_X1 U595 ( .A1(n528), .A2(n545), .ZN(n529) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n538) );
  NOR2_X1 U597 ( .A1(n531), .A2(n538), .ZN(n532) );
  XOR2_X1 U598 ( .A(G113GAT), .B(n532), .Z(G1340GAT) );
  NOR2_X1 U599 ( .A1(n562), .A2(n538), .ZN(n534) );
  XNOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT111), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n535), .Z(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n537) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(KEYINPUT113), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n541) );
  INV_X1 U606 ( .A(n538), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n542), .A2(n568), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n539), .B(KEYINPUT112), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U611 ( .A1(n542), .A2(n570), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n545), .A2(n575), .ZN(n547) );
  NOR2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(KEYINPUT115), .ZN(n559) );
  NOR2_X1 U616 ( .A1(n578), .A2(n559), .ZN(n549) );
  XOR2_X1 U617 ( .A(KEYINPUT116), .B(n549), .Z(n550) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  NOR2_X1 U619 ( .A1(n562), .A2(n559), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n552) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n551) );
  XNOR2_X1 U622 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U623 ( .A(KEYINPUT52), .B(n553), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n556), .A2(n559), .ZN(n558) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  NOR2_X1 U630 ( .A1(n567), .A2(n562), .ZN(n566) );
  XOR2_X1 U631 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n563) );
  XNOR2_X1 U633 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  INV_X1 U635 ( .A(n567), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n571), .A2(n568), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(KEYINPUT58), .ZN(n573) );
  XNOR2_X1 U640 ( .A(G190GAT), .B(n573), .ZN(G1351GAT) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n582) );
  NOR2_X1 U643 ( .A1(n578), .A2(n582), .ZN(n581) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n579), .B(KEYINPUT59), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n585) );
  INV_X1 U648 ( .A(n582), .ZN(n592) );
  NAND2_X1 U649 ( .A1(n592), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(n586), .ZN(G1353GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n589) );
  NAND2_X1 U653 ( .A1(n592), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(G211GAT), .B(n590), .ZN(G1354GAT) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n594) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

