//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  INV_X1    g0005(.A(G264), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI22_X1  g0008(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G97), .C2(G257), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G244), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G68), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(new_n216), .B1(new_n217), .B2(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n215), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(G20), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n222), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n224), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n208), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n205), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n207), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n248), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT73), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n201), .B1(new_n217), .B2(G58), .ZN(new_n255));
  INV_X1    g0055(.A(G20), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT7), .B1(new_n258), .B2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT7), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n260), .B(new_n256), .C1(new_n262), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n259), .A2(new_n217), .A3(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G159), .ZN(new_n268));
  INV_X1    g0068(.A(G68), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT64), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT64), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G68), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n272), .A3(G58), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n202), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(KEYINPUT73), .A3(G20), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n257), .A2(new_n266), .A3(new_n268), .A4(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT16), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT74), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n227), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n256), .B1(new_n273), .B2(new_n202), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n283), .B(new_n254), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n261), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n263), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT72), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(new_n263), .B2(G33), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT7), .B1(new_n289), .B2(G20), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n263), .A3(G33), .ZN(new_n291));
  AOI21_X1  g0091(.A(KEYINPUT72), .B1(new_n261), .B2(KEYINPUT3), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(new_n262), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(new_n260), .A3(new_n256), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n290), .A2(G68), .A3(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n284), .A2(new_n295), .A3(KEYINPUT16), .A4(new_n268), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n276), .A2(KEYINPUT74), .A3(new_n277), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n280), .A2(new_n282), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n281), .A2(new_n227), .ZN(new_n299));
  INV_X1    g0099(.A(G1), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(G13), .A3(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT69), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n301), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n282), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT69), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n304), .B(new_n307), .C1(G1), .C2(new_n256), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT8), .B(G58), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n305), .B2(new_n310), .ZN(new_n312));
  INV_X1    g0112(.A(G41), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n228), .B1(new_n261), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n288), .A2(new_n286), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n211), .A2(G1698), .ZN(new_n316));
  OR2_X1    g0116(.A1(G223), .A2(G1698), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n291), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G87), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n314), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n300), .B1(G41), .B2(G45), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n220), .ZN(new_n323));
  INV_X1    g0123(.A(G274), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n320), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G200), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(G190), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n298), .A2(new_n312), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT17), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n298), .A2(new_n312), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  NOR4_X1   g0133(.A1(new_n320), .A2(new_n323), .A3(new_n333), .A4(new_n325), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n327), .B2(G169), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT18), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n332), .A2(KEYINPUT18), .A3(new_n336), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n309), .B(KEYINPUT70), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n261), .A2(G20), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT15), .B(G87), .Z(new_n344));
  AOI22_X1  g0144(.A1(new_n342), .A2(new_n267), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n256), .B2(new_n247), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(new_n282), .B1(new_n247), .B2(new_n305), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n299), .B1(G1), .B2(new_n256), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n247), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n205), .B2(new_n258), .ZN(new_n352));
  INV_X1    g0152(.A(new_n258), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n353), .A2(new_n220), .A3(G1698), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n350), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n325), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n314), .A2(new_n216), .A3(new_n321), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n349), .B1(G200), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G190), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n360), .B2(new_n358), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n331), .A2(new_n341), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n308), .A2(new_n210), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n305), .A2(new_n210), .ZN(new_n364));
  INV_X1    g0164(.A(new_n343), .ZN(new_n365));
  INV_X1    g0165(.A(G150), .ZN(new_n366));
  INV_X1    g0166(.A(new_n267), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n309), .A2(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n256), .B1(new_n201), .B2(new_n210), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n282), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n363), .A2(new_n364), .A3(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(KEYINPUT9), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n356), .B1(new_n322), .B2(new_n211), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT68), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n375));
  INV_X1    g0175(.A(G1698), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n258), .A2(G222), .A3(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n375), .B(new_n377), .C1(new_n247), .C2(new_n258), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n350), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n371), .A2(KEYINPUT9), .B1(G200), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n374), .A2(G190), .A3(new_n379), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n372), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT10), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT10), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n372), .A2(new_n381), .A3(new_n385), .A4(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n371), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n380), .B2(G179), .ZN(new_n389));
  AOI21_X1  g0189(.A(G169), .B1(new_n374), .B2(new_n379), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n217), .A2(new_n256), .B1(new_n210), .B2(new_n367), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n365), .A2(new_n247), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n282), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT11), .ZN(new_n397));
  INV_X1    g0197(.A(new_n217), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(KEYINPUT12), .A3(new_n305), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n269), .B1(new_n348), .B2(KEYINPUT12), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT12), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(new_n301), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n397), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT13), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n286), .A2(new_n405), .A3(G226), .A4(new_n376), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n286), .A2(new_n405), .A3(G232), .A4(G1698), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G97), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n350), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n314), .A2(G238), .A3(new_n321), .ZN(new_n411));
  AND4_X1   g0211(.A1(new_n404), .A2(new_n410), .A3(new_n356), .A4(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n325), .B1(new_n409), .B2(new_n350), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n404), .B1(new_n413), .B2(new_n411), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n403), .B1(new_n416), .B2(G200), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n360), .B2(new_n416), .ZN(new_n418));
  OAI21_X1  g0218(.A(G169), .B1(new_n412), .B2(new_n414), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT14), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n415), .A2(G179), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT14), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n422), .B(G169), .C1(new_n412), .C2(new_n414), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n403), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT71), .ZN(new_n427));
  INV_X1    g0227(.A(G169), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n358), .A2(new_n428), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n358), .A2(G179), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n349), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NOR4_X1   g0232(.A1(new_n362), .A2(new_n393), .A3(new_n427), .A4(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n315), .B(new_n291), .C1(G250), .C2(G1698), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n376), .A2(G257), .ZN(new_n435));
  INV_X1    g0235(.A(G294), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n434), .A2(new_n435), .B1(new_n261), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n300), .A2(G45), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT5), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT76), .B1(new_n439), .B2(G41), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT76), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(new_n313), .A3(KEYINPUT5), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n438), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n439), .A2(G41), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n350), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n437), .A2(new_n350), .B1(G264), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(G274), .A3(new_n444), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n428), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n333), .A3(new_n447), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n289), .A2(KEYINPUT81), .A3(new_n256), .A4(G87), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT81), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n256), .B(new_n291), .C1(new_n292), .C2(new_n262), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(new_n212), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n455), .A3(KEYINPUT22), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT22), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n258), .A2(new_n457), .A3(new_n256), .A4(G87), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT82), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G116), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G20), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n256), .A2(G107), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n465), .B(KEYINPUT23), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT24), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n463), .B1(new_n456), .B2(new_n460), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT24), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n466), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n299), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n306), .B1(G1), .B2(new_n261), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT25), .B1(new_n305), .B2(new_n205), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n305), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n474), .A2(G107), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n451), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT83), .ZN(new_n481));
  AND4_X1   g0281(.A1(new_n470), .A2(new_n461), .A3(new_n464), .A4(new_n466), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n470), .B1(new_n469), .B2(new_n466), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n282), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G200), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n448), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(G190), .B2(new_n448), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(new_n487), .A3(new_n478), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n480), .A2(new_n481), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n481), .B1(new_n480), .B2(new_n488), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT78), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n314), .A2(G250), .A3(new_n438), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  OR2_X1    g0293(.A1(G238), .A2(G1698), .ZN(new_n494));
  INV_X1    g0294(.A(G244), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G1698), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n462), .B1(new_n293), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT77), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(KEYINPUT77), .B(new_n462), .C1(new_n293), .C2(new_n497), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n493), .B1(new_n502), .B2(new_n350), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n438), .A2(new_n324), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n491), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n314), .B1(new_n500), .B2(new_n501), .ZN(new_n507));
  NOR4_X1   g0307(.A1(new_n507), .A2(KEYINPUT78), .A3(new_n504), .A4(new_n493), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n333), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n501), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n315), .A2(new_n291), .A3(new_n494), .A4(new_n496), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT77), .B1(new_n511), .B2(new_n462), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n350), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(new_n505), .A3(new_n492), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT78), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n503), .A2(new_n491), .A3(new_n505), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n428), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n315), .A2(new_n256), .A3(G68), .A4(new_n291), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT19), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n256), .B1(new_n408), .B2(new_n519), .ZN(new_n520));
  NOR4_X1   g0320(.A1(KEYINPUT79), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT79), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G87), .A2(G97), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(new_n205), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n520), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(G97), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n519), .B1(new_n365), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n518), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n282), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n344), .A2(new_n301), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT80), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT80), .ZN(new_n533));
  AOI211_X1 g0333(.A(new_n533), .B(new_n530), .C1(new_n528), .C2(new_n282), .ZN(new_n534));
  INV_X1    g0334(.A(new_n344), .ZN(new_n535));
  OAI22_X1  g0335(.A1(new_n532), .A2(new_n534), .B1(new_n535), .B2(new_n473), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n509), .A2(new_n517), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(G190), .B1(new_n506), .B2(new_n508), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n515), .A2(new_n516), .A3(G200), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n474), .A2(G87), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n532), .B2(new_n534), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n206), .A2(G1698), .ZN(new_n544));
  INV_X1    g0344(.A(G257), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n376), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n289), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n353), .A2(G303), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n314), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n447), .ZN(new_n550));
  AOI211_X1 g0350(.A(new_n208), .B(new_n350), .C1(new_n443), .C2(new_n444), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n306), .B(G116), .C1(G1), .C2(new_n261), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n300), .A2(new_n207), .A3(G13), .A4(G20), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n281), .A2(new_n227), .B1(G20), .B2(new_n207), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G283), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n556), .B(new_n256), .C1(G33), .C2(new_n526), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT20), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n555), .A2(KEYINPUT20), .A3(new_n557), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n553), .B(new_n554), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n552), .A2(G179), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n547), .A2(new_n548), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n350), .ZN(new_n563));
  INV_X1    g0363(.A(new_n551), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n563), .A2(G190), .A3(new_n447), .A4(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n560), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n565), .B(new_n566), .C1(new_n552), .C2(new_n485), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n560), .A2(G169), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n552), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n563), .A2(new_n447), .A3(new_n564), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n571), .A2(KEYINPUT21), .A3(G169), .A4(new_n560), .ZN(new_n572));
  AND4_X1   g0372(.A1(new_n561), .A2(new_n567), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n301), .A2(G97), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n259), .A2(G107), .A3(new_n265), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT75), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n205), .A2(KEYINPUT6), .A3(G97), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n526), .A2(new_n205), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G97), .A2(G107), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n578), .B1(new_n581), .B2(KEYINPUT6), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G20), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n259), .A2(KEYINPUT75), .A3(new_n265), .A4(G107), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n267), .A2(G77), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n577), .A2(new_n583), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n574), .B1(new_n586), .B2(new_n282), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n473), .A2(new_n526), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n376), .B(new_n291), .C1(new_n292), .C2(new_n262), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n495), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n286), .A2(new_n405), .A3(G250), .A4(G1698), .ZN(new_n593));
  AND2_X1   g0393(.A1(KEYINPUT4), .A2(G244), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n286), .A2(new_n405), .A3(new_n594), .A4(new_n376), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n593), .A2(new_n595), .A3(new_n556), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n350), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n545), .B(new_n350), .C1(new_n443), .C2(new_n444), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n447), .A3(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n587), .A2(new_n589), .B1(new_n428), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n314), .B1(new_n592), .B2(new_n596), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n603), .A2(new_n550), .A3(new_n599), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n333), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n550), .B1(new_n597), .B2(new_n350), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n485), .B1(new_n606), .B2(new_n600), .ZN(new_n607));
  NOR4_X1   g0407(.A1(new_n603), .A2(new_n550), .A3(new_n599), .A4(new_n360), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI211_X1 g0409(.A(new_n574), .B(new_n588), .C1(new_n586), .C2(new_n282), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n602), .A2(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n537), .A2(new_n543), .A3(new_n573), .A4(new_n611), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n489), .A2(new_n490), .A3(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n433), .A2(new_n613), .ZN(G372));
  NAND2_X1  g0414(.A1(new_n514), .A2(new_n428), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n509), .A2(new_n536), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n360), .B1(new_n515), .B2(new_n516), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT84), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n541), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(KEYINPUT84), .B(new_n540), .C1(new_n532), .C2(new_n534), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n514), .A2(G200), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n617), .B1(new_n622), .B2(KEYINPUT85), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT85), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n619), .A2(new_n620), .A3(new_n624), .A4(new_n621), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n616), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n488), .A2(new_n611), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n572), .A2(new_n570), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n561), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT86), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n628), .A2(KEYINPUT86), .A3(new_n561), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n480), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n626), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n623), .A2(new_n625), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n602), .A2(new_n605), .ZN(new_n637));
  INV_X1    g0437(.A(new_n616), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n537), .A2(new_n543), .A3(new_n637), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n616), .B1(new_n640), .B2(KEYINPUT26), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n634), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n433), .A2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n432), .A2(new_n418), .B1(new_n403), .B2(new_n424), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT17), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n330), .B(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n341), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n391), .B1(new_n647), .B2(new_n387), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n643), .A2(new_n648), .ZN(G369));
  AND2_X1   g0449(.A1(new_n631), .A2(new_n632), .ZN(new_n650));
  INV_X1    g0450(.A(G13), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(G20), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n300), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n566), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n650), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n573), .B(KEYINPUT87), .Z(new_n662));
  OAI211_X1 g0462(.A(new_n661), .B(G330), .C1(new_n660), .C2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n489), .A2(new_n490), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n658), .B1(new_n472), .B2(new_n479), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n449), .B1(G179), .B2(new_n448), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n484), .B2(new_n478), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n658), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n659), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n484), .A2(new_n478), .A3(new_n487), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT83), .B1(new_n674), .B2(new_n669), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n480), .A2(new_n481), .A3(new_n488), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n629), .A4(new_n659), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n672), .A2(new_n673), .A3(new_n677), .ZN(G399));
  INV_X1    g0478(.A(new_n230), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G1), .ZN(new_n682));
  OR3_X1    g0482(.A1(new_n521), .A2(new_n524), .A3(G116), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n682), .A2(new_n683), .B1(new_n225), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G330), .ZN(new_n687));
  AND4_X1   g0487(.A1(new_n573), .A2(new_n537), .A3(new_n543), .A4(new_n611), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(new_n675), .A3(new_n676), .A4(new_n659), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT89), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT89), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n665), .A2(new_n691), .A3(new_n688), .A4(new_n659), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n604), .A2(new_n552), .A3(G179), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n694), .B(new_n446), .C1(new_n506), .C2(new_n508), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n604), .A2(new_n552), .A3(G179), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(new_n448), .A3(new_n514), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n515), .A2(new_n516), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(KEYINPUT30), .A3(new_n446), .A4(new_n694), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n697), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n702), .A2(new_n703), .A3(new_n658), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(new_n702), .B2(new_n658), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n687), .B1(new_n693), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n537), .A2(new_n543), .A3(new_n636), .A4(new_n637), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n622), .A2(KEYINPUT85), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n711), .A2(new_n538), .A3(new_n625), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n488), .B(new_n611), .C1(new_n669), .C2(new_n629), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n638), .B(new_n710), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n636), .B1(new_n626), .B2(new_n637), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n709), .B1(new_n716), .B2(new_n659), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n642), .A2(new_n659), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(KEYINPUT29), .ZN(new_n719));
  OR3_X1    g0519(.A1(new_n708), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n686), .B1(new_n720), .B2(new_n300), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT90), .ZN(G364));
  AOI21_X1  g0522(.A(new_n300), .B1(new_n652), .B2(G45), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n680), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n664), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n662), .A2(new_n660), .ZN(new_n727));
  INV_X1    g0527(.A(new_n661), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n726), .B1(G330), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n289), .A2(new_n679), .ZN(new_n731));
  INV_X1    g0531(.A(G45), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n226), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n731), .B(new_n733), .C1(new_n248), .C2(new_n732), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n353), .A2(new_n679), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G355), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n734), .B(new_n736), .C1(G116), .C2(new_n230), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n227), .B1(G20), .B2(new_n428), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n256), .A2(new_n360), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n333), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n256), .A2(G190), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n744), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(G58), .A2(new_n746), .B1(new_n749), .B2(G77), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n333), .A2(new_n485), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n485), .A2(G179), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n743), .A2(new_n753), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n750), .B1(new_n210), .B2(new_n752), .C1(new_n212), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n747), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n353), .B(new_n755), .C1(G107), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n256), .B1(new_n759), .B2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G97), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n751), .A2(new_n747), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n269), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT91), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n747), .A2(new_n759), .ZN(new_n766));
  INV_X1    g0566(.A(G159), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n758), .A2(new_n765), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n760), .A2(new_n436), .ZN(new_n771));
  INV_X1    g0571(.A(G326), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n752), .A2(new_n772), .B1(new_n748), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n766), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n771), .B(new_n774), .C1(G329), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n757), .A2(G283), .ZN(new_n777));
  XOR2_X1   g0577(.A(KEYINPUT33), .B(G317), .Z(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n778), .A2(new_n763), .B1(new_n745), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT93), .ZN(new_n781));
  INV_X1    g0581(.A(G303), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n353), .B1(new_n754), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT92), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n776), .A2(new_n777), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n770), .A2(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n737), .A2(new_n742), .B1(new_n741), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n740), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n725), .B(new_n787), .C1(new_n729), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n730), .A2(new_n789), .ZN(G396));
  INV_X1    g0590(.A(KEYINPUT96), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n431), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n349), .A2(new_n658), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n792), .A2(new_n361), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n432), .A2(new_n658), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n718), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n792), .A2(new_n361), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n642), .A2(new_n659), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(new_n708), .ZN(new_n802));
  INV_X1    g0602(.A(new_n725), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n754), .A2(new_n210), .B1(new_n756), .B2(new_n269), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT95), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n289), .B1(new_n219), .B2(new_n760), .ZN(new_n807));
  INV_X1    g0607(.A(new_n752), .ZN(new_n808));
  INV_X1    g0608(.A(new_n763), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G137), .A2(new_n808), .B1(new_n809), .B2(G150), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n767), .B2(new_n748), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G143), .B2(new_n746), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT94), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n806), .B(new_n807), .C1(new_n813), .C2(KEYINPUT34), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(KEYINPUT34), .B2(new_n813), .C1(new_n815), .C2(new_n766), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n745), .A2(new_n436), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n752), .A2(new_n782), .B1(new_n754), .B2(new_n205), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G311), .B2(new_n775), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n749), .A2(G116), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n353), .B1(new_n756), .B2(new_n212), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G283), .B2(new_n809), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n819), .A2(new_n762), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n816), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n741), .A2(new_n738), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n824), .A2(new_n741), .B1(new_n247), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n826), .B(new_n725), .C1(new_n739), .C2(new_n796), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n804), .A2(new_n827), .ZN(G384));
  AOI21_X1  g0628(.A(new_n691), .B1(new_n613), .B2(new_n659), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n689), .A2(KEYINPUT89), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n707), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n403), .A2(new_n658), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n424), .A2(KEYINPUT99), .A3(new_n403), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT99), .B1(new_n424), .B2(new_n403), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n418), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT100), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n424), .A2(new_n403), .A3(new_n658), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n836), .B1(new_n835), .B2(new_n837), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n796), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT102), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT40), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n831), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n706), .B1(new_n690), .B2(new_n692), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n842), .B1(new_n845), .B2(new_n840), .ZN(new_n846));
  INV_X1    g0646(.A(new_n294), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n260), .B1(new_n293), .B2(new_n256), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n847), .A2(new_n848), .A3(new_n269), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n257), .A2(new_n268), .A3(new_n275), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n277), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(new_n296), .A3(new_n282), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n312), .ZN(new_n853));
  INV_X1    g0653(.A(new_n656), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT18), .B1(new_n332), .B2(new_n336), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n338), .B(new_n335), .C1(new_n298), .C2(new_n312), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n856), .B1(new_n646), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n853), .A2(new_n336), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n330), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT101), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n856), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n330), .A2(new_n862), .A3(KEYINPUT101), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n332), .B1(new_n336), .B2(new_n854), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n868), .A2(new_n861), .A3(new_n330), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n860), .B(KEYINPUT38), .C1(new_n867), .C2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n332), .A2(new_n854), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n331), .B2(new_n341), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n861), .B1(new_n868), .B2(new_n330), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n871), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n844), .A2(new_n846), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT40), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n840), .B1(new_n693), .B2(new_n707), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n863), .A2(new_n864), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n855), .A3(new_n866), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n869), .B1(new_n882), .B2(KEYINPUT37), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n855), .B1(new_n331), .B2(new_n341), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n871), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n870), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(new_n886), .A3(new_n843), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT103), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n831), .A2(new_n433), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n889), .B(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(G330), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n433), .B1(new_n717), .B2(new_n719), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n648), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n833), .A2(new_n834), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n659), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n885), .B2(new_n870), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n870), .A2(new_n876), .A3(new_n898), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n792), .A2(new_n658), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n800), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n838), .A2(new_n839), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n903), .A2(new_n886), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n341), .A2(new_n854), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n901), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n894), .B(new_n909), .Z(new_n910));
  XNOR2_X1  g0710(.A(new_n892), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n300), .B2(new_n652), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n226), .A2(G77), .A3(new_n273), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n210), .A2(G68), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT98), .ZN(new_n915));
  OAI211_X1 g0715(.A(G1), .B(new_n651), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(G20), .B(new_n228), .C1(new_n582), .C2(KEYINPUT35), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n207), .B(new_n917), .C1(KEYINPUT35), .C2(new_n582), .ZN(new_n918));
  XNOR2_X1  g0718(.A(KEYINPUT97), .B(KEYINPUT36), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n912), .A2(new_n916), .A3(new_n920), .ZN(G367));
  OAI21_X1  g0721(.A(new_n611), .B1(new_n610), .B2(new_n659), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n637), .A2(new_n658), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT105), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n926), .A2(new_n677), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT42), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n926), .A2(new_n480), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n659), .B1(new_n929), .B2(new_n637), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n659), .B1(new_n619), .B2(new_n620), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n638), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n626), .B2(new_n932), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT104), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n672), .A2(new_n926), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n680), .B(KEYINPUT41), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT45), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n677), .A2(new_n673), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n945), .B1(new_n926), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n924), .B(KEYINPUT105), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n948), .A2(new_n677), .A3(KEYINPUT45), .A4(new_n673), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n926), .A2(new_n946), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT44), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(KEYINPUT106), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n947), .A2(new_n949), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n926), .A2(new_n946), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n672), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT107), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n956), .A2(new_n960), .A3(new_n957), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n629), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(new_n658), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n677), .B1(new_n671), .B2(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n663), .A2(KEYINPUT108), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT109), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n708), .A2(new_n717), .A3(new_n719), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT109), .B1(new_n720), .B2(new_n967), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT110), .B1(new_n956), .B2(new_n957), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT110), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n953), .A2(new_n974), .A3(new_n672), .A4(new_n955), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n962), .A2(new_n971), .A3(new_n972), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n944), .B1(new_n977), .B2(new_n970), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n941), .B(new_n942), .C1(new_n978), .C2(new_n724), .ZN(new_n979));
  INV_X1    g0779(.A(new_n731), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n742), .B1(new_n230), .B2(new_n535), .C1(new_n242), .C2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n754), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(G116), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT46), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n984), .B(new_n293), .C1(new_n205), .C2(new_n760), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G311), .A2(new_n808), .B1(new_n746), .B2(G303), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT111), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(KEYINPUT111), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G283), .A2(new_n749), .B1(new_n775), .B2(G317), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n757), .A2(G97), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n985), .B(new_n991), .C1(G294), .C2(new_n809), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n353), .B1(new_n757), .B2(G77), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n210), .B2(new_n748), .C1(new_n269), .C2(new_n760), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G143), .A2(new_n808), .B1(new_n746), .B2(G150), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n219), .B2(new_n754), .C1(new_n767), .C2(new_n763), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(G137), .C2(new_n775), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT113), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n998), .B(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n803), .B1(new_n1001), .B2(new_n741), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n981), .B(new_n1002), .C1(new_n935), .C2(new_n788), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n979), .A2(new_n1003), .ZN(G387));
  NAND2_X1  g0804(.A1(new_n971), .A2(new_n972), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n720), .A2(new_n967), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(new_n680), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n293), .B1(new_n207), .B2(new_n756), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G317), .A2(new_n746), .B1(new_n749), .B2(G303), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n773), .B2(new_n763), .C1(new_n779), .C2(new_n752), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT48), .ZN(new_n1011));
  INV_X1    g0811(.A(G283), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(new_n1012), .B2(new_n760), .C1(new_n436), .C2(new_n754), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT49), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n1014), .B2(new_n1013), .C1(new_n772), .C2(new_n766), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G50), .A2(new_n746), .B1(new_n809), .B2(new_n310), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n247), .B2(new_n754), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n990), .B1(new_n269), .B2(new_n748), .C1(new_n366), .C2(new_n766), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n289), .B1(new_n535), .B2(new_n760), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n767), .B2(new_n752), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n803), .B1(new_n1023), .B2(new_n741), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n671), .B2(new_n788), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n342), .A2(new_n210), .ZN(new_n1026));
  AOI21_X1  g0826(.A(G45), .B1(new_n1026), .B2(KEYINPUT50), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n683), .B1(G68), .B2(G77), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(KEYINPUT50), .C2(new_n1026), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n731), .C1(new_n732), .C2(new_n239), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n683), .A2(new_n735), .B1(new_n205), .B2(new_n679), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT114), .Z(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1025), .B1(new_n742), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n968), .B2(new_n724), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1007), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT115), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1007), .A2(KEYINPUT115), .A3(new_n1035), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(G393));
  NAND2_X1  g0840(.A1(new_n926), .A2(new_n740), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n742), .B1(new_n526), .B2(new_n230), .C1(new_n252), .C2(new_n980), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n760), .A2(new_n247), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n752), .A2(new_n366), .B1(new_n745), .B2(new_n767), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT51), .Z(new_n1045));
  AOI211_X1 g0845(.A(new_n1043), .B(new_n1045), .C1(new_n342), .C2(new_n749), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n293), .B1(G143), .B2(new_n775), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n212), .B2(new_n756), .C1(new_n398), .C2(new_n754), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT116), .Z(new_n1049));
  OAI211_X1 g0849(.A(new_n1046), .B(new_n1049), .C1(new_n210), .C2(new_n763), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G283), .A2(new_n982), .B1(new_n749), .B2(G294), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n782), .B2(new_n763), .C1(new_n779), .C2(new_n766), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n258), .B(new_n1052), .C1(G116), .C2(new_n761), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G317), .A2(new_n808), .B1(new_n746), .B2(G311), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT52), .Z(new_n1055));
  OAI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(new_n205), .C2(new_n756), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1050), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n803), .B1(new_n1057), .B2(new_n741), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1041), .A2(new_n1042), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n976), .A2(new_n958), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n1060), .B2(new_n723), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n977), .A2(new_n680), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1060), .A2(new_n1005), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(G390));
  INV_X1    g0865(.A(new_n899), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n900), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n904), .B1(new_n800), .B2(new_n902), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1066), .B(new_n1067), .C1(new_n1068), .C2(new_n897), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n659), .B(new_n799), .C1(new_n714), .C2(new_n715), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT117), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1070), .A2(new_n1071), .A3(new_n902), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n1070), .B2(new_n902), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1072), .A2(new_n1073), .A3(new_n904), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n877), .A2(new_n896), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1069), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NOR4_X1   g0876(.A1(new_n845), .A2(new_n687), .A3(new_n797), .A4(new_n904), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n708), .A2(new_n796), .A3(new_n905), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1069), .B(new_n1079), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n831), .A2(G330), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n904), .B1(new_n1082), .B2(new_n797), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1073), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1070), .A2(new_n1071), .A3(new_n902), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1086), .A3(new_n1079), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n905), .B1(new_n708), .B2(new_n796), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n903), .B1(new_n1088), .B2(new_n1077), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n831), .A2(G330), .A3(new_n433), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n893), .A2(new_n1091), .A3(new_n648), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1081), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1078), .A2(new_n1080), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n680), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1078), .A2(new_n724), .A3(new_n1080), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT119), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1066), .A2(new_n1067), .A3(new_n738), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n760), .A2(new_n767), .ZN(new_n1101));
  INV_X1    g0901(.A(G137), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n258), .B1(new_n756), .B2(new_n210), .C1(new_n1102), .C2(new_n763), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(G125), .C2(new_n775), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n745), .A2(new_n815), .B1(new_n748), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n982), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT53), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n754), .B2(new_n366), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1106), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(G128), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1104), .B(new_n1110), .C1(new_n1111), .C2(new_n752), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n752), .A2(new_n1012), .B1(new_n763), .B2(new_n205), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G97), .B2(new_n749), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n1115), .A2(KEYINPUT118), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(KEYINPUT118), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n745), .A2(new_n207), .B1(new_n756), .B2(new_n269), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1043), .B(new_n1118), .C1(G294), .C2(new_n775), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1116), .A2(new_n353), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n754), .A2(new_n212), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1112), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1122), .A2(new_n741), .B1(new_n309), .B2(new_n825), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1100), .A2(new_n725), .A3(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1098), .A2(new_n1099), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1099), .B1(new_n1098), .B2(new_n1124), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1097), .B1(new_n1125), .B2(new_n1126), .ZN(G378));
  INV_X1    g0927(.A(KEYINPUT40), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n877), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n880), .B2(new_n843), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1128), .B1(new_n1130), .B2(new_n846), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n887), .ZN(new_n1132));
  OAI21_X1  g0932(.A(G330), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n371), .A2(new_n656), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n387), .B2(new_n392), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n391), .B(new_n1134), .C1(new_n384), .C2(new_n386), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT55), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT55), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT56), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1140), .A2(new_n1141), .A3(KEYINPUT56), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n909), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1148), .A2(new_n906), .A3(new_n901), .A4(new_n908), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1133), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n888), .A2(G330), .A3(new_n1149), .A4(new_n1147), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1096), .A2(new_n1093), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n680), .B1(new_n1153), .B2(KEYINPUT57), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1096), .A2(new_n1093), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1155), .A2(KEYINPUT57), .A3(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n825), .A2(new_n210), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n748), .A2(new_n1102), .B1(new_n760), .B2(new_n366), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G125), .A2(new_n808), .B1(new_n809), .B2(G132), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n754), .B2(new_n1105), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G128), .C2(new_n746), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT59), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n775), .B2(G124), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G33), .B1(new_n757), .B2(G159), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n313), .B1(new_n247), .B2(new_n754), .C1(new_n535), .C2(new_n748), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n289), .B(new_n1168), .C1(G68), .C2(new_n761), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n745), .A2(new_n205), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n752), .A2(new_n207), .B1(new_n763), .B2(new_n526), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(G283), .C2(new_n775), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1169), .B(new_n1172), .C1(new_n219), .C2(new_n756), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT58), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G41), .B1(new_n289), .B2(G33), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1167), .B(new_n1174), .C1(G50), .C2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n803), .B1(new_n1176), .B2(new_n741), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1159), .B(new_n1177), .C1(new_n1148), .C2(new_n739), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT120), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n1156), .B2(new_n724), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1158), .A2(new_n1180), .ZN(G375));
  INV_X1    g0981(.A(KEYINPUT122), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1090), .B2(new_n724), .ZN(new_n1183));
  AOI211_X1 g0983(.A(KEYINPUT122), .B(new_n723), .C1(new_n1087), .C2(new_n1089), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n904), .A2(new_n738), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n535), .A2(new_n760), .B1(new_n1012), .B2(new_n745), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G107), .A2(new_n749), .B1(new_n775), .B2(G303), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n436), .B2(new_n752), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(G97), .C2(new_n982), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n258), .B1(new_n757), .B2(G77), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT123), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1189), .B(new_n1191), .C1(new_n207), .C2(new_n763), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n745), .A2(new_n1102), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n756), .A2(new_n219), .B1(new_n760), .B2(new_n210), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n293), .B(new_n1194), .C1(G150), .C2(new_n749), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n808), .A2(G132), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT124), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n763), .A2(new_n1105), .B1(new_n766), .B2(new_n1111), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G159), .B2(new_n982), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1195), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1192), .B1(new_n1193), .B2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1201), .A2(new_n741), .B1(new_n269), .B2(new_n825), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1185), .A2(new_n725), .A3(new_n1202), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1183), .A2(new_n1184), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1087), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n943), .B(KEYINPUT121), .Z(new_n1206));
  NAND3_X1  g1006(.A1(new_n1094), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1204), .A2(new_n1207), .ZN(G381));
  AND3_X1   g1008(.A1(new_n1097), .A2(new_n1098), .A3(new_n1124), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1158), .A2(new_n1180), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(G396), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1038), .A2(new_n1211), .A3(new_n1039), .ZN(new_n1212));
  INV_X1    g1012(.A(G390), .ZN(new_n1213));
  INV_X1    g1013(.A(G384), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1213), .A2(new_n979), .A3(new_n1214), .A4(new_n1003), .ZN(new_n1215));
  OR4_X1    g1015(.A1(G381), .A2(new_n1210), .A3(new_n1212), .A4(new_n1215), .ZN(G407));
  OAI211_X1 g1016(.A(G407), .B(G213), .C1(G343), .C2(new_n1210), .ZN(G409));
  INV_X1    g1017(.A(new_n1212), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1211), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(G387), .A2(new_n1213), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n979), .A2(new_n1003), .A3(G390), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1212), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1222), .ZN(new_n1226));
  AOI21_X1  g1026(.A(G390), .B1(new_n979), .B2(new_n1003), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1223), .A2(new_n1228), .A3(KEYINPUT127), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT127), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(G213), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(G343), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G378), .B(new_n1180), .C1(new_n1154), .C2(new_n1157), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1153), .A2(new_n1206), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1180), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1209), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1233), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT126), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1205), .A2(KEYINPUT125), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT60), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1205), .A2(KEYINPUT125), .A3(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1241), .A2(new_n680), .A3(new_n1094), .A4(new_n1243), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1244), .A2(G384), .A3(new_n1204), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1244), .B2(new_n1204), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1238), .A2(new_n1239), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1239), .B1(new_n1238), .B2(new_n1247), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1248), .A2(new_n1249), .A3(KEYINPUT62), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1233), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1233), .A2(G2897), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1244), .A2(new_n1204), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1214), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1244), .A2(G384), .A3(new_n1204), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1254), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1247), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT62), .B1(new_n1253), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1231), .B1(new_n1250), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1226), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1220), .B1(new_n1222), .B2(new_n1221), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1238), .A2(KEYINPUT63), .A3(new_n1247), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1268), .A2(new_n1271), .A3(new_n1262), .A4(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1266), .A2(new_n1273), .ZN(G405));
  NAND2_X1  g1074(.A1(G375), .A2(new_n1209), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1263), .B1(new_n1275), .B2(new_n1234), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1223), .A2(new_n1228), .A3(KEYINPUT127), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1275), .A2(new_n1263), .A3(new_n1234), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1277), .A2(new_n1279), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1281), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n1283), .A2(new_n1276), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1282), .A2(new_n1284), .ZN(G402));
endmodule


