//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT77), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(new_n193), .ZN(new_n195));
  XOR2_X1   g009(.A(G119), .B(G128), .Z(new_n196));
  OR3_X1    g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G128), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n200), .B(new_n202), .C1(G119), .C2(new_n201), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G110), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n197), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G125), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G140), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT75), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n207), .A2(KEYINPUT75), .A3(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT76), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT16), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n208), .A2(KEYINPUT16), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT16), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n220), .B1(new_n212), .B2(new_n213), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(new_n215), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n207), .A2(KEYINPUT75), .A3(G125), .ZN(new_n224));
  XNOR2_X1  g038(.A(G125), .B(G140), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(new_n211), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT76), .B1(new_n226), .B2(new_n220), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n227), .A2(G146), .A3(new_n218), .A4(new_n216), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n205), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n196), .B1(new_n194), .B2(new_n195), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n203), .A2(G110), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n230), .A2(new_n231), .B1(new_n206), .B2(new_n225), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n232), .A2(new_n228), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n191), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT78), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n223), .A2(new_n228), .ZN(new_n237));
  INV_X1    g051(.A(new_n205), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n232), .A2(new_n228), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(new_n190), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT78), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n242), .B(new_n191), .C1(new_n229), .C2(new_n233), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n235), .A2(new_n236), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n241), .A2(new_n243), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(KEYINPUT25), .A3(new_n236), .A4(new_n235), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G217), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(G234), .B2(new_n236), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n247), .A2(new_n235), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n251), .A2(G902), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT79), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(G210), .B1(G237), .B2(G902), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT88), .ZN(new_n261));
  XNOR2_X1  g075(.A(G110), .B(G122), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(G116), .B(G119), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT5), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n199), .A2(G116), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n266), .B(G113), .C1(KEYINPUT5), .C2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n270));
  OAI22_X1  g084(.A1(new_n269), .A2(new_n270), .B1(KEYINPUT2), .B2(G113), .ZN(new_n271));
  XOR2_X1   g085(.A(G116), .B(G119), .Z(new_n272));
  NOR3_X1   g086(.A1(new_n271), .A2(new_n272), .A3(KEYINPUT70), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT2), .A2(G113), .ZN(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT2), .A2(G113), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n274), .B1(new_n280), .B2(new_n265), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n268), .B1(new_n273), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G104), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT3), .B1(new_n283), .B2(G107), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n285));
  INV_X1    g099(.A(G107), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(G104), .ZN(new_n287));
  INV_X1    g101(.A(G101), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n283), .A2(G107), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n284), .A2(new_n287), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n283), .A2(G107), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n286), .A2(G104), .ZN(new_n292));
  OAI21_X1  g106(.A(G101), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n264), .B1(new_n282), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G113), .B1(new_n267), .B2(KEYINPUT5), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(KEYINPUT86), .B(G113), .C1(new_n267), .C2(KEYINPUT5), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(new_n266), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n273), .B2(new_n281), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT87), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n300), .B(KEYINPUT87), .C1(new_n273), .C2(new_n281), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n295), .B1(new_n305), .B2(new_n294), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT0), .A2(G128), .ZN(new_n307));
  OR2_X1    g121(.A1(KEYINPUT0), .A2(G128), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n206), .A2(G143), .ZN(new_n309));
  INV_X1    g123(.A(G143), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(G146), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n307), .B(new_n308), .C1(new_n309), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT64), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n313), .B1(new_n310), .B2(G146), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n206), .A2(KEYINPUT64), .A3(G143), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n310), .A2(G146), .ZN(new_n316));
  INV_X1    g130(.A(new_n307), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n314), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT1), .ZN(new_n321));
  OAI21_X1  g135(.A(G128), .B1(new_n311), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n206), .A2(G143), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n314), .A2(new_n315), .A3(new_n326), .A4(new_n316), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n209), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G224), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n329), .A2(KEYINPUT83), .A3(G953), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT83), .B1(new_n329), .B2(G953), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n330), .A2(KEYINPUT7), .A3(new_n331), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n320), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n332), .B1(new_n320), .B2(new_n328), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n268), .B(new_n294), .C1(new_n273), .C2(new_n281), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n284), .A2(new_n287), .A3(new_n289), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G101), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT4), .A3(new_n290), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n340), .A3(G101), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT70), .B1(new_n271), .B2(new_n272), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n280), .A2(new_n274), .A3(new_n265), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n343), .A2(new_n344), .B1(new_n271), .B2(new_n272), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n336), .B(new_n262), .C1(new_n342), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n335), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n261), .B(new_n236), .C1(new_n306), .C2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n336), .B1(new_n342), .B2(new_n345), .ZN(new_n349));
  INV_X1    g163(.A(new_n262), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT6), .A3(new_n346), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n320), .A2(new_n328), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n330), .A2(new_n331), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT84), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n353), .B(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n349), .A2(new_n357), .A3(new_n350), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n352), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n290), .A2(new_n293), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n303), .B2(new_n304), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n346), .B(new_n335), .C1(new_n362), .C2(new_n295), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n261), .B1(new_n363), .B2(new_n236), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n260), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT89), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n236), .B1(new_n306), .B2(new_n347), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT88), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n368), .A2(new_n259), .A3(new_n359), .A4(new_n348), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT89), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n370), .B(new_n260), .C1(new_n360), .C2(new_n364), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(G234), .A2(G237), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(G952), .A3(new_n188), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(G902), .A3(G953), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT21), .B(G898), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n375), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G214), .B1(G237), .B2(G902), .ZN(new_n381));
  XOR2_X1   g195(.A(new_n381), .B(KEYINPUT82), .Z(new_n382));
  NAND3_X1  g196(.A1(new_n372), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G137), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT11), .A3(G134), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT11), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G137), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(KEYINPUT11), .ZN(new_n389));
  INV_X1    g203(.A(G134), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT65), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT65), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G134), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(KEYINPUT66), .A2(G131), .ZN(new_n395));
  NOR2_X1   g209(.A1(KEYINPUT66), .A2(G131), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n388), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n388), .A2(new_n394), .ZN(new_n399));
  INV_X1    g213(.A(G131), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n314), .A2(new_n316), .A3(new_n315), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n322), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n327), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n294), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT10), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n312), .A2(new_n318), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n339), .A2(new_n409), .A3(new_n341), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n407), .B1(new_n325), .B2(new_n327), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n294), .ZN(new_n412));
  AND4_X1   g226(.A1(new_n402), .A2(new_n408), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n406), .A2(new_n407), .B1(new_n294), .B2(new_n411), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n402), .B1(new_n414), .B2(new_n410), .ZN(new_n415));
  XNOR2_X1  g229(.A(G110), .B(G140), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n188), .A2(G227), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n413), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n402), .A3(new_n410), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n325), .A2(new_n327), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(new_n294), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n361), .B1(new_n327), .B2(new_n404), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n401), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT80), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT12), .B1(new_n401), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AND4_X1   g241(.A1(new_n394), .A2(new_n385), .A3(new_n387), .A4(new_n397), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n400), .B1(new_n388), .B2(new_n394), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT12), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n406), .B1(new_n421), .B2(new_n294), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(new_n433), .B2(new_n401), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n420), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n419), .B1(new_n435), .B2(new_n418), .ZN(new_n436));
  OAI21_X1  g250(.A(G469), .B1(new_n436), .B2(G902), .ZN(new_n437));
  INV_X1    g251(.A(new_n418), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n420), .B(new_n438), .C1(new_n427), .C2(new_n434), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n418), .B1(new_n413), .B2(new_n415), .ZN(new_n440));
  AOI21_X1  g254(.A(G902), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G469), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n441), .A2(KEYINPUT81), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT81), .B1(new_n441), .B2(new_n442), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n437), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT9), .B(G234), .ZN(new_n446));
  OAI21_X1  g260(.A(G221), .B1(new_n446), .B2(G902), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n391), .A2(new_n393), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n310), .A2(G128), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n201), .A2(G143), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT93), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G128), .B(G143), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT93), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n448), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G116), .B(G122), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(new_n286), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n454), .A2(KEYINPUT13), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n460), .B(G134), .C1(KEYINPUT13), .C2(new_n449), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT14), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G122), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(G116), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n286), .B1(new_n466), .B2(KEYINPUT14), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT94), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n458), .A2(new_n286), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n453), .A2(new_n455), .A3(new_n448), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n456), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n462), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n446), .A2(new_n250), .A3(G953), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n462), .B(new_n474), .C1(new_n469), .C2(new_n472), .ZN(new_n477));
  AOI21_X1  g291(.A(G902), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(KEYINPUT15), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  AOI211_X1 g296(.A(G902), .B(new_n480), .C1(new_n476), .C2(new_n477), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G475), .ZN(new_n485));
  INV_X1    g299(.A(new_n397), .ZN(new_n486));
  NOR2_X1   g300(.A1(G237), .A2(G953), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(G143), .A3(G214), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(G143), .B1(new_n487), .B2(G214), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT17), .ZN(new_n492));
  INV_X1    g306(.A(G237), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n188), .A3(G214), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n310), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n397), .A3(new_n488), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n488), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT17), .A3(new_n486), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n223), .A2(new_n500), .A3(new_n228), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n225), .A2(new_n206), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n214), .B2(new_n206), .ZN(new_n503));
  NAND2_X1  g317(.A1(KEYINPUT18), .A2(G131), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n495), .A2(new_n488), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n498), .A2(KEYINPUT18), .A3(G131), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT92), .B(G104), .Z(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n501), .A2(new_n511), .A3(new_n507), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n485), .B1(new_n515), .B2(new_n236), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n501), .A2(new_n511), .A3(new_n507), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n212), .A2(KEYINPUT19), .A3(new_n213), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT19), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT90), .B1(new_n225), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n212), .A2(KEYINPUT90), .A3(KEYINPUT19), .A4(new_n213), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n206), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n228), .A3(KEYINPUT91), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n491), .A2(new_n496), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT91), .B1(new_n524), .B2(new_n228), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n507), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n517), .B1(new_n529), .B2(new_n512), .ZN(new_n530));
  NOR2_X1   g344(.A1(G475), .A2(G902), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT20), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT20), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n524), .A2(new_n228), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n526), .A3(new_n525), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n511), .B1(new_n538), .B2(new_n507), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n534), .B(new_n531), .C1(new_n539), .C2(new_n517), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n516), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n445), .A2(new_n447), .A3(new_n484), .A4(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n383), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n345), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n409), .B1(new_n428), .B2(new_n429), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n400), .B1(G134), .B2(G137), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n448), .B2(G137), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n421), .A2(new_n398), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n548), .A3(KEYINPUT30), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n545), .A2(KEYINPUT67), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT67), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n409), .B(new_n551), .C1(new_n428), .C2(new_n429), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n398), .A2(new_n547), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT68), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n553), .A2(new_n554), .B1(new_n325), .B2(new_n327), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n398), .A2(KEYINPUT68), .A3(new_n547), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n550), .A2(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n544), .B(new_n549), .C1(new_n557), .C2(KEYINPUT30), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT31), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n545), .A2(new_n548), .A3(new_n345), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n487), .A2(G210), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT27), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT26), .B(G101), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n558), .A2(new_n559), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n559), .B1(new_n558), .B2(new_n567), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n550), .A2(new_n552), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n555), .A2(new_n556), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n544), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT28), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n560), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n545), .A2(new_n548), .A3(new_n345), .A4(KEYINPUT28), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n565), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n568), .A2(new_n569), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(G472), .A2(G902), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT71), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT32), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n558), .A2(new_n567), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT31), .ZN(new_n584));
  INV_X1    g398(.A(new_n577), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n558), .A2(new_n559), .A3(new_n567), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT71), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n579), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n581), .A2(new_n582), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n545), .A2(new_n548), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n544), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n576), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT29), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n566), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(G902), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n574), .B(new_n575), .C1(new_n557), .C2(new_n345), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT72), .B1(new_n598), .B2(new_n566), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT72), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n572), .A2(new_n576), .A3(new_n600), .A4(new_n565), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n595), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n565), .B1(new_n558), .B2(new_n560), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n583), .A2(KEYINPUT31), .B1(new_n566), .B2(new_n598), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n580), .B1(new_n605), .B2(new_n586), .ZN(new_n606));
  AOI22_X1  g420(.A1(G472), .A2(new_n604), .B1(new_n606), .B2(KEYINPUT32), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n590), .A2(new_n607), .A3(KEYINPUT73), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT73), .B1(new_n590), .B2(new_n607), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n258), .B(new_n543), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  OAI21_X1  g425(.A(G472), .B1(new_n578), .B2(G902), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n581), .A2(new_n612), .A3(new_n589), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n614));
  INV_X1    g428(.A(new_n447), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n439), .A2(new_n440), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n442), .A3(new_n236), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT81), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n441), .A2(KEYINPUT81), .A3(new_n442), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n615), .B1(new_n621), .B2(new_n437), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n613), .A2(new_n258), .A3(new_n614), .A4(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n445), .A2(new_n252), .A3(new_n256), .A4(new_n447), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n581), .A2(new_n612), .A3(new_n589), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT95), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n476), .A2(new_n477), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT33), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n476), .A2(new_n630), .A3(new_n477), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n479), .A2(G902), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(KEYINPUT96), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n633), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n629), .B2(new_n631), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(new_n478), .B2(G478), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n634), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n541), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n365), .A2(new_n369), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n381), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n641), .A2(new_n379), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n627), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NAND2_X1  g461(.A1(new_n533), .A2(new_n540), .ZN(new_n648));
  INV_X1    g462(.A(new_n484), .ZN(new_n649));
  INV_X1    g463(.A(new_n516), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n648), .A2(new_n380), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT97), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n643), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n541), .A2(KEYINPUT97), .A3(new_n380), .A4(new_n649), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n627), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n239), .A2(new_n240), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n255), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n252), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n251), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n246), .B2(new_n248), .ZN(new_n667));
  INV_X1    g481(.A(new_n664), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT98), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n543), .A2(new_n613), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  AND2_X1   g487(.A1(new_n665), .A2(new_n669), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n590), .A2(new_n607), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT73), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n590), .A2(new_n607), .A3(KEYINPUT73), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n674), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n648), .A2(new_n650), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT99), .B(G900), .Z(new_n681));
  AOI21_X1  g495(.A(new_n375), .B1(new_n681), .B2(new_n377), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n680), .A2(new_n484), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n445), .A2(new_n447), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n643), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n679), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  INV_X1    g501(.A(KEYINPUT100), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n680), .A2(new_n381), .A3(new_n649), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n688), .B1(new_n670), .B2(new_n689), .ZN(new_n690));
  OR3_X1    g504(.A1(new_n670), .A2(new_n688), .A3(new_n689), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n558), .A2(new_n567), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n565), .B1(new_n592), .B2(new_n560), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n236), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n606), .A2(KEYINPUT32), .B1(G472), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n590), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n372), .B(KEYINPUT38), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n690), .A2(new_n691), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n682), .B(KEYINPUT39), .Z(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n684), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT40), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n700), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  NAND2_X1  g521(.A1(new_n677), .A2(new_n678), .ZN(new_n708));
  INV_X1    g522(.A(new_n682), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT102), .B1(new_n640), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n541), .A2(new_n639), .A3(new_n711), .A4(new_n682), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n708), .A2(new_n670), .A3(new_n685), .A4(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT103), .B(G146), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G48));
  INV_X1    g530(.A(new_n616), .ZN(new_n717));
  OAI211_X1 g531(.A(KEYINPUT104), .B(G469), .C1(new_n717), .C2(G902), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n441), .B2(new_n442), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n621), .A3(new_n447), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n257), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n644), .B(new_n723), .C1(new_n608), .C2(new_n609), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  OAI211_X1 g540(.A(new_n656), .B(new_n723), .C1(new_n608), .C2(new_n609), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  NAND3_X1  g542(.A1(new_n541), .A2(new_n380), .A3(new_n484), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n722), .A2(new_n729), .A3(new_n643), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n670), .B(new_n730), .C1(new_n608), .C2(new_n609), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT105), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n708), .A2(new_n733), .A3(new_n670), .A4(new_n730), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  INV_X1    g550(.A(new_n642), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n689), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n722), .A2(new_n379), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n565), .B1(new_n576), .B2(new_n592), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n584), .A2(KEYINPUT106), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n569), .B2(new_n740), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n586), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n579), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n612), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n738), .A2(new_n739), .A3(new_n258), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n612), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n669), .B2(new_n665), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n722), .A2(new_n643), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n713), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n209), .ZN(G27));
  AND2_X1   g568(.A1(new_n369), .A2(new_n381), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n366), .A3(new_n371), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT107), .B1(new_n684), .B2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n366), .A2(new_n371), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n622), .A2(new_n758), .A3(new_n759), .A4(new_n755), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n710), .A2(new_n712), .A3(KEYINPUT42), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n708), .A2(new_n761), .A3(new_n258), .A4(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n607), .B1(KEYINPUT32), .B2(new_n606), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n636), .A2(new_n638), .ZN(new_n765));
  AOI211_X1 g579(.A(new_n637), .B(new_n635), .C1(new_n629), .C2(new_n631), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n680), .A2(new_n767), .A3(new_n709), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n711), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n640), .A2(KEYINPUT102), .A3(new_n709), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n764), .A2(new_n769), .A3(new_n258), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n757), .A2(new_n760), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT42), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n763), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n400), .ZN(G33));
  NAND4_X1  g589(.A1(new_n708), .A2(new_n761), .A3(new_n258), .A4(new_n683), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  OAI21_X1  g591(.A(G469), .B1(new_n436), .B2(KEYINPUT45), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n778), .A2(KEYINPUT108), .B1(KEYINPUT45), .B2(new_n436), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(KEYINPUT108), .B2(new_n778), .ZN(new_n780));
  NAND2_X1  g594(.A1(G469), .A2(G902), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n783));
  OR3_X1    g597(.A1(new_n782), .A2(new_n783), .A3(KEYINPUT46), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n783), .B1(new_n782), .B2(KEYINPUT46), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(KEYINPUT46), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n784), .A2(new_n621), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n447), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n703), .ZN(new_n789));
  INV_X1    g603(.A(new_n756), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n767), .A2(new_n541), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n791), .B(KEYINPUT43), .Z(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n625), .A3(new_n670), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT44), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  INV_X1    g610(.A(KEYINPUT47), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n788), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n787), .A2(KEYINPUT47), .A3(new_n447), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n708), .A2(new_n258), .A3(new_n756), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n713), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  AND4_X1   g617(.A1(new_n670), .A2(new_n769), .A3(new_n747), .A4(new_n770), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n761), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n541), .A2(new_n484), .A3(new_n709), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n541), .A2(KEYINPUT111), .A3(new_n484), .A4(new_n709), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n622), .A2(new_n808), .A3(new_n790), .A4(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n708), .A2(new_n670), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n776), .A2(new_n805), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n774), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n727), .A2(new_n724), .A3(new_n748), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n734), .B2(new_n732), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n516), .B(new_n484), .C1(new_n533), .C2(new_n540), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n640), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n383), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n623), .A2(new_n626), .A3(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n610), .A2(new_n820), .A3(new_n671), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n813), .A2(new_n814), .A3(new_n816), .A4(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n727), .A2(new_n724), .A3(new_n748), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n735), .A2(new_n823), .A3(new_n821), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n679), .A2(new_n810), .B1(new_n804), .B2(new_n761), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n773), .A3(new_n763), .A4(new_n776), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT112), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n670), .B(new_n685), .C1(new_n608), .C2(new_n609), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n753), .B1(new_n829), .B2(new_n683), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n684), .B1(new_n590), .B2(new_n695), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n667), .A2(new_n668), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n832), .A2(KEYINPUT113), .A3(new_n709), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT113), .B1(new_n832), .B2(new_n709), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n831), .B(new_n738), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n830), .A2(KEYINPUT52), .A3(new_n714), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n804), .A2(new_n752), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n686), .A2(new_n714), .A3(new_n837), .A4(new_n835), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n822), .A2(new_n827), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(KEYINPUT114), .A3(new_n845), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n842), .A2(KEYINPUT114), .A3(new_n843), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n774), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n816), .B2(KEYINPUT115), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n735), .A2(new_n823), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT116), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n774), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n816), .A2(KEYINPUT115), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n821), .A2(new_n825), .A3(KEYINPUT53), .A4(new_n776), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n836), .B2(new_n840), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n854), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n845), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n848), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n188), .A2(G952), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n258), .A2(new_n792), .A3(new_n375), .A4(new_n747), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(new_n752), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n756), .A2(new_n374), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n723), .A2(new_n590), .A3(new_n868), .A4(new_n695), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n641), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n722), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n792), .A2(new_n871), .A3(new_n868), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n764), .A2(new_n258), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(KEYINPUT118), .A3(KEYINPUT48), .ZN(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n721), .A2(new_n621), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT110), .Z(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n447), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n790), .B(new_n866), .C1(new_n800), .C2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n697), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n722), .A2(new_n381), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT117), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n866), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT50), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n872), .A2(new_n674), .A3(new_n750), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n869), .A2(new_n680), .A3(new_n767), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n881), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n870), .B(new_n877), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n864), .A2(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n879), .B(KEYINPUT49), .Z(new_n895));
  NAND3_X1  g709(.A1(new_n258), .A2(new_n382), .A3(new_n447), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n896), .A2(new_n696), .A3(new_n791), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n882), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(G75));
  AOI21_X1  g713(.A(new_n236), .B1(new_n861), .B2(new_n845), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n901), .A3(G210), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n352), .A2(new_n358), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n356), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n901), .B1(new_n900), .B2(G210), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n188), .A2(G952), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT56), .B1(new_n900), .B2(G210), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(new_n906), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n909), .A2(new_n913), .ZN(G51));
  AOI211_X1 g728(.A(new_n236), .B(new_n780), .C1(new_n861), .C2(new_n845), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n861), .A2(new_n845), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT54), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n863), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n781), .B(KEYINPUT57), .Z(new_n919));
  AOI21_X1  g733(.A(new_n717), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n915), .B1(new_n920), .B2(KEYINPUT120), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n922));
  INV_X1    g736(.A(new_n919), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n917), .B2(new_n863), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n924), .B2(new_n717), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n910), .B1(new_n921), .B2(new_n925), .ZN(G54));
  NAND3_X1  g740(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n530), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n530), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n910), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT59), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n632), .B1(new_n864), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n918), .A2(new_n632), .A3(new_n932), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n933), .A2(new_n910), .A3(new_n934), .ZN(G63));
  XNOR2_X1  g749(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n250), .A2(new_n236), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n861), .B2(new_n845), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n253), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n941), .A2(new_n910), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n940), .A2(new_n943), .A3(new_n663), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n940), .B2(new_n663), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n942), .B(KEYINPUT61), .C1(new_n944), .C2(new_n945), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(G66));
  INV_X1    g764(.A(new_n378), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n188), .B1(new_n951), .B2(G224), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n824), .B2(new_n188), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n904), .B1(G898), .B2(new_n188), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT123), .Z(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G69));
  NAND2_X1  g770(.A1(new_n830), .A2(new_n714), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT124), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n873), .A2(new_n737), .A3(new_n689), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n787), .A2(new_n447), .A3(new_n702), .A4(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n960), .A2(new_n849), .A3(new_n776), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n802), .A2(new_n795), .A3(new_n958), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n188), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n188), .A2(G900), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT125), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n549), .B1(new_n557), .B2(KEYINPUT30), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(new_n523), .Z(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n958), .A2(new_n706), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n971));
  NOR4_X1   g785(.A1(new_n818), .A2(new_n684), .A3(new_n703), .A4(new_n756), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n708), .A2(new_n972), .A3(new_n258), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n802), .A2(new_n795), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n971), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n976), .A2(new_n188), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n969), .B1(new_n977), .B2(new_n968), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n968), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n969), .B(new_n982), .C1(new_n977), .C2(new_n968), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(G72));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n976), .B2(new_n824), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n558), .A2(new_n560), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT127), .Z(new_n991));
  NAND3_X1  g805(.A1(new_n989), .A2(new_n565), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n846), .A2(new_n847), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n993), .B(new_n988), .C1(new_n692), .C2(new_n603), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n988), .B1(new_n962), .B2(new_n824), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n991), .A2(new_n565), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n910), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n992), .A2(new_n994), .A3(new_n997), .ZN(G57));
endmodule


