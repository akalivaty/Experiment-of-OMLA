

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592;

  AND2_X2 U328 ( .A1(n568), .A2(n567), .ZN(n576) );
  AND2_X2 U329 ( .A1(n366), .A2(n511), .ZN(n371) );
  XNOR2_X2 U330 ( .A(n372), .B(KEYINPUT48), .ZN(n534) );
  NOR2_X2 U331 ( .A1(n371), .A2(n370), .ZN(n372) );
  XNOR2_X2 U332 ( .A(n465), .B(KEYINPUT41), .ZN(n554) );
  XNOR2_X2 U333 ( .A(n345), .B(n344), .ZN(n465) );
  XNOR2_X1 U334 ( .A(KEYINPUT78), .B(n560), .ZN(n577) );
  XOR2_X1 U335 ( .A(n329), .B(n328), .Z(n586) );
  XOR2_X1 U336 ( .A(G148GAT), .B(G78GAT), .Z(n432) );
  AND2_X1 U337 ( .A1(n368), .A2(n296), .ZN(n369) );
  NOR2_X1 U338 ( .A1(n560), .A2(n586), .ZN(n296) );
  XOR2_X1 U339 ( .A(n315), .B(n314), .Z(n560) );
  XOR2_X1 U340 ( .A(n365), .B(n364), .Z(n583) );
  XNOR2_X1 U341 ( .A(n377), .B(n306), .ZN(n307) );
  XNOR2_X1 U342 ( .A(n308), .B(n307), .ZN(n313) );
  INV_X1 U343 ( .A(G204GAT), .ZN(n461) );
  XNOR2_X1 U344 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U345 ( .A(n464), .B(n463), .ZN(G1353GAT) );
  INV_X1 U346 ( .A(KEYINPUT54), .ZN(n394) );
  XOR2_X1 U347 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n298) );
  XNOR2_X1 U348 ( .A(KEYINPUT8), .B(G29GAT), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U350 ( .A(KEYINPUT7), .B(n299), .Z(n364) );
  INV_X1 U351 ( .A(n364), .ZN(n303) );
  XOR2_X1 U352 ( .A(KEYINPUT72), .B(G106GAT), .Z(n301) );
  XNOR2_X1 U353 ( .A(G99GAT), .B(G92GAT), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U355 ( .A(G85GAT), .B(n302), .Z(n340) );
  XOR2_X1 U356 ( .A(n303), .B(n340), .Z(n315) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G190GAT), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n304), .B(G134GAT), .ZN(n451) );
  INV_X1 U359 ( .A(KEYINPUT76), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n451), .B(n305), .ZN(n308) );
  XOR2_X1 U361 ( .A(G36GAT), .B(G218GAT), .Z(n377) );
  NAND2_X1 U362 ( .A1(G232GAT), .A2(G233GAT), .ZN(n306) );
  XOR2_X1 U363 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n310) );
  XNOR2_X1 U364 ( .A(KEYINPUT10), .B(KEYINPUT77), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U366 ( .A(G50GAT), .B(G162GAT), .Z(n430) );
  XOR2_X1 U367 ( .A(n311), .B(n430), .Z(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U369 ( .A(KEYINPUT36), .B(n577), .Z(n590) );
  XOR2_X1 U370 ( .A(G15GAT), .B(G127GAT), .Z(n444) );
  XNOR2_X1 U371 ( .A(n444), .B(G155GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n316), .B(G211GAT), .ZN(n329) );
  XOR2_X1 U373 ( .A(G57GAT), .B(KEYINPUT13), .Z(n333) );
  XOR2_X1 U374 ( .A(n333), .B(KEYINPUT79), .Z(n318) );
  NAND2_X1 U375 ( .A1(G231GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U377 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n320) );
  XNOR2_X1 U378 ( .A(G22GAT), .B(KEYINPUT14), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U380 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U381 ( .A(G1GAT), .B(G8GAT), .Z(n359) );
  XOR2_X1 U382 ( .A(G78GAT), .B(G64GAT), .Z(n324) );
  XNOR2_X1 U383 ( .A(G183GAT), .B(G71GAT), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n359), .B(n325), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n328) );
  INV_X1 U387 ( .A(n586), .ZN(n466) );
  NOR2_X1 U388 ( .A1(n590), .A2(n466), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n330), .B(KEYINPUT45), .ZN(n346) );
  XOR2_X1 U390 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n332) );
  XNOR2_X1 U391 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n337) );
  XOR2_X1 U393 ( .A(KEYINPUT71), .B(KEYINPUT75), .Z(n335) );
  XNOR2_X1 U394 ( .A(n333), .B(n432), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U396 ( .A(n337), .B(n336), .Z(n339) );
  NAND2_X1 U397 ( .A1(G230GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U399 ( .A(n341), .B(n340), .Z(n345) );
  XNOR2_X1 U400 ( .A(G120GAT), .B(G176GAT), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n342), .B(G71GAT), .ZN(n443) );
  XNOR2_X1 U402 ( .A(G64GAT), .B(KEYINPUT73), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n343), .B(G204GAT), .ZN(n378) );
  XNOR2_X1 U404 ( .A(n443), .B(n378), .ZN(n344) );
  NAND2_X1 U405 ( .A1(n346), .A2(n465), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n347), .B(KEYINPUT117), .ZN(n366) );
  XOR2_X1 U407 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n349) );
  XNOR2_X1 U408 ( .A(KEYINPUT67), .B(KEYINPUT70), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n363) );
  XOR2_X1 U410 ( .A(G113GAT), .B(G36GAT), .Z(n351) );
  XNOR2_X1 U411 ( .A(G43GAT), .B(G50GAT), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U413 ( .A(KEYINPUT30), .B(G15GAT), .Z(n353) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(G197GAT), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U416 ( .A(n355), .B(n354), .Z(n361) );
  XOR2_X1 U417 ( .A(G141GAT), .B(G22GAT), .Z(n427) );
  XOR2_X1 U418 ( .A(n427), .B(KEYINPUT29), .Z(n357) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n365) );
  INV_X1 U424 ( .A(n583), .ZN(n511) );
  NAND2_X1 U425 ( .A1(n583), .A2(n554), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n367), .B(KEYINPUT46), .ZN(n368) );
  XOR2_X1 U427 ( .A(KEYINPUT47), .B(n369), .Z(n370) );
  XOR2_X1 U428 ( .A(KEYINPUT83), .B(G183GAT), .Z(n374) );
  XNOR2_X1 U429 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n376) );
  XOR2_X1 U431 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n375) );
  XOR2_X1 U432 ( .A(n376), .B(n375), .Z(n455) );
  INV_X1 U433 ( .A(n455), .ZN(n392) );
  XNOR2_X1 U434 ( .A(G92GAT), .B(n377), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n385) );
  XOR2_X1 U436 ( .A(G211GAT), .B(KEYINPUT21), .Z(n381) );
  XNOR2_X1 U437 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n433) );
  XOR2_X1 U439 ( .A(n433), .B(G8GAT), .Z(n383) );
  NAND2_X1 U440 ( .A1(G226GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U442 ( .A(n385), .B(n384), .Z(n390) );
  XOR2_X1 U443 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n387) );
  XNOR2_X1 U444 ( .A(G176GAT), .B(KEYINPUT97), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U446 ( .A(G190GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U448 ( .A(n392), .B(n391), .Z(n470) );
  NOR2_X1 U449 ( .A1(n534), .A2(n470), .ZN(n393) );
  XNOR2_X1 U450 ( .A(n394), .B(n393), .ZN(n422) );
  XOR2_X1 U451 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n399) );
  XOR2_X1 U452 ( .A(KEYINPUT88), .B(KEYINPUT2), .Z(n396) );
  XNOR2_X1 U453 ( .A(KEYINPUT89), .B(G155GAT), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U455 ( .A(KEYINPUT3), .B(n397), .Z(n440) );
  XNOR2_X1 U456 ( .A(n440), .B(KEYINPUT92), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U458 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n401) );
  XNOR2_X1 U459 ( .A(G148GAT), .B(KEYINPUT5), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U461 ( .A(n403), .B(n402), .Z(n408) );
  XOR2_X1 U462 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n405) );
  XNOR2_X1 U463 ( .A(G120GAT), .B(KEYINPUT91), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U465 ( .A(G127GAT), .B(n406), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U467 ( .A(KEYINPUT76), .B(G85GAT), .Z(n410) );
  XNOR2_X1 U468 ( .A(G29GAT), .B(G134GAT), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U470 ( .A(n412), .B(n411), .Z(n421) );
  XNOR2_X1 U471 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n413), .B(KEYINPUT80), .ZN(n452) );
  XOR2_X1 U473 ( .A(n452), .B(G141GAT), .Z(n415) );
  NAND2_X1 U474 ( .A1(G225GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U476 ( .A(KEYINPUT4), .B(G57GAT), .Z(n417) );
  XNOR2_X1 U477 ( .A(G1GAT), .B(G162GAT), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U480 ( .A(n421), .B(n420), .Z(n476) );
  INV_X1 U481 ( .A(n476), .ZN(n525) );
  NOR2_X1 U482 ( .A1(n422), .A2(n525), .ZN(n423) );
  XOR2_X1 U483 ( .A(KEYINPUT64), .B(n423), .Z(n564) );
  INV_X1 U484 ( .A(n564), .ZN(n460) );
  XOR2_X1 U485 ( .A(KEYINPUT103), .B(KEYINPUT26), .Z(n458) );
  XOR2_X1 U486 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n425) );
  XNOR2_X1 U487 ( .A(G204GAT), .B(KEYINPUT86), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U489 ( .A(n426), .B(G106GAT), .Z(n429) );
  XNOR2_X1 U490 ( .A(n427), .B(G218GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n431) );
  XOR2_X1 U492 ( .A(n431), .B(n430), .Z(n435) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U495 ( .A(KEYINPUT90), .B(KEYINPUT85), .Z(n437) );
  NAND2_X1 U496 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U498 ( .A(n439), .B(n438), .Z(n442) );
  XNOR2_X1 U499 ( .A(n440), .B(KEYINPUT22), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n563) );
  XOR2_X1 U501 ( .A(n444), .B(n443), .Z(n446) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U504 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n448) );
  XNOR2_X1 U505 ( .A(G99GAT), .B(KEYINPUT81), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U507 ( .A(n450), .B(n449), .Z(n454) );
  XNOR2_X1 U508 ( .A(n451), .B(n452), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n454), .B(n453), .ZN(n456) );
  XOR2_X1 U510 ( .A(n456), .B(n455), .Z(n535) );
  NAND2_X1 U511 ( .A1(n563), .A2(n535), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U513 ( .A(KEYINPUT102), .B(n459), .Z(n472) );
  INV_X1 U514 ( .A(n472), .ZN(n550) );
  NAND2_X1 U515 ( .A1(n460), .A2(n472), .ZN(n589) );
  OR2_X1 U516 ( .A1(n589), .A2(n465), .ZN(n464) );
  XOR2_X1 U517 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n462) );
  XOR2_X1 U518 ( .A(KEYINPUT105), .B(KEYINPUT34), .Z(n485) );
  NAND2_X1 U519 ( .A1(n465), .A2(n583), .ZN(n499) );
  NOR2_X1 U520 ( .A1(n577), .A2(n466), .ZN(n467) );
  XNOR2_X1 U521 ( .A(n467), .B(KEYINPUT16), .ZN(n483) );
  NOR2_X1 U522 ( .A1(n535), .A2(n470), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n563), .A2(n468), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n469), .B(KEYINPUT25), .ZN(n474) );
  INV_X1 U525 ( .A(n470), .ZN(n527) );
  XOR2_X1 U526 ( .A(KEYINPUT27), .B(KEYINPUT100), .Z(n471) );
  XOR2_X1 U527 ( .A(n527), .B(n471), .Z(n478) );
  NAND2_X1 U528 ( .A1(n478), .A2(n472), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U530 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U531 ( .A(KEYINPUT104), .B(n477), .ZN(n482) );
  INV_X1 U532 ( .A(n535), .ZN(n567) );
  XOR2_X1 U533 ( .A(n567), .B(KEYINPUT84), .Z(n479) );
  NAND2_X1 U534 ( .A1(n525), .A2(n478), .ZN(n552) );
  XNOR2_X1 U535 ( .A(n563), .B(KEYINPUT28), .ZN(n531) );
  NOR2_X1 U536 ( .A1(n552), .A2(n531), .ZN(n536) );
  NAND2_X1 U537 ( .A1(n479), .A2(n536), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT101), .B(n480), .Z(n481) );
  NAND2_X1 U539 ( .A1(n482), .A2(n481), .ZN(n496) );
  NAND2_X1 U540 ( .A1(n483), .A2(n496), .ZN(n512) );
  NOR2_X1 U541 ( .A1(n499), .A2(n512), .ZN(n490) );
  NAND2_X1 U542 ( .A1(n490), .A2(n525), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n490), .A2(n527), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT35), .Z(n489) );
  NAND2_X1 U548 ( .A1(n490), .A2(n567), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  NAND2_X1 U550 ( .A1(n531), .A2(n490), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n491), .B(KEYINPUT106), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G22GAT), .B(n492), .ZN(G1327GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT109), .B(KEYINPUT39), .Z(n494) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n502) );
  NOR2_X1 U556 ( .A1(n590), .A2(n586), .ZN(n495) );
  NAND2_X1 U557 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U558 ( .A(KEYINPUT108), .B(n497), .ZN(n498) );
  XOR2_X1 U559 ( .A(KEYINPUT37), .B(n498), .Z(n524) );
  NOR2_X1 U560 ( .A1(n524), .A2(n499), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(KEYINPUT38), .ZN(n508) );
  NAND2_X1 U562 ( .A1(n525), .A2(n508), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(KEYINPUT110), .ZN(n504) );
  NAND2_X1 U565 ( .A1(n527), .A2(n508), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(G1329GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT40), .B(KEYINPUT111), .Z(n506) );
  NAND2_X1 U568 ( .A1(n508), .A2(n567), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NAND2_X1 U571 ( .A1(n508), .A2(n531), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n509), .B(KEYINPUT112), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(n510), .ZN(G1331GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT114), .B(KEYINPUT42), .Z(n514) );
  XOR2_X1 U575 ( .A(KEYINPUT113), .B(n554), .Z(n571) );
  NAND2_X1 U576 ( .A1(n511), .A2(n571), .ZN(n523) );
  NOR2_X1 U577 ( .A1(n523), .A2(n512), .ZN(n519) );
  NAND2_X1 U578 ( .A1(n519), .A2(n525), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U580 ( .A(G57GAT), .B(n515), .Z(G1332GAT) );
  XOR2_X1 U581 ( .A(G64GAT), .B(KEYINPUT115), .Z(n517) );
  NAND2_X1 U582 ( .A1(n519), .A2(n527), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1333GAT) );
  NAND2_X1 U584 ( .A1(n567), .A2(n519), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n518), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT116), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U587 ( .A1(n519), .A2(n531), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(n522), .ZN(G1335GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n530) );
  NAND2_X1 U591 ( .A1(n525), .A2(n530), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n567), .A2(n530), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  XOR2_X1 U600 ( .A(G113GAT), .B(KEYINPUT119), .Z(n540) );
  NOR2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n537) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U603 ( .A(KEYINPUT118), .B(n538), .Z(n547) );
  NAND2_X1 U604 ( .A1(n547), .A2(n583), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT120), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U607 ( .A1(n547), .A2(n571), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(KEYINPUT121), .Z(n545) );
  NAND2_X1 U611 ( .A1(n586), .A2(n547), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U615 ( .A1(n577), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  OR2_X1 U617 ( .A1(n534), .A2(n550), .ZN(n551) );
  NOR2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n559), .A2(n583), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U622 ( .A1(n559), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n586), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT122), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(n562), .ZN(G1347GAT) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n570) );
  XNOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT55), .ZN(n566) );
  NOR2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n576), .A2(n583), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1348GAT) );
  NAND2_X1 U636 ( .A1(n576), .A2(n571), .ZN(n573) );
  XOR2_X1 U637 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G176GAT), .B(n574), .ZN(G1349GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n586), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT58), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U648 ( .A(KEYINPUT125), .B(n582), .Z(n585) );
  INV_X1 U649 ( .A(n589), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n587), .A2(n583), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

