//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(G137), .A3(new_n460), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT69), .B1(new_n466), .B2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(new_n460), .A3(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  OR2_X1    g046(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n460), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT70), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n461), .A2(new_n460), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AND3_X1   g058(.A1(new_n478), .A2(new_n480), .A3(new_n483), .ZN(G162));
  AND2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI211_X1 g061(.A(G138), .B(new_n460), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n461), .A2(KEYINPUT72), .A3(G138), .A4(new_n460), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(new_n460), .B2(G114), .ZN(new_n493));
  NOR2_X1   g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n494), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT71), .A4(G2104), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n495), .A2(new_n499), .B1(new_n476), .B2(G126), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n487), .A2(new_n488), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n491), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT73), .A3(G62), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(new_n508), .ZN(new_n513));
  INV_X1    g088(.A(G62), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n510), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n509), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n517), .A2(new_n527), .ZN(G166));
  AND2_X1   g103(.A1(new_n509), .A2(new_n522), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n522), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n530), .A2(new_n532), .A3(new_n533), .A4(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n523), .A2(new_n538), .B1(new_n525), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT74), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n518), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n541), .A2(KEYINPUT75), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(KEYINPUT75), .B1(new_n541), .B2(new_n543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n523), .A2(new_n548), .B1(new_n525), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n509), .A2(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n518), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT76), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n513), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n529), .A2(G91), .B1(new_n564), .B2(G651), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n519), .A2(new_n521), .A3(G53), .A4(G543), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND2_X1  g144(.A1(new_n529), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n531), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n513), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT77), .ZN(new_n578));
  AOI22_X1  g153(.A1(G86), .A2(new_n529), .B1(new_n531), .B2(G48), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G305));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n523), .A2(new_n581), .B1(new_n525), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n518), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  AND3_X1   g162(.A1(new_n509), .A2(new_n522), .A3(G92), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n531), .A2(G54), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(new_n518), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G171), .B2(new_n594), .ZN(G321));
  XOR2_X1   g171(.A(G321), .B(KEYINPUT78), .Z(G284));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G299), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G297));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G280));
  INV_X1    g176(.A(new_n593), .ZN(new_n602));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n467), .A2(new_n469), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(new_n461), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(G2100), .ZN(new_n616));
  AOI21_X1  g191(.A(KEYINPUT79), .B1(new_n482), .B2(G135), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(G123), .B2(new_n476), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n482), .A2(KEYINPUT79), .A3(G135), .ZN(new_n619));
  NOR2_X1   g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(new_n460), .B2(G111), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2096), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n615), .A2(new_n616), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT80), .Z(G156));
  XNOR2_X1  g201(.A(KEYINPUT82), .B(G1341), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2435), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2438), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G1348), .ZN(new_n634));
  INV_X1    g209(.A(G1348), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n634), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n638), .B1(new_n634), .B2(new_n636), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n628), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n634), .A2(new_n636), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(new_n637), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n634), .A2(new_n636), .A3(new_n638), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n627), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n647), .B(new_n648), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n641), .A2(new_n645), .A3(new_n649), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT83), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT84), .Z(G401));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2067), .B(G2678), .Z(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(KEYINPUT18), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n623), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n661), .A2(new_n664), .A3(KEYINPUT17), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT86), .B(G2100), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n673), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  AOI22_X1  g254(.A1(new_n677), .A2(KEYINPUT20), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n679), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n681), .A2(new_n673), .A3(new_n676), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n680), .B(new_n682), .C1(KEYINPUT20), .C2(new_n677), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT87), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G25), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n482), .A2(G131), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n476), .A2(G119), .ZN(new_n695));
  OR2_X1    g270(.A1(G95), .A2(G2105), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n696), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n693), .B1(new_n699), .B2(new_n692), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G1986), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n586), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n704), .B2(G24), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n702), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n709));
  XNOR2_X1  g284(.A(G288), .B(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n708), .B1(new_n710), .B2(new_n704), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G6), .B(G305), .S(G16), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n704), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n704), .ZN(new_n718));
  INV_X1    g293(.A(G1971), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n713), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n707), .B1(new_n721), .B2(KEYINPUT34), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(KEYINPUT34), .B2(new_n721), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n703), .B2(new_n706), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT36), .Z(new_n725));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G4), .B2(G16), .ZN(new_n727));
  OR3_X1    g302(.A1(new_n726), .A2(G4), .A3(G16), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n727), .B(new_n728), .C1(new_n593), .C2(new_n704), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(new_n635), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT90), .B(KEYINPUT91), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G5), .A2(G16), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G171), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G164), .A2(new_n692), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G27), .B2(new_n692), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT96), .B(G2078), .Z(new_n739));
  OAI21_X1  g314(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(KEYINPUT24), .A2(G34), .ZN(new_n741));
  NOR2_X1   g316(.A1(KEYINPUT24), .A2(G34), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n692), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT93), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n472), .B2(new_n692), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n744), .B2(new_n743), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G2084), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n692), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n692), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT29), .B(G2090), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT31), .B(G11), .Z(new_n753));
  NOR2_X1   g328(.A1(new_n622), .A2(new_n692), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n692), .A2(G33), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n482), .A2(G139), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT25), .Z(new_n758));
  AOI22_X1  g333(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n756), .B(new_n758), .C1(new_n460), .C2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n755), .B1(new_n760), .B2(G29), .ZN(new_n761));
  INV_X1    g336(.A(G2072), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n692), .B1(new_n764), .B2(G28), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n764), .B2(G28), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n754), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n762), .B2(new_n761), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n752), .A2(new_n753), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n704), .A2(G19), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n555), .B2(new_n704), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT92), .B(G1341), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n738), .A2(new_n739), .B1(new_n750), .B2(new_n751), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n769), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G29), .A2(G32), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n482), .A2(G141), .B1(G129), .B2(new_n476), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n610), .A2(G105), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT94), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT26), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n776), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT27), .B(G1996), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G286), .A2(new_n704), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT95), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(KEYINPUT95), .B1(G16), .B2(G21), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G1966), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT28), .ZN(new_n794));
  INV_X1    g369(.A(G26), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G29), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(G29), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n476), .A2(G128), .ZN(new_n798));
  NOR2_X1   g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(new_n460), .B2(G116), .ZN(new_n800));
  INV_X1    g375(.A(G140), .ZN(new_n801));
  OAI221_X1 g376(.A(new_n798), .B1(new_n799), .B2(new_n800), .C1(new_n801), .C2(new_n481), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n797), .B1(new_n802), .B2(G29), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(new_n794), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n792), .A2(G1966), .B1(G2067), .B2(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(G2067), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n704), .A2(G20), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT97), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT23), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G299), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1956), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n793), .A2(new_n805), .A3(new_n806), .A4(new_n811), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n740), .A2(new_n775), .A3(new_n787), .A4(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n725), .A2(new_n732), .A3(new_n813), .ZN(G150));
  INV_X1    g389(.A(G150), .ZN(G311));
  NAND2_X1  g390(.A1(new_n529), .A2(G93), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT99), .B(G55), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n816), .B1(new_n518), .B2(new_n817), .C1(new_n525), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G860), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT100), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT37), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n819), .A2(new_n554), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n555), .B2(new_n819), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n593), .A2(new_n603), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT39), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n822), .B1(new_n829), .B2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT101), .Z(G145));
  XNOR2_X1  g406(.A(G162), .B(KEYINPUT102), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G160), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n622), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n476), .A2(G130), .ZN(new_n836));
  NOR2_X1   g411(.A1(G106), .A2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(new_n460), .B2(G118), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G142), .B2(new_n482), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n698), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT104), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n612), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n783), .B(new_n503), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT103), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n760), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n802), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n844), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n843), .A2(new_n848), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n835), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n843), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n848), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n851), .B(new_n852), .C1(new_n855), .C2(new_n835), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g432(.A1(new_n710), .A2(G290), .ZN(new_n858));
  XNOR2_X1  g433(.A(G288), .B(KEYINPUT88), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n586), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(G305), .A2(G166), .ZN(new_n862));
  NAND2_X1  g437(.A1(G305), .A2(G166), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT108), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n861), .A2(KEYINPUT108), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n858), .A2(new_n860), .A3(new_n862), .A4(new_n863), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT107), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n870), .A2(KEYINPUT107), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(KEYINPUT109), .A3(KEYINPUT42), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n870), .B(KEYINPUT107), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n867), .A3(new_n868), .ZN(new_n876));
  OR2_X1    g451(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n877));
  NAND2_X1  g452(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n824), .B(new_n605), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n593), .B(G299), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT41), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n882), .B(KEYINPUT106), .Z(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n885), .B2(new_n881), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT110), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n880), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n874), .A2(new_n887), .A3(new_n879), .A4(new_n886), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(G868), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n819), .A2(new_n594), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  MUX2_X1   g469(.A(new_n892), .B(new_n894), .S(KEYINPUT111), .Z(G295));
  MUX2_X1   g470(.A(new_n892), .B(new_n894), .S(KEYINPUT111), .Z(G331));
  INV_X1    g471(.A(new_n824), .ZN(new_n897));
  OAI21_X1  g472(.A(G168), .B1(new_n544), .B2(new_n545), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n544), .A2(new_n545), .A3(G168), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n824), .A3(new_n898), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n903), .A3(new_n883), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n903), .ZN(new_n905));
  INV_X1    g480(.A(new_n882), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n876), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT112), .B1(new_n908), .B2(G37), .ZN(new_n909));
  INV_X1    g484(.A(new_n904), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n882), .B1(new_n901), .B2(new_n903), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n873), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT112), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n913), .A3(new_n852), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(new_n876), .A3(new_n904), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n885), .B1(new_n901), .B2(new_n903), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n873), .B1(new_n919), .B2(new_n910), .ZN(new_n920));
  AND4_X1   g495(.A1(KEYINPUT43), .A2(new_n920), .A3(new_n852), .A4(new_n915), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT44), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n920), .A2(new_n917), .A3(new_n852), .A4(new_n915), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n922), .A2(new_n927), .ZN(G397));
  XNOR2_X1  g503(.A(KEYINPUT113), .B(G1384), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n503), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n931));
  INV_X1    g506(.A(G40), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n464), .A2(new_n471), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(G290), .A2(G1986), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT48), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n934), .A2(G1996), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n784), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n939), .B(KEYINPUT114), .Z(new_n940));
  INV_X1    g515(.A(G2067), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n802), .B(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G1996), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n784), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n940), .B1(new_n935), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n698), .B(new_n701), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(new_n934), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT125), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n937), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n935), .A2(KEYINPUT48), .A3(new_n936), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n949), .B(new_n950), .C1(new_n948), .C2(new_n947), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n938), .A2(KEYINPUT46), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n938), .A2(KEYINPUT46), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n934), .B1(new_n784), .B2(new_n942), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT47), .Z(new_n956));
  NAND3_X1  g531(.A1(new_n945), .A2(new_n701), .A3(new_n699), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G2067), .B2(new_n802), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n935), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n951), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n936), .ZN(new_n961));
  NAND2_X1  g536(.A1(G290), .A2(G1986), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n934), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n947), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n503), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT115), .B1(new_n966), .B2(new_n931), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n968), .B(KEYINPUT45), .C1(new_n503), .C2(new_n965), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n971), .A2(new_n933), .ZN(new_n972));
  AOI21_X1  g547(.A(G1971), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n503), .B2(new_n965), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G2090), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n503), .A2(new_n965), .A3(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n977), .A2(new_n978), .A3(new_n933), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT117), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n982), .A2(KEYINPUT117), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n974), .A2(KEYINPUT118), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT118), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n982), .B(KEYINPUT117), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(new_n987), .B2(new_n973), .ZN(new_n988));
  INV_X1    g563(.A(G8), .ZN(new_n989));
  NOR2_X1   g564(.A1(G166), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n990), .B(KEYINPUT55), .Z(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n985), .A2(new_n988), .A3(G8), .A4(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(G305), .A2(G1981), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n579), .A2(new_n577), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G1981), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n933), .A2(new_n503), .A3(new_n965), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n994), .A2(KEYINPUT49), .A3(new_n996), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n999), .A2(G8), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(G8), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n710), .B2(G1976), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G288), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1004), .B(new_n1005), .C1(G1976), .C2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n993), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1976), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1002), .A2(new_n1011), .A3(new_n1007), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1003), .B1(new_n1012), .B2(new_n994), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT56), .B(G2072), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n972), .B(new_n1016), .C1(new_n967), .C2(new_n969), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n565), .A2(new_n1019), .A3(new_n567), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1019), .B1(new_n565), .B2(new_n567), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1018), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1022), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(KEYINPUT57), .A3(new_n1020), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1956), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n933), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n980), .B1(new_n503), .B2(new_n965), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1017), .A2(new_n1026), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1026), .B1(new_n1017), .B2(new_n1030), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n981), .A2(new_n933), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n635), .B1(new_n1033), .B2(new_n976), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1000), .A2(KEYINPUT121), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n933), .A2(new_n503), .A3(new_n1036), .A4(new_n965), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n941), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n593), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1031), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1017), .A2(new_n1030), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1026), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT61), .A3(new_n1031), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n972), .B(new_n943), .C1(new_n967), .C2(new_n969), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1047));
  XOR2_X1   g622(.A(KEYINPUT58), .B(G1341), .Z(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1045), .B1(new_n1050), .B2(new_n555), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1050), .A2(new_n1045), .A3(new_n555), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1044), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT61), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1017), .A2(new_n1026), .A3(new_n1030), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(new_n1055), .B2(new_n1032), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT60), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n593), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1034), .A2(new_n1038), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n602), .A2(KEYINPUT60), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1040), .B1(new_n1053), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G2078), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n972), .B(new_n1064), .C1(new_n967), .C2(new_n969), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n977), .A2(new_n933), .A3(new_n981), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n735), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1064), .A2(KEYINPUT53), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n930), .B2(new_n931), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n972), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1067), .A2(G301), .A3(new_n1069), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT122), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n966), .A2(new_n931), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n933), .A3(new_n1076), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1077), .A2(new_n1070), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1067), .A2(new_n1069), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G171), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1065), .A2(new_n1066), .B1(new_n735), .B2(new_n1068), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(G301), .A4(new_n1072), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1074), .A2(new_n1080), .A3(new_n1081), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1079), .A2(G301), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(G171), .A3(new_n1072), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(KEYINPUT54), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G286), .A2(G8), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1033), .A2(new_n976), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT119), .B(G2084), .Z(new_n1093));
  INV_X1    g668(.A(G1966), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1092), .A2(new_n1093), .B1(new_n1077), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1090), .B(new_n1091), .C1(new_n1095), .C2(new_n989), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1077), .A2(new_n1094), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n977), .A2(new_n933), .A3(new_n981), .A4(new_n1093), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT51), .B(G8), .C1(new_n1099), .C2(G286), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1095), .A2(new_n1091), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1063), .A2(new_n1089), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1102), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1080), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1106), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1105), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1009), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n993), .A2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1028), .A2(G2090), .A3(new_n1029), .ZN(new_n1116));
  OAI21_X1  g691(.A(G8), .B1(new_n973), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n991), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1015), .B1(new_n1113), .B2(new_n1119), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1095), .A2(new_n989), .A3(G286), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n985), .A2(new_n988), .A3(G8), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(new_n991), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1115), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n993), .A2(new_n1114), .A3(new_n1118), .A4(new_n1121), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1122), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g703(.A(KEYINPUT124), .B(new_n964), .C1(new_n1120), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(new_n1014), .A3(new_n1128), .ZN(new_n1132));
  INV_X1    g707(.A(new_n964), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n960), .B1(new_n1129), .B2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g710(.A(KEYINPUT83), .ZN(new_n1137));
  AND3_X1   g711(.A1(new_n641), .A2(new_n645), .A3(new_n649), .ZN(new_n1138));
  AOI21_X1  g712(.A(new_n649), .B1(new_n641), .B2(new_n645), .ZN(new_n1139));
  NOR2_X1   g713(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1140), .B2(G14), .ZN(new_n1141));
  NOR2_X1   g715(.A1(new_n653), .A2(KEYINPUT83), .ZN(new_n1142));
  OAI211_X1 g716(.A(G319), .B(new_n670), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g717(.A1(new_n1143), .A2(KEYINPUT126), .ZN(new_n1144));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n1145));
  NAND4_X1  g719(.A1(new_n654), .A2(new_n1145), .A3(G319), .A4(new_n670), .ZN(new_n1146));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n1146), .A3(new_n690), .ZN(new_n1147));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n1148));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g723(.A1(new_n1144), .A2(new_n1146), .A3(KEYINPUT127), .A4(new_n690), .ZN(new_n1150));
  AND4_X1   g724(.A1(new_n856), .A2(new_n1149), .A3(new_n925), .A4(new_n1150), .ZN(G308));
  NAND4_X1  g725(.A1(new_n1149), .A2(new_n925), .A3(new_n856), .A4(new_n1150), .ZN(G225));
endmodule


