

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747;

  NAND2_X1 U366 ( .A1(n439), .A2(n438), .ZN(n603) );
  INV_X2 U367 ( .A(n524), .ZN(n429) );
  XNOR2_X2 U368 ( .A(n523), .B(n522), .ZN(n524) );
  OR2_X2 U369 ( .A1(n706), .A2(G902), .ZN(n496) );
  NOR2_X2 U370 ( .A1(n418), .A2(n414), .ZN(n455) );
  AND2_X2 U371 ( .A1(n525), .A2(n433), .ZN(n432) );
  XNOR2_X2 U372 ( .A(n520), .B(n519), .ZN(n634) );
  XOR2_X2 U373 ( .A(KEYINPUT76), .B(n511), .Z(n525) );
  NOR2_X2 U374 ( .A1(n594), .A2(n541), .ZN(n511) );
  XNOR2_X2 U375 ( .A(n413), .B(G125), .ZN(n530) );
  AND2_X1 U376 ( .A1(n604), .A2(n670), .ZN(n390) );
  INV_X2 U377 ( .A(G143), .ZN(n406) );
  AND2_X1 U378 ( .A1(n404), .A2(n402), .ZN(n400) );
  NAND2_X1 U379 ( .A1(n670), .A2(n562), .ZN(n594) );
  NOR2_X1 U380 ( .A1(n447), .A2(KEYINPUT6), .ZN(n385) );
  INV_X1 U381 ( .A(n598), .ZN(n345) );
  NAND2_X1 U382 ( .A1(n400), .A2(n399), .ZN(n398) );
  NAND2_X1 U383 ( .A1(n401), .A2(n635), .ZN(n399) );
  AND2_X1 U384 ( .A1(n372), .A2(n371), .ZN(n370) );
  XNOR2_X1 U385 ( .A(n453), .B(n452), .ZN(n745) );
  NAND2_X1 U386 ( .A1(n431), .A2(n430), .ZN(n453) );
  OR2_X1 U387 ( .A1(n525), .A2(n424), .ZN(n430) );
  XNOR2_X1 U388 ( .A(n381), .B(n380), .ZN(n698) );
  XNOR2_X1 U389 ( .A(n409), .B(n510), .ZN(n598) );
  INV_X1 U390 ( .A(G146), .ZN(n413) );
  NAND2_X1 U391 ( .A1(n624), .A2(n623), .ZN(n443) );
  OR2_X2 U392 ( .A1(n743), .A2(KEYINPUT44), .ZN(n616) );
  XNOR2_X2 U393 ( .A(n550), .B(KEYINPUT86), .ZN(n559) );
  XNOR2_X2 U394 ( .A(n731), .B(n450), .ZN(n520) );
  XNOR2_X2 U395 ( .A(n451), .B(n491), .ZN(n731) );
  OR2_X1 U396 ( .A1(n634), .A2(n446), .ZN(n445) );
  NOR2_X1 U397 ( .A1(n636), .A2(KEYINPUT84), .ZN(n373) );
  NOR2_X1 U398 ( .A1(KEYINPUT71), .A2(KEYINPUT44), .ZN(n612) );
  NOR2_X1 U399 ( .A1(n445), .A2(KEYINPUT6), .ZN(n389) );
  INV_X1 U400 ( .A(KEYINPUT4), .ZN(n488) );
  XOR2_X1 U401 ( .A(KEYINPUT88), .B(n497), .Z(n619) );
  XNOR2_X1 U402 ( .A(n378), .B(KEYINPUT15), .ZN(n497) );
  INV_X1 U403 ( .A(G902), .ZN(n378) );
  OR2_X1 U404 ( .A1(G237), .A2(G902), .ZN(n537) );
  NAND2_X1 U405 ( .A1(n568), .A2(n358), .ZN(n405) );
  INV_X1 U406 ( .A(KEYINPUT48), .ZN(n421) );
  NOR2_X1 U407 ( .A1(n369), .A2(n349), .ZN(n368) );
  NAND2_X1 U408 ( .A1(n374), .A2(n373), .ZN(n371) );
  NOR2_X1 U409 ( .A1(G953), .A2(G237), .ZN(n470) );
  XNOR2_X1 U410 ( .A(G113), .B(G143), .ZN(n471) );
  XOR2_X1 U411 ( .A(G104), .B(G122), .Z(n472) );
  INV_X1 U412 ( .A(G146), .ZN(n450) );
  NOR2_X1 U413 ( .A1(n715), .A2(G902), .ZN(n409) );
  XNOR2_X1 U414 ( .A(n477), .B(n476), .ZN(n478) );
  NOR2_X1 U415 ( .A1(n389), .A2(n385), .ZN(n387) );
  AND2_X1 U416 ( .A1(n445), .A2(KEYINPUT6), .ZN(n388) );
  XNOR2_X1 U417 ( .A(n500), .B(n352), .ZN(n411) );
  XOR2_X1 U418 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n466) );
  XNOR2_X1 U419 ( .A(n530), .B(G140), .ZN(n412) );
  XNOR2_X1 U420 ( .A(n459), .B(n353), .ZN(n382) );
  AND2_X1 U421 ( .A1(n628), .A2(G210), .ZN(n417) );
  INV_X1 U422 ( .A(KEYINPUT1), .ZN(n407) );
  NAND2_X1 U423 ( .A1(n426), .A2(n350), .ZN(n425) );
  NAND2_X1 U424 ( .A1(n524), .A2(n433), .ZN(n426) );
  OR2_X1 U425 ( .A1(n683), .A2(KEYINPUT39), .ZN(n428) );
  XNOR2_X1 U426 ( .A(n556), .B(KEYINPUT107), .ZN(n611) );
  XNOR2_X1 U427 ( .A(n465), .B(n464), .ZN(n566) );
  INV_X1 U428 ( .A(n397), .ZN(n394) );
  AND2_X1 U429 ( .A1(n665), .A2(G475), .ZN(n442) );
  XNOR2_X1 U430 ( .A(n498), .B(KEYINPUT20), .ZN(n507) );
  NAND2_X1 U431 ( .A1(n619), .A2(G234), .ZN(n498) );
  XOR2_X1 U432 ( .A(KEYINPUT18), .B(KEYINPUT87), .Z(n534) );
  XNOR2_X1 U433 ( .A(G116), .B(G101), .ZN(n515) );
  XNOR2_X1 U434 ( .A(n532), .B(G137), .ZN(n451) );
  NAND2_X1 U435 ( .A1(G234), .A2(G237), .ZN(n481) );
  XNOR2_X1 U436 ( .A(n539), .B(n538), .ZN(n549) );
  OR2_X1 U437 ( .A1(n351), .A2(G902), .ZN(n446) );
  NAND2_X1 U438 ( .A1(n351), .A2(G902), .ZN(n448) );
  AND2_X1 U439 ( .A1(n600), .A2(n383), .ZN(n438) );
  AND2_X1 U440 ( .A1(n420), .A2(n419), .ZN(n577) );
  INV_X1 U441 ( .A(n746), .ZN(n419) );
  XNOR2_X1 U442 ( .A(n422), .B(n421), .ZN(n420) );
  XNOR2_X1 U443 ( .A(n513), .B(G119), .ZN(n527) );
  XNOR2_X1 U444 ( .A(n376), .B(n363), .ZN(n725) );
  INV_X1 U445 ( .A(KEYINPUT45), .ZN(n618) );
  XNOR2_X1 U446 ( .A(n475), .B(n474), .ZN(n632) );
  XNOR2_X1 U447 ( .A(n473), .B(n354), .ZN(n474) );
  INV_X1 U448 ( .A(KEYINPUT41), .ZN(n380) );
  NAND2_X1 U449 ( .A1(n690), .A2(n571), .ZN(n381) );
  NOR2_X1 U450 ( .A1(n403), .A2(n717), .ZN(n402) );
  NOR2_X1 U451 ( .A1(n454), .A2(G472), .ZN(n403) );
  XNOR2_X1 U452 ( .A(G101), .B(G110), .ZN(n492) );
  XNOR2_X1 U453 ( .A(n367), .B(n527), .ZN(n719) );
  XNOR2_X1 U454 ( .A(n526), .B(KEYINPUT16), .ZN(n367) );
  XNOR2_X1 U455 ( .A(n506), .B(n505), .ZN(n715) );
  XNOR2_X1 U456 ( .A(n732), .B(n410), .ZN(n506) );
  XNOR2_X1 U457 ( .A(n411), .B(n503), .ZN(n410) );
  XNOR2_X1 U458 ( .A(n461), .B(n382), .ZN(n462) );
  NAND2_X1 U459 ( .A1(n713), .A2(n417), .ZN(n416) );
  INV_X1 U460 ( .A(KEYINPUT40), .ZN(n452) );
  NAND2_X1 U461 ( .A1(n347), .A2(n396), .ZN(n395) );
  AND2_X1 U462 ( .A1(n610), .A2(n435), .ZN(n646) );
  AND2_X1 U463 ( .A1(n611), .A2(n436), .ZN(n435) );
  INV_X1 U464 ( .A(n345), .ZN(n436) );
  XNOR2_X1 U465 ( .A(n480), .B(KEYINPUT105), .ZN(n655) );
  NAND2_X1 U466 ( .A1(n394), .A2(n396), .ZN(n393) );
  XNOR2_X1 U467 ( .A(n377), .B(n364), .ZN(G60) );
  XNOR2_X1 U468 ( .A(n392), .B(n709), .ZN(n391) );
  NAND2_X1 U469 ( .A1(n713), .A2(G469), .ZN(n392) );
  AND2_X1 U470 ( .A1(n683), .A2(KEYINPUT39), .ZN(n346) );
  AND2_X1 U471 ( .A1(n666), .A2(n397), .ZN(n347) );
  NAND2_X2 U472 ( .A1(n387), .A2(n386), .ZN(n604) );
  NOR2_X1 U473 ( .A1(n432), .A2(n359), .ZN(n348) );
  AND2_X1 U474 ( .A1(n608), .A2(KEYINPUT84), .ZN(n349) );
  AND2_X1 U475 ( .A1(n428), .A2(n427), .ZN(n350) );
  XNOR2_X1 U476 ( .A(G472), .B(KEYINPUT72), .ZN(n351) );
  XOR2_X1 U477 ( .A(G128), .B(G110), .Z(n352) );
  XOR2_X1 U478 ( .A(n458), .B(n457), .Z(n353) );
  XOR2_X1 U479 ( .A(n472), .B(n471), .Z(n354) );
  XOR2_X2 U480 ( .A(G104), .B(G107), .Z(n355) );
  NOR2_X1 U481 ( .A1(n525), .A2(n524), .ZN(n356) );
  AND2_X1 U482 ( .A1(n669), .A2(n670), .ZN(n357) );
  XNOR2_X1 U483 ( .A(KEYINPUT82), .B(n660), .ZN(n358) );
  AND2_X1 U484 ( .A1(n434), .A2(n433), .ZN(n359) );
  AND2_X1 U485 ( .A1(n454), .A2(G472), .ZN(n360) );
  INV_X1 U486 ( .A(KEYINPUT39), .ZN(n433) );
  AND2_X1 U487 ( .A1(n415), .A2(n629), .ZN(n361) );
  INV_X1 U488 ( .A(n653), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n632), .B(KEYINPUT59), .ZN(n362) );
  XOR2_X1 U490 ( .A(n618), .B(KEYINPUT65), .Z(n363) );
  NOR2_X1 U491 ( .A1(n739), .A2(G952), .ZN(n717) );
  XOR2_X1 U492 ( .A(n633), .B(KEYINPUT60), .Z(n364) );
  XNOR2_X1 U493 ( .A(n366), .B(n365), .ZN(n625) );
  XNOR2_X1 U494 ( .A(n535), .B(n719), .ZN(n365) );
  XNOR2_X1 U495 ( .A(n536), .B(n528), .ZN(n366) );
  XNOR2_X2 U496 ( .A(n718), .B(KEYINPUT70), .ZN(n528) );
  XNOR2_X2 U497 ( .A(n355), .B(n492), .ZN(n718) );
  NAND2_X1 U498 ( .A1(n370), .A2(n368), .ZN(n376) );
  NAND2_X1 U499 ( .A1(n617), .A2(n375), .ZN(n369) );
  NAND2_X1 U500 ( .A1(n615), .A2(n614), .ZN(n372) );
  INV_X1 U501 ( .A(n608), .ZN(n374) );
  NAND2_X1 U502 ( .A1(n636), .A2(KEYINPUT84), .ZN(n375) );
  NAND2_X1 U503 ( .A1(n379), .A2(n629), .ZN(n377) );
  AND2_X1 U504 ( .A1(n391), .A2(n629), .ZN(G54) );
  XNOR2_X1 U505 ( .A(n444), .B(n362), .ZN(n379) );
  NAND2_X1 U506 ( .A1(n713), .A2(n360), .ZN(n404) );
  NOR2_X2 U507 ( .A1(n607), .A2(n666), .ZN(n636) );
  NOR2_X2 U508 ( .A1(n609), .A2(n395), .ZN(n437) );
  XNOR2_X2 U509 ( .A(n603), .B(n602), .ZN(n609) );
  NAND2_X1 U510 ( .A1(n345), .A2(n383), .ZN(n408) );
  INV_X1 U511 ( .A(n667), .ZN(n383) );
  OR2_X1 U512 ( .A1(n599), .A2(n556), .ZN(n593) );
  XNOR2_X2 U513 ( .A(n440), .B(KEYINPUT0), .ZN(n599) );
  NAND2_X1 U514 ( .A1(n507), .A2(G221), .ZN(n499) );
  NAND2_X1 U515 ( .A1(n388), .A2(n447), .ZN(n386) );
  NOR2_X2 U516 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U517 ( .A1(n384), .A2(n684), .ZN(n596) );
  NAND2_X1 U518 ( .A1(n640), .A2(n656), .ZN(n384) );
  NAND2_X1 U519 ( .A1(n634), .A2(n351), .ZN(n449) );
  NAND2_X2 U520 ( .A1(n447), .A2(n445), .ZN(n556) );
  NAND2_X1 U521 ( .A1(n669), .A2(n390), .ZN(n586) );
  AND2_X4 U522 ( .A1(n443), .A2(n665), .ZN(n713) );
  NOR2_X1 U523 ( .A1(n609), .A2(n393), .ZN(n606) );
  INV_X1 U524 ( .A(n604), .ZN(n396) );
  INV_X1 U525 ( .A(n605), .ZN(n397) );
  XNOR2_X1 U526 ( .A(n398), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U527 ( .A(n713), .ZN(n401) );
  NAND2_X1 U528 ( .A1(n357), .A2(n556), .ZN(n678) );
  XNOR2_X1 U529 ( .A(n532), .B(n531), .ZN(n536) );
  NOR2_X1 U530 ( .A1(n564), .A2(n405), .ZN(n569) );
  XNOR2_X2 U531 ( .A(KEYINPUT79), .B(n553), .ZN(n651) );
  OR2_X2 U532 ( .A1(n584), .A2(n583), .ZN(n440) );
  INV_X2 U533 ( .A(G116), .ZN(n441) );
  NAND2_X1 U534 ( .A1(n662), .A2(n620), .ZN(n624) );
  NOR2_X2 U535 ( .A1(n725), .A2(n737), .ZN(n662) );
  NAND2_X1 U536 ( .A1(n443), .A2(n442), .ZN(n444) );
  XNOR2_X2 U537 ( .A(n489), .B(n488), .ZN(n532) );
  XNOR2_X2 U538 ( .A(n406), .B(G128), .ZN(n489) );
  XNOR2_X2 U539 ( .A(n562), .B(n407), .ZN(n605) );
  XNOR2_X2 U540 ( .A(n496), .B(G469), .ZN(n562) );
  XNOR2_X2 U541 ( .A(n408), .B(KEYINPUT67), .ZN(n670) );
  XNOR2_X2 U542 ( .A(n412), .B(n466), .ZN(n732) );
  NAND2_X1 U543 ( .A1(n416), .A2(n361), .ZN(n414) );
  OR2_X1 U544 ( .A1(n628), .A2(G210), .ZN(n415) );
  NOR2_X1 U545 ( .A1(n713), .A2(n628), .ZN(n418) );
  NAND2_X1 U546 ( .A1(n423), .A2(n569), .ZN(n422) );
  XNOR2_X1 U547 ( .A(n548), .B(KEYINPUT46), .ZN(n423) );
  NAND2_X1 U548 ( .A1(n429), .A2(n683), .ZN(n434) );
  NAND2_X1 U549 ( .A1(n429), .A2(n346), .ZN(n424) );
  NOR2_X1 U550 ( .A1(n425), .A2(n432), .ZN(n431) );
  NAND2_X1 U551 ( .A1(n348), .A2(n430), .ZN(n547) );
  XNOR2_X1 U552 ( .A(n613), .B(n612), .ZN(n615) );
  NOR2_X2 U553 ( .A1(n744), .A2(n646), .ZN(n613) );
  XNOR2_X2 U554 ( .A(n437), .B(KEYINPUT32), .ZN(n744) );
  INV_X1 U555 ( .A(n599), .ZN(n439) );
  XNOR2_X2 U556 ( .A(n441), .B(G122), .ZN(n526) );
  AND2_X2 U557 ( .A1(n449), .A2(n448), .ZN(n447) );
  NOR2_X1 U558 ( .A1(n611), .A2(n687), .ZN(n523) );
  NOR2_X1 U559 ( .A1(n745), .A2(n747), .ZN(n548) );
  INV_X1 U560 ( .A(n635), .ZN(n454) );
  XNOR2_X1 U561 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U562 ( .A(n514), .B(n527), .ZN(n518) );
  INV_X1 U563 ( .A(KEYINPUT95), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n503) );
  INV_X1 U566 ( .A(G475), .ZN(n476) );
  XNOR2_X1 U567 ( .A(n601), .B(KEYINPUT22), .ZN(n602) );
  XNOR2_X1 U568 ( .A(n479), .B(n478), .ZN(n565) );
  INV_X1 U569 ( .A(n655), .ZN(n647) );
  XNOR2_X1 U570 ( .A(KEYINPUT104), .B(G478), .ZN(n465) );
  XNOR2_X1 U571 ( .A(n526), .B(G134), .ZN(n463) );
  XNOR2_X1 U572 ( .A(n489), .B(G107), .ZN(n456) );
  XNOR2_X1 U573 ( .A(n456), .B(KEYINPUT101), .ZN(n459) );
  XOR2_X1 U574 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n458) );
  XNOR2_X1 U575 ( .A(KEYINPUT103), .B(KEYINPUT9), .ZN(n457) );
  XNOR2_X1 U576 ( .A(KEYINPUT64), .B(G953), .ZN(n484) );
  INV_X1 U577 ( .A(n484), .ZN(n739) );
  NAND2_X1 U578 ( .A1(n739), .A2(G234), .ZN(n460) );
  XOR2_X1 U579 ( .A(KEYINPUT8), .B(n460), .Z(n504) );
  NAND2_X1 U580 ( .A1(G217), .A2(n504), .ZN(n461) );
  XNOR2_X1 U581 ( .A(n463), .B(n462), .ZN(n711) );
  NOR2_X1 U582 ( .A1(G902), .A2(n711), .ZN(n464) );
  XOR2_X1 U583 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n468) );
  XOR2_X1 U584 ( .A(KEYINPUT69), .B(G131), .Z(n490) );
  XNOR2_X1 U585 ( .A(n490), .B(KEYINPUT11), .ZN(n467) );
  XNOR2_X1 U586 ( .A(n468), .B(n467), .ZN(n469) );
  XOR2_X1 U587 ( .A(n732), .B(n469), .Z(n475) );
  XOR2_X1 U588 ( .A(KEYINPUT75), .B(n470), .Z(n512) );
  NAND2_X1 U589 ( .A1(G214), .A2(n512), .ZN(n473) );
  NOR2_X1 U590 ( .A1(G902), .A2(n632), .ZN(n479) );
  XNOR2_X1 U591 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n477) );
  INV_X1 U592 ( .A(n565), .ZN(n546) );
  NOR2_X1 U593 ( .A1(n566), .A2(n546), .ZN(n480) );
  XNOR2_X1 U594 ( .A(n481), .B(KEYINPUT14), .ZN(n483) );
  NAND2_X1 U595 ( .A1(n483), .A2(G952), .ZN(n482) );
  XOR2_X1 U596 ( .A(KEYINPUT91), .B(n482), .Z(n697) );
  NOR2_X1 U597 ( .A1(G953), .A2(n697), .ZN(n581) );
  NAND2_X1 U598 ( .A1(G902), .A2(n483), .ZN(n578) );
  NOR2_X1 U599 ( .A1(G900), .A2(n578), .ZN(n485) );
  NAND2_X1 U600 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U601 ( .A(KEYINPUT109), .B(n486), .ZN(n487) );
  NOR2_X1 U602 ( .A1(n581), .A2(n487), .ZN(n541) );
  XOR2_X1 U603 ( .A(n490), .B(G134), .Z(n491) );
  XNOR2_X1 U604 ( .A(n528), .B(G140), .ZN(n494) );
  NAND2_X1 U605 ( .A1(G227), .A2(n739), .ZN(n493) );
  XNOR2_X1 U606 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U607 ( .A(n520), .B(n495), .ZN(n706) );
  XNOR2_X1 U608 ( .A(KEYINPUT21), .B(n499), .ZN(n667) );
  XOR2_X1 U609 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n500) );
  XNOR2_X1 U610 ( .A(G119), .B(G137), .ZN(n502) );
  NAND2_X1 U611 ( .A1(G221), .A2(n504), .ZN(n505) );
  XOR2_X1 U612 ( .A(KEYINPUT78), .B(KEYINPUT25), .Z(n509) );
  NAND2_X1 U613 ( .A1(n507), .A2(G217), .ZN(n508) );
  XNOR2_X1 U614 ( .A(n509), .B(n508), .ZN(n510) );
  AND2_X1 U615 ( .A1(n512), .A2(G210), .ZN(n514) );
  XNOR2_X1 U616 ( .A(G113), .B(KEYINPUT3), .ZN(n513) );
  XOR2_X1 U617 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n516) );
  XNOR2_X1 U618 ( .A(n516), .B(n515), .ZN(n517) );
  NAND2_X1 U619 ( .A1(G214), .A2(n537), .ZN(n521) );
  XNOR2_X1 U620 ( .A(KEYINPUT90), .B(n521), .ZN(n571) );
  INV_X1 U621 ( .A(n571), .ZN(n687) );
  XNOR2_X1 U622 ( .A(KEYINPUT30), .B(KEYINPUT111), .ZN(n522) );
  XOR2_X1 U623 ( .A(KEYINPUT17), .B(KEYINPUT89), .Z(n529) );
  NAND2_X1 U624 ( .A1(G224), .A2(n739), .ZN(n533) );
  XNOR2_X1 U625 ( .A(n534), .B(n533), .ZN(n535) );
  NAND2_X1 U626 ( .A1(n625), .A2(n619), .ZN(n539) );
  NAND2_X1 U627 ( .A1(G210), .A2(n537), .ZN(n538) );
  BUF_X1 U628 ( .A(n549), .Z(n575) );
  XNOR2_X1 U629 ( .A(KEYINPUT38), .B(n575), .ZN(n683) );
  NOR2_X1 U630 ( .A1(n655), .A2(n547), .ZN(n540) );
  XNOR2_X1 U631 ( .A(n540), .B(KEYINPUT112), .ZN(n746) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n685) );
  INV_X1 U633 ( .A(n685), .ZN(n600) );
  AND2_X1 U634 ( .A1(n683), .A2(n600), .ZN(n690) );
  NOR2_X1 U635 ( .A1(n541), .A2(n667), .ZN(n542) );
  NAND2_X1 U636 ( .A1(n542), .A2(n598), .ZN(n555) );
  NOR2_X1 U637 ( .A1(n611), .A2(n555), .ZN(n543) );
  XNOR2_X1 U638 ( .A(KEYINPUT28), .B(n543), .ZN(n544) );
  NAND2_X1 U639 ( .A1(n544), .A2(n562), .ZN(n552) );
  NOR2_X1 U640 ( .A1(n698), .A2(n552), .ZN(n545) );
  XNOR2_X1 U641 ( .A(KEYINPUT42), .B(n545), .ZN(n747) );
  NAND2_X1 U642 ( .A1(n566), .A2(n546), .ZN(n653) );
  NOR2_X2 U643 ( .A1(n549), .A2(n687), .ZN(n550) );
  XOR2_X1 U644 ( .A(KEYINPUT19), .B(KEYINPUT77), .Z(n551) );
  XNOR2_X1 U645 ( .A(n559), .B(n551), .ZN(n584) );
  OR2_X1 U646 ( .A1(n552), .A2(n584), .ZN(n553) );
  NAND2_X1 U647 ( .A1(n653), .A2(n655), .ZN(n684) );
  NAND2_X1 U648 ( .A1(n651), .A2(n684), .ZN(n554) );
  XNOR2_X1 U649 ( .A(KEYINPUT47), .B(n554), .ZN(n564) );
  INV_X1 U650 ( .A(n555), .ZN(n557) );
  NAND2_X1 U651 ( .A1(n557), .A2(n604), .ZN(n558) );
  NOR2_X1 U652 ( .A1(n653), .A2(n558), .ZN(n570) );
  NAND2_X1 U653 ( .A1(n559), .A2(n570), .ZN(n561) );
  XNOR2_X1 U654 ( .A(KEYINPUT36), .B(KEYINPUT85), .ZN(n560) );
  XNOR2_X1 U655 ( .A(n561), .B(n560), .ZN(n563) );
  INV_X2 U656 ( .A(n605), .ZN(n669) );
  NAND2_X1 U657 ( .A1(n563), .A2(n669), .ZN(n660) );
  NOR2_X1 U658 ( .A1(n566), .A2(n565), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n356), .A2(n588), .ZN(n567) );
  NOR2_X1 U660 ( .A1(n575), .A2(n567), .ZN(n650) );
  INV_X1 U661 ( .A(n650), .ZN(n568) );
  AND2_X1 U662 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U663 ( .A(KEYINPUT110), .B(n572), .ZN(n573) );
  NAND2_X1 U664 ( .A1(n573), .A2(n605), .ZN(n574) );
  XNOR2_X1 U665 ( .A(n574), .B(KEYINPUT43), .ZN(n576) );
  NAND2_X1 U666 ( .A1(n576), .A2(n575), .ZN(n661) );
  NAND2_X1 U667 ( .A1(n577), .A2(n661), .ZN(n737) );
  XOR2_X1 U668 ( .A(G898), .B(KEYINPUT92), .Z(n724) );
  NAND2_X1 U669 ( .A1(G953), .A2(n724), .ZN(n721) );
  NOR2_X1 U670 ( .A1(n578), .A2(n721), .ZN(n579) );
  XOR2_X1 U671 ( .A(KEYINPUT93), .B(n579), .Z(n580) );
  NOR2_X1 U672 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U673 ( .A(n582), .B(KEYINPUT94), .ZN(n583) );
  XOR2_X1 U674 ( .A(KEYINPUT108), .B(KEYINPUT33), .Z(n585) );
  XNOR2_X1 U675 ( .A(n586), .B(n585), .ZN(n699) );
  NOR2_X1 U676 ( .A1(n599), .A2(n699), .ZN(n587) );
  XNOR2_X1 U677 ( .A(n587), .B(KEYINPUT34), .ZN(n589) );
  NAND2_X1 U678 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X2 U679 ( .A(n590), .B(KEYINPUT35), .ZN(n743) );
  NAND2_X1 U680 ( .A1(n743), .A2(KEYINPUT44), .ZN(n597) );
  NOR2_X1 U681 ( .A1(n599), .A2(n678), .ZN(n592) );
  XNOR2_X1 U682 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n591) );
  XNOR2_X1 U683 ( .A(n592), .B(n591), .ZN(n656) );
  XNOR2_X1 U684 ( .A(KEYINPUT97), .B(n595), .ZN(n640) );
  NAND2_X1 U685 ( .A1(n597), .A2(n596), .ZN(n608) );
  XOR2_X1 U686 ( .A(KEYINPUT106), .B(n345), .Z(n666) );
  XOR2_X1 U687 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n601) );
  XNOR2_X1 U688 ( .A(n606), .B(KEYINPUT83), .ZN(n607) );
  NOR2_X1 U689 ( .A1(n669), .A2(n609), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n613), .A2(n743), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n616), .A2(KEYINPUT71), .ZN(n617) );
  INV_X1 U692 ( .A(n619), .ZN(n620) );
  XOR2_X1 U693 ( .A(n620), .B(KEYINPUT81), .Z(n621) );
  NAND2_X1 U694 ( .A1(n621), .A2(KEYINPUT2), .ZN(n622) );
  XNOR2_X1 U695 ( .A(KEYINPUT66), .B(n622), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n662), .A2(KEYINPUT2), .ZN(n665) );
  XOR2_X1 U697 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n627) );
  XNOR2_X1 U698 ( .A(n625), .B(KEYINPUT55), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n627), .B(n626), .ZN(n628) );
  INV_X1 U700 ( .A(n717), .ZN(n629) );
  INV_X1 U701 ( .A(KEYINPUT123), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n630), .B(KEYINPUT56), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n455), .B(n631), .ZN(G51) );
  INV_X1 U704 ( .A(KEYINPUT125), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n634), .B(KEYINPUT62), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n636), .B(G101), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT113), .ZN(G3) );
  NOR2_X1 U708 ( .A1(n653), .A2(n640), .ZN(n638) );
  XOR2_X1 U709 ( .A(KEYINPUT114), .B(n638), .Z(n639) );
  XNOR2_X1 U710 ( .A(G104), .B(n639), .ZN(G6) );
  NOR2_X1 U711 ( .A1(n655), .A2(n640), .ZN(n645) );
  XOR2_X1 U712 ( .A(KEYINPUT27), .B(KEYINPUT116), .Z(n642) );
  XNOR2_X1 U713 ( .A(G107), .B(KEYINPUT115), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U715 ( .A(KEYINPUT26), .B(n643), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(G9) );
  XOR2_X1 U717 ( .A(G110), .B(n646), .Z(G12) );
  XOR2_X1 U718 ( .A(G128), .B(KEYINPUT29), .Z(n649) );
  NAND2_X1 U719 ( .A1(n651), .A2(n647), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(G30) );
  XOR2_X1 U721 ( .A(G143), .B(n650), .Z(G45) );
  NAND2_X1 U722 ( .A1(n427), .A2(n651), .ZN(n652) );
  XNOR2_X1 U723 ( .A(G146), .B(n652), .ZN(G48) );
  NOR2_X1 U724 ( .A1(n656), .A2(n653), .ZN(n654) );
  XOR2_X1 U725 ( .A(G113), .B(n654), .Z(G15) );
  NOR2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n658) );
  XNOR2_X1 U727 ( .A(G116), .B(KEYINPUT117), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n658), .B(n657), .ZN(G18) );
  XOR2_X1 U729 ( .A(G125), .B(KEYINPUT37), .Z(n659) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(G27) );
  XNOR2_X1 U731 ( .A(G140), .B(n661), .ZN(G42) );
  NOR2_X1 U732 ( .A1(n662), .A2(KEYINPUT2), .ZN(n663) );
  XOR2_X1 U733 ( .A(KEYINPUT80), .B(n663), .Z(n664) );
  NAND2_X1 U734 ( .A1(n665), .A2(n664), .ZN(n703) );
  NAND2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U736 ( .A(KEYINPUT49), .B(n668), .ZN(n675) );
  NOR2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n672) );
  XNOR2_X1 U738 ( .A(KEYINPUT119), .B(KEYINPUT50), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n672), .B(n671), .ZN(n673) );
  XOR2_X1 U740 ( .A(KEYINPUT118), .B(n673), .Z(n674) );
  NOR2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n677) );
  INV_X1 U742 ( .A(n556), .ZN(n676) );
  NAND2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U745 ( .A(n680), .B(KEYINPUT120), .ZN(n681) );
  XNOR2_X1 U746 ( .A(n681), .B(KEYINPUT51), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n698), .A2(n682), .ZN(n693) );
  NAND2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n686) );
  AND2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U752 ( .A1(n699), .A2(n691), .ZN(n692) );
  NOR2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U754 ( .A(n694), .B(KEYINPUT52), .Z(n695) );
  XNOR2_X1 U755 ( .A(KEYINPUT121), .B(n695), .ZN(n696) );
  NOR2_X1 U756 ( .A1(n697), .A2(n696), .ZN(n701) );
  NOR2_X1 U757 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U758 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U759 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n704), .A2(G953), .ZN(n705) );
  XNOR2_X1 U761 ( .A(n705), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U762 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n706), .B(KEYINPUT57), .ZN(n707) );
  XNOR2_X1 U764 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U765 ( .A1(G478), .A2(n713), .ZN(n710) );
  XNOR2_X1 U766 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U767 ( .A1(n717), .A2(n712), .ZN(G63) );
  NAND2_X1 U768 ( .A1(G217), .A2(n713), .ZN(n714) );
  XNOR2_X1 U769 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U770 ( .A1(n717), .A2(n716), .ZN(G66) );
  XOR2_X1 U771 ( .A(n719), .B(n718), .Z(n720) );
  NAND2_X1 U772 ( .A1(n721), .A2(n720), .ZN(n730) );
  NAND2_X1 U773 ( .A1(G953), .A2(G224), .ZN(n722) );
  XOR2_X1 U774 ( .A(KEYINPUT61), .B(n722), .Z(n723) );
  NOR2_X1 U775 ( .A1(n724), .A2(n723), .ZN(n728) );
  NOR2_X1 U776 ( .A1(G953), .A2(n725), .ZN(n726) );
  XNOR2_X1 U777 ( .A(n726), .B(KEYINPUT126), .ZN(n727) );
  NOR2_X1 U778 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(G69) );
  XNOR2_X1 U780 ( .A(n732), .B(n731), .ZN(n736) );
  INV_X1 U781 ( .A(n736), .ZN(n733) );
  XOR2_X1 U782 ( .A(G227), .B(n733), .Z(n734) );
  NAND2_X1 U783 ( .A1(n734), .A2(G900), .ZN(n735) );
  NAND2_X1 U784 ( .A1(n735), .A2(G953), .ZN(n742) );
  XOR2_X1 U785 ( .A(n737), .B(n736), .Z(n738) );
  XNOR2_X1 U786 ( .A(n738), .B(KEYINPUT127), .ZN(n740) );
  NAND2_X1 U787 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U788 ( .A1(n742), .A2(n741), .ZN(G72) );
  XOR2_X1 U789 ( .A(n743), .B(G122), .Z(G24) );
  XOR2_X1 U790 ( .A(n744), .B(G119), .Z(G21) );
  XOR2_X1 U791 ( .A(n745), .B(G131), .Z(G33) );
  XOR2_X1 U792 ( .A(n746), .B(G134), .Z(G36) );
  XOR2_X1 U793 ( .A(n747), .B(G137), .Z(G39) );
endmodule

