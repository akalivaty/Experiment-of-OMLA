//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  NAND2_X1  g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G68), .A2(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n217), .B(new_n218), .C1(new_n202), .C2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n216), .B(new_n220), .C1(G97), .C2(G257), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G1), .B2(G20), .ZN(new_n222));
  XOR2_X1   g0022(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n223));
  XNOR2_X1  g0023(.A(new_n222), .B(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n210), .B(new_n224), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G226), .B(G232), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G232), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G1698), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G226), .B2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G97), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n249), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT70), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n248), .A2(G238), .A3(new_n263), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n261), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT13), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT71), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT13), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n261), .B(new_n273), .C1(new_n268), .C2(new_n269), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n270), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(G169), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT72), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT73), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n275), .A2(new_n280), .A3(G169), .A4(new_n276), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n279), .B(KEYINPUT14), .C1(new_n278), .C2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n271), .A2(new_n274), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G179), .ZN(new_n284));
  INV_X1    g0084(.A(new_n281), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n282), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT67), .B1(new_n207), .B2(new_n255), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n225), .A3(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n226), .A2(G33), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n294), .A2(new_n202), .B1(new_n295), .B2(new_n212), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n226), .A2(G68), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT11), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n292), .B1(new_n262), .B2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G68), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(new_n299), .ZN(new_n303));
  INV_X1    g0103(.A(G13), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G1), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT12), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n300), .A2(new_n302), .A3(new_n303), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n288), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n283), .A2(G190), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n275), .A2(G200), .A3(new_n276), .ZN(new_n311));
  INV_X1    g0111(.A(new_n308), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G20), .A2(G77), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT8), .B(G58), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT15), .B(G87), .Z(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n314), .B1(new_n294), .B2(new_n315), .C1(new_n317), .C2(new_n295), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(new_n292), .B1(G77), .B2(new_n301), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n305), .A2(G20), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(G77), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT3), .B(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G238), .A2(G1698), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n322), .B(new_n323), .C1(new_n250), .C2(G1698), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n324), .B(new_n249), .C1(G107), .C2(new_n322), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n248), .A2(new_n263), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n325), .B(new_n265), .C1(new_n213), .C2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n321), .B1(G200), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(new_n327), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n309), .A2(new_n313), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G58), .ZN(new_n332));
  INV_X1    g0132(.A(G68), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(G20), .B1(new_n334), .B2(new_n201), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n293), .A2(G159), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n322), .B2(G20), .ZN(new_n339));
  INV_X1    g0139(.A(new_n256), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n255), .A2(KEYINPUT74), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT74), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n340), .B1(new_n344), .B2(new_n253), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n338), .A2(G20), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n339), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n337), .B1(new_n348), .B2(G68), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT75), .B1(new_n349), .B2(KEYINPUT16), .ZN(new_n350));
  INV_X1    g0150(.A(new_n254), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT74), .B(G33), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(KEYINPUT3), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT7), .B1(new_n353), .B2(G20), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n254), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(new_n338), .A3(new_n226), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(G68), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n337), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT75), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT16), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT3), .B1(new_n341), .B2(new_n343), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n346), .B1(new_n363), .B2(new_n340), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n333), .B1(new_n364), .B2(new_n339), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n361), .B(new_n362), .C1(new_n365), .C2(new_n337), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n350), .A2(new_n292), .A3(new_n360), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n320), .A2(new_n315), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n301), .B2(new_n315), .ZN(new_n369));
  INV_X1    g0169(.A(new_n265), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n219), .A2(G1698), .ZN(new_n371));
  OR2_X1    g0171(.A1(G223), .A2(G1698), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n355), .A2(new_n254), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G87), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n370), .B1(new_n375), .B2(new_n249), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n326), .A2(new_n250), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n329), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n248), .B1(new_n373), .B2(new_n374), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n380), .A2(new_n370), .A3(new_n377), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n379), .B1(new_n381), .B2(G200), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n367), .A2(new_n369), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT76), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT17), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n385), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n386), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n367), .A2(new_n369), .ZN(new_n390));
  INV_X1    g0190(.A(G169), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n376), .B2(new_n378), .ZN(new_n392));
  INV_X1    g0192(.A(G179), .ZN(new_n393));
  NOR4_X1   g0193(.A1(new_n380), .A2(new_n393), .A3(new_n370), .A4(new_n377), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT18), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n398), .B(new_n395), .C1(new_n367), .C2(new_n369), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n387), .A2(new_n389), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G223), .A2(G1698), .ZN(new_n402));
  INV_X1    g0202(.A(G1698), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G222), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n322), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(new_n249), .C1(G77), .C2(new_n322), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n406), .B(new_n265), .C1(new_n219), .C2(new_n326), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n407), .A2(G179), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n203), .A2(G20), .ZN(new_n409));
  INV_X1    g0209(.A(G150), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n409), .B1(new_n410), .B2(new_n294), .C1(new_n315), .C2(new_n295), .ZN(new_n411));
  INV_X1    g0211(.A(new_n320), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n411), .A2(new_n292), .B1(new_n202), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n292), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n202), .B1(new_n262), .B2(G20), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(KEYINPUT68), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(KEYINPUT68), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n414), .A2(new_n416), .A3(new_n320), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n407), .A2(new_n391), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n408), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n327), .A2(G179), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n327), .A2(new_n391), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n321), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n413), .A2(new_n418), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(KEYINPUT9), .B1(G200), .B2(new_n407), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n407), .A2(new_n329), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT69), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT9), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n419), .B2(new_n430), .ZN(new_n431));
  AOI211_X1 g0231(.A(KEYINPUT69), .B(KEYINPUT9), .C1(new_n413), .C2(new_n418), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n427), .B(new_n428), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT10), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT9), .B1(new_n413), .B2(new_n418), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n435), .B(new_n429), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT10), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n428), .A4(new_n427), .ZN(new_n438));
  AOI211_X1 g0238(.A(new_n421), .B(new_n425), .C1(new_n434), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n401), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n331), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n305), .ZN(new_n442));
  INV_X1    g0242(.A(G107), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G20), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT25), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n442), .A2(KEYINPUT25), .A3(new_n444), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n255), .A2(G1), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n292), .A2(new_n412), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n446), .B1(new_n448), .B2(G107), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n214), .A2(G20), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n254), .A3(new_n256), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT22), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n344), .A2(new_n226), .A3(G116), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT23), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n444), .B(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n355), .A2(KEYINPUT22), .A3(new_n254), .A4(new_n450), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT84), .B(KEYINPUT24), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT85), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n455), .A2(new_n457), .A3(new_n458), .A4(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n458), .A2(new_n453), .A3(new_n457), .A4(new_n454), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n461), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n463), .A2(new_n465), .B1(new_n460), .B2(new_n459), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n445), .B(new_n449), .C1(new_n466), .C2(new_n414), .ZN(new_n467));
  INV_X1    g0267(.A(G257), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n215), .A2(new_n403), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n355), .A2(new_n254), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n344), .A2(G294), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n248), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G45), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G1), .ZN(new_n475));
  AND2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  NOR2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n248), .ZN(new_n479));
  INV_X1    g0279(.A(G264), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n475), .B(G274), .C1(new_n477), .C2(new_n476), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NOR4_X1   g0283(.A1(new_n473), .A2(new_n481), .A3(G190), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G200), .ZN(new_n485));
  INV_X1    g0285(.A(new_n481), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n471), .A2(new_n472), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n482), .C1(new_n487), .C2(new_n248), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n484), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n467), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n473), .A2(new_n483), .A3(new_n481), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(KEYINPUT86), .A3(G179), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT86), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n488), .B2(G169), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n488), .A2(new_n393), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n467), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G238), .A2(G1698), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n213), .B2(G1698), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(new_n355), .A3(new_n254), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n344), .A2(G116), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n248), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n475), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G250), .A3(new_n248), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n505), .A2(new_n264), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(G169), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NOR4_X1   g0311(.A1(new_n504), .A2(G179), .A3(new_n509), .A4(new_n507), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n355), .A2(new_n226), .A3(G68), .A4(new_n254), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n259), .A2(KEYINPUT77), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT77), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G97), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n515), .B1(new_n519), .B2(new_n295), .ZN(new_n520));
  AOI21_X1  g0320(.A(G87), .B1(new_n516), .B2(new_n518), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n521), .A2(new_n443), .ZN(new_n522));
  AOI21_X1  g0322(.A(G20), .B1(new_n260), .B2(KEYINPUT19), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n514), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(new_n292), .B1(new_n412), .B2(new_n317), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n448), .A2(new_n316), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT81), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n514), .A2(new_n520), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n523), .B1(new_n443), .B2(new_n521), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n292), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n317), .A2(new_n412), .ZN(new_n531));
  AND4_X1   g0331(.A1(KEYINPUT81), .A2(new_n530), .A3(new_n526), .A4(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n513), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n448), .A2(G87), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n525), .A2(new_n534), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n504), .A2(new_n509), .A3(new_n507), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G190), .ZN(new_n537));
  INV_X1    g0337(.A(new_n536), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G200), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n293), .A2(G77), .ZN(new_n542));
  XOR2_X1   g0342(.A(G97), .B(G107), .Z(new_n543));
  NAND2_X1  g0343(.A1(new_n443), .A2(KEYINPUT6), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n543), .A2(KEYINPUT6), .B1(new_n519), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G20), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n256), .B1(new_n352), .B2(KEYINPUT3), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n257), .A2(new_n226), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n547), .A2(new_n346), .B1(new_n548), .B2(new_n338), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n542), .B(new_n546), .C1(new_n549), .C2(new_n443), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n292), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n320), .A2(G97), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n447), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n414), .A2(new_n320), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n555), .B2(new_n259), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n355), .A2(G244), .A3(new_n254), .ZN(new_n559));
  XNOR2_X1  g0359(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(new_n257), .B2(new_n215), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G1698), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n403), .A2(KEYINPUT4), .A3(G244), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n322), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G283), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT79), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n562), .A2(new_n564), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n249), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n482), .B1(new_n479), .B2(new_n468), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n391), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  AOI211_X1 g0377(.A(new_n393), .B(new_n575), .C1(new_n573), .C2(new_n249), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n558), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n556), .B1(new_n550), .B2(new_n292), .ZN(new_n580));
  AOI21_X1  g0380(.A(G200), .B1(new_n574), .B2(new_n576), .ZN(new_n581));
  AOI211_X1 g0381(.A(G190), .B(new_n575), .C1(new_n573), .C2(new_n249), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n579), .A2(new_n583), .A3(KEYINPUT80), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n541), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT82), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n499), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n480), .A2(G1698), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n468), .A2(new_n403), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n355), .A2(new_n254), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(new_n322), .ZN(new_n595));
  INV_X1    g0395(.A(new_n479), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n595), .A2(new_n249), .B1(G270), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n597), .A2(new_n482), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT20), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n516), .A2(new_n518), .A3(new_n255), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n600), .A2(new_n571), .A3(new_n226), .ZN(new_n601));
  INV_X1    g0401(.A(G116), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n292), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n599), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n600), .A2(new_n571), .A3(new_n226), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT20), .A3(new_n292), .A4(new_n603), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n305), .A2(G20), .A3(new_n602), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n414), .A2(G116), .A3(new_n320), .A4(new_n554), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT83), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n448), .A2(KEYINPUT83), .A3(G116), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n608), .A2(new_n609), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n598), .A2(new_n614), .A3(G179), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n391), .B1(new_n597), .B2(new_n482), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n614), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT21), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n615), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n598), .A2(G190), .ZN(new_n622));
  INV_X1    g0422(.A(new_n614), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n622), .B(new_n623), .C1(new_n485), .C2(new_n598), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n533), .A2(new_n540), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n579), .A2(new_n583), .A3(KEYINPUT80), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT80), .B1(new_n579), .B2(new_n583), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n625), .B1(new_n629), .B2(KEYINPUT82), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n441), .A2(new_n590), .A3(new_n630), .ZN(G372));
  NAND2_X1  g0431(.A1(new_n434), .A2(new_n438), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n313), .A2(new_n425), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n383), .A2(new_n386), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n383), .A2(new_n388), .ZN(new_n635));
  INV_X1    g0435(.A(new_n386), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n309), .A2(new_n633), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n397), .A2(new_n399), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n632), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n421), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n618), .A2(new_n620), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n598), .A2(new_n614), .A3(G179), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n498), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n584), .A2(new_n490), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n626), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n566), .A2(new_n571), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(G1698), .B2(new_n563), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n248), .B1(new_n650), .B2(new_n562), .ZN(new_n651));
  OAI21_X1  g0451(.A(G169), .B1(new_n651), .B2(new_n575), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n574), .A2(G179), .A3(new_n576), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n580), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n533), .A2(new_n540), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n533), .A2(new_n540), .A3(new_n654), .A4(KEYINPUT26), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n648), .A2(new_n659), .A3(new_n533), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n441), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n643), .A2(new_n661), .ZN(G369));
  INV_X1    g0462(.A(new_n467), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT87), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n304), .A2(G20), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(new_n262), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n262), .A2(new_n226), .A3(G13), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n667), .A2(new_n669), .A3(G213), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n664), .B1(new_n670), .B2(G343), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(new_n664), .A3(G343), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n663), .A2(new_n675), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n499), .A2(new_n676), .B1(new_n498), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n614), .A2(new_n674), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT88), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT89), .B1(new_n621), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n620), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n619), .B1(new_n616), .B2(new_n614), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n645), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT88), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n678), .B(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT89), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n621), .A2(new_n679), .A3(new_n624), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n680), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n689), .A2(KEYINPUT90), .A3(G330), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT90), .B1(new_n689), .B2(G330), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n677), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n498), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT91), .ZN(new_n694));
  INV_X1    g0494(.A(new_n673), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n671), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n672), .A2(KEYINPUT91), .A3(new_n673), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n683), .A2(new_n491), .A3(new_n498), .A4(new_n675), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n692), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0503(.A(new_n208), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G1), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n522), .A2(new_n602), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n707), .A2(new_n708), .B1(new_n228), .B2(new_n706), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT93), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n590), .A2(new_n630), .A3(new_n699), .ZN(new_n712));
  XNOR2_X1  g0512(.A(KEYINPUT94), .B(KEYINPUT31), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n574), .A2(new_n536), .A3(new_n576), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n492), .A2(new_n597), .A3(G179), .ZN(new_n716));
  OR3_X1    g0516(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT30), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT30), .B1(new_n715), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n598), .B1(new_n574), .B2(new_n576), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n393), .A3(new_n538), .A4(new_n488), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n714), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n722), .A2(KEYINPUT95), .A3(new_n698), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT95), .B1(new_n722), .B2(new_n698), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n675), .B1(new_n719), .B2(new_n721), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT31), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n712), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n660), .A2(new_n675), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT96), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT96), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n660), .A2(new_n732), .A3(new_n675), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(KEYINPUT29), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n660), .A2(new_n699), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n729), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n711), .B1(new_n738), .B2(G1), .ZN(G364));
  NOR2_X1   g0539(.A1(new_n226), .A2(G190), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G179), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT101), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(KEYINPUT101), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n226), .A2(new_n329), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n393), .A2(new_n485), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT99), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n749), .B1(new_n747), .B2(new_n748), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n746), .A2(G329), .B1(new_n753), .B2(G326), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n485), .A2(G179), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n740), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n322), .B1(new_n757), .B2(G283), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n747), .A2(new_n755), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n393), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n747), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G303), .A2(new_n760), .B1(new_n763), .B2(G322), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n748), .A2(new_n740), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G317), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(KEYINPUT33), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n767), .A2(KEYINPUT33), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AND4_X1   g0570(.A1(new_n754), .A2(new_n758), .A3(new_n764), .A4(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G294), .ZN(new_n772));
  INV_X1    g0572(.A(new_n741), .ZN(new_n773));
  OAI21_X1  g0573(.A(G20), .B1(new_n773), .B2(new_n329), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT102), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n774), .A2(new_n775), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n740), .A2(new_n761), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n771), .B1(new_n772), .B2(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n781), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n753), .A2(G50), .B1(G77), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n332), .B2(new_n762), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT100), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n746), .A2(G159), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT32), .ZN(new_n788));
  INV_X1    g0588(.A(new_n779), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G97), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n322), .B1(new_n756), .B2(new_n443), .C1(new_n333), .C2(new_n765), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n787), .B2(KEYINPUT32), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n786), .A2(new_n788), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n759), .A2(new_n214), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n782), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n225), .B1(G20), .B2(new_n391), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G13), .A2(G33), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT98), .Z(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G20), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n796), .ZN(new_n800));
  NAND3_X1  g0600(.A1(G355), .A2(new_n208), .A3(new_n322), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n242), .A2(G45), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n353), .A2(new_n704), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G45), .B2(new_n228), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n801), .B1(G116), .B2(new_n208), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n795), .A2(new_n796), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n665), .A2(G45), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n706), .A2(G1), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT97), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n799), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n806), .B(new_n810), .C1(new_n689), .C2(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n690), .A2(new_n691), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n808), .B1(new_n689), .B2(G330), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(G396));
  NOR2_X1   g0615(.A1(new_n424), .A2(new_n674), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n321), .A2(new_n674), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n330), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n816), .B1(new_n818), .B2(new_n424), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n735), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n660), .A2(new_n699), .A3(new_n819), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n729), .B(new_n823), .Z(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n808), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n757), .A2(G87), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n826), .B1(new_n602), .B2(new_n781), .C1(new_n827), .C2(new_n765), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n322), .B(new_n828), .C1(G294), .C2(new_n763), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n760), .A2(G107), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n746), .A2(G311), .B1(new_n753), .B2(G303), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n829), .A2(new_n790), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G143), .ZN(new_n833));
  INV_X1    g0633(.A(G159), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n762), .A2(new_n833), .B1(new_n781), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n753), .B2(G137), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n410), .B2(new_n765), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n757), .A2(G68), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n789), .A2(G58), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n746), .A2(G132), .B1(G50), .B2(new_n760), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n832), .B1(new_n842), .B2(new_n356), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n796), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n798), .B2(new_n819), .ZN(new_n845));
  INV_X1    g0645(.A(new_n798), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n796), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT103), .Z(new_n848));
  OAI21_X1  g0648(.A(new_n810), .B1(new_n848), .B2(G77), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT104), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n825), .B1(new_n845), .B2(new_n850), .ZN(G384));
  INV_X1    g0651(.A(KEYINPUT40), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n714), .A2(KEYINPUT108), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n726), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT31), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n713), .B2(KEYINPUT108), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n854), .B1(new_n726), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n712), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n308), .A2(new_n674), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n309), .A2(new_n313), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n313), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n308), .B(new_n674), .C1(new_n288), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n858), .A2(new_n819), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n360), .A2(new_n292), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT16), .B1(new_n358), .B2(new_n359), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n369), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n400), .A2(new_n670), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n396), .B2(new_n670), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n383), .ZN(new_n870));
  INV_X1    g0670(.A(new_n383), .ZN(new_n871));
  INV_X1    g0671(.A(new_n670), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n367), .A2(new_n369), .B1(new_n395), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  MUX2_X1   g0675(.A(new_n870), .B(new_n874), .S(new_n875), .Z(new_n876));
  AND3_X1   g0676(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n868), .B2(new_n876), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n852), .B1(new_n864), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n876), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT106), .B1(new_n390), .B2(new_n670), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n882), .A2(new_n875), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n874), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n882), .A2(new_n875), .B1(new_n871), .B2(new_n873), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT107), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n637), .A2(new_n887), .A3(new_n634), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT107), .B1(new_n387), .B2(new_n389), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n639), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n390), .A2(new_n670), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n886), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n881), .B1(new_n893), .B2(KEYINPUT38), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n820), .B1(new_n712), .B2(new_n857), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n894), .A2(KEYINPUT40), .A3(new_n863), .A4(new_n895), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n880), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n858), .A2(new_n441), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n897), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(G330), .ZN(new_n900));
  INV_X1    g0700(.A(new_n816), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT105), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n901), .A2(KEYINPUT105), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n822), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n863), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n905), .A2(new_n879), .B1(new_n639), .B2(new_n670), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n877), .A2(new_n878), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n907), .B2(new_n894), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n309), .A2(new_n674), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n734), .A2(new_n736), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n441), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n643), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n911), .B(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n900), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n262), .B2(new_n665), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n602), .B1(new_n545), .B2(KEYINPUT35), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(new_n227), .C1(KEYINPUT35), .C2(new_n545), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT36), .ZN(new_n920));
  OAI21_X1  g0720(.A(G77), .B1(new_n332), .B2(new_n333), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n921), .A2(new_n228), .B1(G50), .B2(new_n333), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(G1), .A3(new_n304), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n917), .A2(new_n920), .A3(new_n923), .ZN(G367));
  NAND2_X1  g0724(.A1(new_n807), .A2(G1), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n692), .A2(KEYINPUT114), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT114), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n928), .B(new_n677), .C1(new_n690), .C2(new_n691), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n701), .A2(new_n700), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT110), .B1(new_n579), .B2(new_n699), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT110), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n654), .A2(new_n932), .A3(new_n698), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n579), .B(new_n583), .C1(new_n580), .C2(new_n699), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT44), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n930), .A2(new_n937), .A3(KEYINPUT44), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT45), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n930), .B2(new_n937), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n936), .A2(new_n701), .A3(KEYINPUT45), .A4(new_n700), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n940), .A2(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n927), .A2(new_n929), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n940), .A2(new_n941), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n943), .A2(new_n944), .ZN(new_n948));
  OAI211_X1 g0748(.A(KEYINPUT114), .B(new_n692), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n683), .A2(new_n675), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n701), .B1(new_n677), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n813), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n737), .B1(new_n950), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n705), .B(KEYINPUT41), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n926), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n535), .A2(new_n675), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n626), .A2(KEYINPUT109), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT109), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n541), .B2(new_n959), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n961), .B(new_n963), .C1(new_n533), .C2(new_n960), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT112), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT111), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n936), .A2(new_n693), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n698), .B1(new_n968), .B2(new_n579), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT42), .ZN(new_n970));
  INV_X1    g0770(.A(new_n701), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n970), .B1(new_n971), .B2(new_n936), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n967), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT42), .B1(new_n937), .B2(new_n701), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n498), .B1(new_n934), .B2(new_n935), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n699), .B1(new_n975), .B2(new_n654), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(new_n976), .A3(KEYINPUT111), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n937), .A2(KEYINPUT42), .A3(new_n701), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n966), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  AOI211_X1 g0781(.A(KEYINPUT112), .B(new_n979), .C1(new_n973), .C2(new_n977), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n965), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n977), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT111), .B1(new_n974), .B2(new_n976), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n980), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT112), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n964), .B(KEYINPUT43), .Z(new_n988));
  NAND3_X1  g0788(.A1(new_n978), .A2(new_n966), .A3(new_n980), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n813), .A2(new_n677), .A3(new_n936), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(KEYINPUT113), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n983), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n991), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT113), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n983), .A2(new_n990), .A3(new_n995), .A4(new_n994), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n958), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT115), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n958), .A2(new_n997), .A3(KEYINPUT115), .A4(new_n998), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n779), .A2(new_n333), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n322), .B1(new_n781), .B2(new_n202), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n762), .A2(new_n410), .B1(new_n756), .B2(new_n212), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G58), .C2(new_n760), .ZN(new_n1007));
  INV_X1    g0807(.A(G137), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n745), .C1(new_n833), .C2(new_n752), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1004), .B(new_n1009), .C1(G159), .C2(new_n766), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G303), .A2(new_n763), .B1(new_n783), .B2(G283), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n519), .B2(new_n756), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n753), .B2(G311), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n772), .B2(new_n765), .C1(new_n767), .C2(new_n745), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n356), .B1(new_n779), .B2(new_n443), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n759), .A2(new_n602), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT46), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1010), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT47), .Z(new_n1020));
  AOI21_X1  g0820(.A(new_n809), .B1(new_n1020), .B2(new_n796), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n803), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n800), .B1(new_n208), .B2(new_n317), .C1(new_n238), .C2(new_n1022), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n964), .A2(new_n811), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1003), .A2(new_n1025), .ZN(G387));
  INV_X1    g0826(.A(new_n954), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n737), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n954), .A2(new_n738), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n705), .A3(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n746), .A2(G326), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G311), .A2(new_n766), .B1(new_n783), .B2(G303), .ZN(new_n1032));
  INV_X1    g0832(.A(G322), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1032), .B1(new_n767), .B2(new_n762), .C1(new_n752), .C2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT48), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n827), .B2(new_n779), .C1(new_n772), .C2(new_n759), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT49), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n353), .B(new_n1031), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n1037), .B2(new_n1036), .C1(new_n602), .C2(new_n756), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n765), .A2(new_n315), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n760), .A2(G77), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n756), .B2(new_n259), .C1(new_n202), .C2(new_n762), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n356), .B(new_n1042), .C1(G68), .C2(new_n783), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n789), .A2(new_n316), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n746), .A2(G150), .B1(new_n753), .B2(G159), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1039), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n809), .B1(new_n1047), .B2(new_n796), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n315), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n202), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT50), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n333), .A2(new_n212), .ZN(new_n1052));
  NOR4_X1   g0852(.A1(new_n1051), .A2(G45), .A3(new_n1052), .A4(new_n708), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n803), .B1(new_n235), .B2(new_n474), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n708), .A2(new_n208), .A3(new_n322), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n208), .A2(G107), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n800), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1048), .B(new_n1058), .C1(new_n677), .C2(new_n811), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1030), .B(new_n1059), .C1(new_n926), .C2(new_n1027), .ZN(G393));
  AND2_X1   g0860(.A1(new_n946), .A2(new_n949), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n706), .B1(new_n1061), .B2(new_n1029), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n1029), .B2(new_n1061), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n937), .A2(new_n799), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n800), .B1(new_n208), .B2(new_n519), .C1(new_n245), .C2(new_n1022), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n826), .B1(new_n202), .B2(new_n765), .C1(new_n315), .C2(new_n781), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n356), .B(new_n1066), .C1(G143), .C2(new_n746), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n760), .A2(G68), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n752), .A2(new_n410), .B1(new_n834), .B2(new_n762), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n779), .A2(new_n212), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n789), .A2(G116), .B1(G303), .B2(new_n766), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n752), .A2(new_n767), .B1(new_n780), .B2(new_n762), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n257), .B1(new_n756), .B2(new_n443), .C1(new_n827), .C2(new_n759), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n746), .B2(G322), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n781), .A2(new_n772), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1073), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n809), .B1(new_n1083), .B2(new_n796), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1064), .A2(new_n1065), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n950), .B2(new_n925), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1063), .A2(new_n1086), .ZN(G390));
  OAI221_X1 g0887(.A(new_n839), .B1(new_n443), .B2(new_n765), .C1(new_n602), .C2(new_n762), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1088), .A2(new_n322), .A3(new_n794), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n827), .B2(new_n752), .C1(new_n772), .C2(new_n745), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n781), .A2(new_n519), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1090), .A2(new_n1071), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n257), .B1(new_n757), .B2(G50), .ZN(new_n1093));
  XOR2_X1   g0893(.A(KEYINPUT54), .B(G143), .Z(new_n1094));
  AOI22_X1  g0894(.A1(G132), .A2(new_n763), .B1(new_n783), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(new_n779), .C2(new_n834), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n746), .A2(G125), .B1(new_n753), .B2(G128), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n759), .A2(new_n410), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT53), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1096), .B(new_n1100), .C1(G137), .C2(new_n766), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n796), .B1(new_n1092), .B2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1102), .A2(new_n810), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n1049), .B2(new_n848), .C1(new_n909), .C2(new_n798), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n895), .A2(G330), .A3(new_n863), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n863), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n818), .A2(new_n424), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n660), .A2(new_n732), .A3(new_n675), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n732), .B1(new_n660), .B2(new_n675), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1106), .B1(new_n1110), .B2(new_n901), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT117), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n910), .B(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n894), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n894), .A2(new_n907), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n878), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n910), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1116), .A2(new_n1118), .B1(new_n1119), .B2(new_n905), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1105), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n905), .A2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1107), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n731), .B2(new_n733), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n863), .B1(new_n1126), .B2(new_n816), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1113), .A2(new_n894), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n728), .A2(G330), .A3(new_n819), .A4(new_n863), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1124), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1121), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1104), .B1(new_n1133), .B2(new_n926), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n858), .A2(new_n441), .A3(G330), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT118), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n858), .A2(new_n441), .A3(KEYINPUT118), .A4(G330), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(new_n913), .A3(new_n643), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1126), .A2(new_n816), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n858), .A2(G330), .A3(new_n819), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1142), .A2(KEYINPUT119), .A3(new_n1106), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT119), .B1(new_n1142), .B2(new_n1106), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1141), .B(new_n1130), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n728), .A2(G330), .A3(new_n819), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1106), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1105), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n904), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1140), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n706), .B1(new_n1151), .B2(new_n1133), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1121), .A2(new_n1132), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1150), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1134), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(G378));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n632), .A2(new_n642), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT121), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n419), .A2(new_n670), .ZN(new_n1160));
  XOR2_X1   g0960(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1161));
  XNOR2_X1  g0961(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1159), .B(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n880), .A2(new_n896), .A3(G330), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT122), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n880), .A2(new_n896), .A3(KEYINPUT122), .A4(G330), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1116), .A2(new_n910), .A3(new_n1118), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n906), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n911), .A2(new_n1168), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1167), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1170), .A2(new_n1169), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1174), .A2(new_n897), .A3(KEYINPUT122), .A4(G330), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n911), .A2(new_n1168), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n1166), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1140), .B1(new_n1153), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1157), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1140), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1154), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1177), .A4(new_n1173), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1181), .A2(new_n705), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1163), .A2(new_n846), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n848), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n202), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G128), .A2(new_n763), .B1(new_n766), .B2(G132), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n1008), .B2(new_n781), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n753), .B2(G125), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1094), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1191), .B1(new_n410), .B2(new_n779), .C1(new_n759), .C2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT59), .Z(new_n1194));
  AOI21_X1  g0994(.A(G41), .B1(new_n746), .B2(G124), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G33), .B1(new_n757), .B2(G159), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n763), .A2(G107), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n766), .A2(G97), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n783), .A2(new_n316), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1041), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NOR4_X1   g1001(.A1(new_n1004), .A2(new_n1201), .A3(G41), .A4(new_n353), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n756), .A2(new_n332), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT120), .Z(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G283), .B2(new_n746), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1202), .B(new_n1206), .C1(new_n602), .C2(new_n752), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT58), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n343), .ZN(new_n1209));
  AOI21_X1  g1009(.A(G41), .B1(new_n1209), .B2(KEYINPUT3), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1197), .B(new_n1208), .C1(G50), .C2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n808), .B1(new_n1211), .B2(new_n796), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1186), .A2(new_n1188), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1214), .B1(new_n1215), .B2(new_n925), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1185), .A2(new_n1216), .ZN(G375));
  OAI21_X1  g1017(.A(new_n353), .B1(new_n834), .B2(new_n759), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1204), .B1(new_n410), .B2(new_n781), .C1(new_n202), .C2(new_n779), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G128), .C2(new_n746), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT124), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n753), .A2(G132), .B1(G137), .B2(new_n763), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(new_n765), .C2(new_n1192), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n762), .A2(new_n827), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n746), .A2(G303), .B1(new_n753), .B2(G294), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n257), .B1(new_n756), .B2(new_n212), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n765), .A2(new_n602), .B1(new_n781), .B2(new_n443), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(G97), .C2(new_n760), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1044), .A2(new_n1225), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1223), .B1(new_n1224), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n809), .B1(new_n1230), .B2(new_n796), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n798), .B2(new_n863), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n333), .B2(new_n1187), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n925), .B(KEYINPUT123), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1179), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1145), .A2(new_n1149), .A3(new_n1140), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n956), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1237), .B2(new_n1150), .ZN(G381));
  NAND3_X1  g1038(.A1(new_n1185), .A2(new_n1155), .A3(new_n1216), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(G381), .A2(G393), .A3(G396), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(G407));
  OAI211_X1 g1043(.A(G407), .B(G213), .C1(G343), .C2(new_n1239), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT125), .Z(G409));
  INV_X1    g1045(.A(G343), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(G213), .A3(G2897), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1155), .B1(new_n1185), .B2(new_n1216), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1234), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n1180), .B2(new_n957), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1215), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(new_n1155), .A3(new_n1213), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1246), .A2(G213), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1247), .B1(new_n1248), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT60), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1151), .B(new_n705), .C1(new_n1256), .C2(new_n1236), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1236), .A2(new_n1256), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1235), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(G384), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1255), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1260), .B(new_n1247), .C1(new_n1248), .C2(new_n1254), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G375), .A2(G378), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1266), .A2(new_n1260), .A3(new_n1253), .A4(new_n1252), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT61), .B1(new_n1267), .B2(KEYINPUT62), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1025), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(G390), .ZN(new_n1272));
  XOR2_X1   g1072(.A(G393), .B(G396), .Z(new_n1273));
  INV_X1    g1073(.A(G390), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT126), .B1(G387), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT126), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1271), .A2(new_n1276), .A3(G390), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1272), .B(new_n1273), .C1(new_n1275), .C2(new_n1277), .ZN(new_n1278));
  OR3_X1    g1078(.A1(new_n1271), .A2(KEYINPUT127), .A3(new_n1274), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1274), .B1(new_n1271), .B2(KEYINPUT127), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1273), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1269), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1283), .B1(new_n1285), .B2(new_n1267), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1262), .A2(KEYINPUT63), .A3(new_n1264), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1284), .A2(new_n1289), .ZN(G405));
  NAND2_X1  g1090(.A1(new_n1266), .A2(new_n1239), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1261), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(new_n1283), .ZN(G402));
endmodule


