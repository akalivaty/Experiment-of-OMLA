

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759;

  AND2_X1 U385 ( .A1(n590), .A2(KEYINPUT44), .ZN(n613) );
  XNOR2_X1 U386 ( .A(n531), .B(KEYINPUT19), .ZN(n568) );
  XNOR2_X1 U387 ( .A(n577), .B(n576), .ZN(n757) );
  INV_X2 U388 ( .A(G116), .ZN(n380) );
  XNOR2_X1 U389 ( .A(n371), .B(n411), .ZN(n673) );
  XNOR2_X1 U390 ( .A(n430), .B(n429), .ZN(n685) );
  XNOR2_X1 U391 ( .A(n511), .B(KEYINPUT4), .ZN(n486) );
  XNOR2_X1 U392 ( .A(G146), .B(G125), .ZN(n491) );
  INV_X2 U393 ( .A(G953), .ZN(n744) );
  NAND2_X1 U394 ( .A1(n495), .A2(n672), .ZN(n531) );
  XNOR2_X1 U395 ( .A(n666), .B(KEYINPUT82), .ZN(n428) );
  XNOR2_X1 U396 ( .A(n493), .B(n492), .ZN(n495) );
  XNOR2_X1 U397 ( .A(n486), .B(n461), .ZN(n740) );
  XNOR2_X1 U398 ( .A(G131), .B(G134), .ZN(n459) );
  OR2_X1 U399 ( .A1(G237), .A2(G902), .ZN(n494) );
  XNOR2_X1 U400 ( .A(n469), .B(KEYINPUT3), .ZN(n485) );
  XNOR2_X1 U401 ( .A(n422), .B(n485), .ZN(n732) );
  XNOR2_X1 U402 ( .A(n484), .B(n501), .ZN(n422) );
  XNOR2_X1 U403 ( .A(n510), .B(n378), .ZN(n484) );
  XNOR2_X1 U404 ( .A(n379), .B(KEYINPUT16), .ZN(n378) );
  NOR2_X1 U405 ( .A1(n709), .A2(n594), .ZN(n584) );
  NAND2_X1 U406 ( .A1(n520), .A2(n538), .ZN(n528) );
  XOR2_X1 U407 ( .A(G122), .B(G104), .Z(n501) );
  XNOR2_X1 U408 ( .A(n491), .B(KEYINPUT10), .ZN(n742) );
  XOR2_X1 U409 ( .A(KEYINPUT11), .B(G140), .Z(n503) );
  XNOR2_X1 U410 ( .A(G113), .B(G143), .ZN(n502) );
  XNOR2_X1 U411 ( .A(n498), .B(n500), .ZN(n398) );
  INV_X1 U412 ( .A(n742), .ZN(n397) );
  XNOR2_X1 U413 ( .A(n536), .B(n535), .ZN(n676) );
  NAND2_X1 U414 ( .A1(n673), .A2(n672), .ZN(n536) );
  BUF_X1 U415 ( .A(n495), .Z(n371) );
  XNOR2_X1 U416 ( .A(n509), .B(n363), .ZN(n537) );
  NOR2_X1 U417 ( .A1(G953), .A2(G237), .ZN(n499) );
  XNOR2_X1 U418 ( .A(n470), .B(n438), .ZN(n437) );
  INV_X1 U419 ( .A(G116), .ZN(n438) );
  XOR2_X1 U420 ( .A(KEYINPUT5), .B(G137), .Z(n470) );
  XNOR2_X1 U421 ( .A(n389), .B(n553), .ZN(n388) );
  XNOR2_X1 U422 ( .A(n740), .B(n462), .ZN(n476) );
  XNOR2_X1 U423 ( .A(n420), .B(n418), .ZN(n417) );
  XNOR2_X1 U424 ( .A(n489), .B(n419), .ZN(n418) );
  XNOR2_X1 U425 ( .A(n486), .B(n421), .ZN(n420) );
  XNOR2_X1 U426 ( .A(n387), .B(KEYINPUT104), .ZN(n578) );
  OR2_X1 U427 ( .A1(n691), .A2(n382), .ZN(n387) );
  AND2_X1 U428 ( .A1(n524), .A2(n523), .ZN(n545) );
  INV_X1 U429 ( .A(KEYINPUT30), .ZN(n369) );
  INV_X1 U430 ( .A(n371), .ZN(n412) );
  XNOR2_X1 U431 ( .A(G478), .B(n519), .ZN(n538) );
  XNOR2_X1 U432 ( .A(n537), .B(n409), .ZN(n520) );
  INV_X1 U433 ( .A(KEYINPUT100), .ZN(n409) );
  XNOR2_X1 U434 ( .A(n433), .B(n367), .ZN(n709) );
  NAND2_X1 U435 ( .A1(n400), .A2(n399), .ZN(n666) );
  NAND2_X1 U436 ( .A1(n659), .A2(KEYINPUT36), .ZN(n399) );
  AND2_X1 U437 ( .A1(n403), .A2(n401), .ZN(n400) );
  NAND2_X1 U438 ( .A1(n618), .A2(KEYINPUT79), .ZN(n394) );
  AND2_X1 U439 ( .A1(n428), .A2(n427), .ZN(n375) );
  INV_X1 U440 ( .A(G110), .ZN(n379) );
  XNOR2_X1 U441 ( .A(G137), .B(G140), .ZN(n475) );
  XOR2_X1 U442 ( .A(KEYINPUT65), .B(G101), .Z(n490) );
  INV_X1 U443 ( .A(n490), .ZN(n421) );
  XNOR2_X1 U444 ( .A(n491), .B(KEYINPUT87), .ZN(n419) );
  NAND2_X1 U445 ( .A1(G234), .A2(G237), .ZN(n453) );
  INV_X1 U446 ( .A(KEYINPUT38), .ZN(n411) );
  AND2_X1 U447 ( .A1(n530), .A2(n407), .ZN(n406) );
  INV_X1 U448 ( .A(n531), .ZN(n407) );
  INV_X1 U449 ( .A(KEYINPUT36), .ZN(n405) );
  XNOR2_X1 U450 ( .A(n532), .B(KEYINPUT1), .ZN(n691) );
  XNOR2_X1 U451 ( .A(n482), .B(G469), .ZN(n532) );
  NOR2_X1 U452 ( .A1(G902), .A2(n716), .ZN(n482) );
  XNOR2_X1 U453 ( .A(n450), .B(n364), .ZN(n429) );
  OR2_X1 U454 ( .A1(n725), .A2(G902), .ZN(n430) );
  NOR2_X2 U455 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U456 ( .A(G119), .B(G110), .ZN(n440) );
  XNOR2_X1 U457 ( .A(n377), .B(KEYINPUT101), .ZN(n376) );
  INV_X1 U458 ( .A(G122), .ZN(n377) );
  XNOR2_X1 U459 ( .A(n507), .B(n506), .ZN(n624) );
  XNOR2_X1 U460 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n507) );
  INV_X1 U462 ( .A(KEYINPUT73), .ZN(n385) );
  XNOR2_X1 U463 ( .A(G104), .B(G107), .ZN(n477) );
  XOR2_X1 U464 ( .A(KEYINPUT91), .B(G110), .Z(n478) );
  NOR2_X1 U465 ( .A1(n676), .A2(n675), .ZN(n540) );
  AND2_X1 U466 ( .A1(n406), .A2(n405), .ZN(n404) );
  AND2_X1 U467 ( .A1(n402), .A2(n533), .ZN(n401) );
  OR2_X1 U468 ( .A1(n406), .A2(n405), .ZN(n402) );
  XNOR2_X1 U469 ( .A(KEYINPUT22), .B(KEYINPUT70), .ZN(n573) );
  BUF_X1 U470 ( .A(n685), .Z(n382) );
  INV_X1 U471 ( .A(KEYINPUT6), .ZN(n434) );
  XNOR2_X1 U472 ( .A(n476), .B(n435), .ZN(n638) );
  XNOR2_X1 U473 ( .A(n485), .B(n436), .ZN(n435) );
  XNOR2_X1 U474 ( .A(n437), .B(n362), .ZN(n436) );
  XNOR2_X1 U475 ( .A(n476), .B(n386), .ZN(n716) );
  XNOR2_X1 U476 ( .A(n481), .B(n739), .ZN(n386) );
  XNOR2_X1 U477 ( .A(n479), .B(n384), .ZN(n481) );
  XNOR2_X1 U478 ( .A(n480), .B(n385), .ZN(n384) );
  XNOR2_X1 U479 ( .A(n632), .B(KEYINPUT54), .ZN(n633) );
  NAND2_X1 U480 ( .A1(n557), .A2(n412), .ZN(n558) );
  XNOR2_X1 U481 ( .A(n381), .B(n548), .ZN(n754) );
  INV_X1 U482 ( .A(KEYINPUT35), .ZN(n432) );
  XNOR2_X1 U483 ( .A(n416), .B(n414), .ZN(n663) );
  XNOR2_X1 U484 ( .A(n415), .B(KEYINPUT31), .ZN(n414) );
  INV_X1 U485 ( .A(KEYINPUT95), .ZN(n415) );
  NOR2_X1 U486 ( .A1(n525), .A2(n412), .ZN(n653) );
  INV_X1 U487 ( .A(KEYINPUT107), .ZN(n408) );
  XOR2_X1 U488 ( .A(G902), .B(KEYINPUT15), .Z(n618) );
  AND2_X1 U489 ( .A1(n499), .A2(G210), .ZN(n362) );
  XNOR2_X1 U490 ( .A(n528), .B(n408), .ZN(n659) );
  XOR2_X1 U491 ( .A(KEYINPUT99), .B(n508), .Z(n363) );
  XOR2_X1 U492 ( .A(KEYINPUT72), .B(KEYINPUT25), .Z(n364) );
  XOR2_X1 U493 ( .A(n445), .B(n444), .Z(n365) );
  NOR2_X1 U494 ( .A1(n552), .A2(n551), .ZN(n366) );
  XOR2_X1 U495 ( .A(KEYINPUT84), .B(KEYINPUT33), .Z(n367) );
  XOR2_X1 U496 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n368) );
  INV_X1 U497 ( .A(KEYINPUT79), .ZN(n413) );
  NAND2_X1 U498 ( .A1(n410), .A2(n589), .ZN(n590) );
  NOR2_X2 U499 ( .A1(n757), .A2(n756), .ZN(n410) );
  INV_X1 U500 ( .A(n616), .ZN(n738) );
  NAND2_X1 U501 ( .A1(n391), .A2(n616), .ZN(n390) );
  AND2_X2 U502 ( .A1(n561), .A2(n670), .ZN(n616) );
  XNOR2_X1 U503 ( .A(n546), .B(KEYINPUT39), .ZN(n560) );
  XNOR2_X1 U504 ( .A(n370), .B(n369), .ZN(n524) );
  NAND2_X1 U505 ( .A1(n688), .A2(n672), .ZN(n370) );
  NAND2_X1 U506 ( .A1(n424), .A2(n375), .ZN(n389) );
  XNOR2_X1 U507 ( .A(n732), .B(n417), .ZN(n631) );
  AND2_X1 U508 ( .A1(n373), .A2(n713), .ZN(G66) );
  XNOR2_X2 U509 ( .A(n614), .B(KEYINPUT45), .ZN(n729) );
  NAND2_X1 U510 ( .A1(n372), .A2(n426), .ZN(n425) );
  INV_X1 U511 ( .A(n753), .ZN(n372) );
  XNOR2_X1 U512 ( .A(n544), .B(n543), .ZN(n753) );
  XNOR2_X1 U513 ( .A(n724), .B(n374), .ZN(n373) );
  INV_X1 U514 ( .A(n725), .ZN(n374) );
  NOR2_X1 U515 ( .A1(n729), .A2(n394), .ZN(n393) );
  XNOR2_X1 U516 ( .A(n511), .B(n376), .ZN(n512) );
  NOR2_X1 U517 ( .A1(n729), .A2(n617), .ZN(n391) );
  XNOR2_X2 U518 ( .A(n380), .B(G107), .ZN(n510) );
  NAND2_X1 U519 ( .A1(n560), .A2(n547), .ZN(n381) );
  NAND2_X1 U520 ( .A1(n759), .A2(n388), .ZN(n559) );
  XNOR2_X1 U521 ( .A(n448), .B(n447), .ZN(n725) );
  XNOR2_X1 U522 ( .A(n425), .B(n368), .ZN(n424) );
  INV_X1 U523 ( .A(n423), .ZN(n621) );
  NAND2_X1 U524 ( .A1(n423), .A2(KEYINPUT76), .ZN(n671) );
  XNOR2_X1 U525 ( .A(n603), .B(KEYINPUT105), .ZN(n575) );
  OR2_X2 U526 ( .A1(n581), .A2(n533), .ZN(n603) );
  NAND2_X1 U527 ( .A1(n383), .A2(n585), .ZN(n586) );
  XNOR2_X1 U528 ( .A(n584), .B(KEYINPUT34), .ZN(n383) );
  NAND2_X1 U529 ( .A1(n390), .A2(n413), .ZN(n395) );
  NAND2_X1 U530 ( .A1(n395), .A2(n392), .ZN(n396) );
  NAND2_X1 U531 ( .A1(n616), .A2(n393), .ZN(n392) );
  NAND2_X1 U532 ( .A1(n396), .A2(n620), .ZN(n623) );
  NAND2_X1 U533 ( .A1(n655), .A2(n530), .ZN(n554) );
  NAND2_X1 U534 ( .A1(n655), .A2(n404), .ZN(n403) );
  NAND2_X1 U535 ( .A1(n410), .A2(n592), .ZN(n611) );
  NOR2_X1 U536 ( .A1(n594), .A2(n695), .ZN(n416) );
  XNOR2_X2 U537 ( .A(n569), .B(KEYINPUT0), .ZN(n594) );
  NAND2_X1 U538 ( .A1(n615), .A2(n616), .ZN(n423) );
  INV_X1 U539 ( .A(n754), .ZN(n426) );
  NOR2_X1 U540 ( .A1(n534), .A2(n366), .ZN(n427) );
  INV_X1 U541 ( .A(n755), .ZN(n606) );
  AND2_X1 U542 ( .A1(n431), .A2(n591), .ZN(n592) );
  XNOR2_X1 U543 ( .A(n755), .B(KEYINPUT66), .ZN(n431) );
  XNOR2_X2 U544 ( .A(n586), .B(n432), .ZN(n755) );
  NAND2_X1 U545 ( .A1(n593), .A2(n600), .ZN(n433) );
  XNOR2_X1 U546 ( .A(n688), .B(n434), .ZN(n600) );
  XNOR2_X2 U547 ( .A(n472), .B(n471), .ZN(n688) );
  XNOR2_X1 U548 ( .A(n718), .B(n717), .ZN(n719) );
  AND2_X1 U549 ( .A1(n596), .A2(n522), .ZN(n523) );
  NOR2_X1 U550 ( .A1(n631), .A2(n618), .ZN(n493) );
  NOR2_X1 U551 ( .A1(n688), .A2(n382), .ZN(n439) );
  INV_X1 U552 ( .A(n691), .ZN(n533) );
  INV_X1 U553 ( .A(KEYINPUT48), .ZN(n553) );
  INV_X1 U554 ( .A(KEYINPUT111), .ZN(n535) );
  XNOR2_X1 U555 ( .A(n446), .B(n365), .ZN(n447) );
  BUF_X1 U556 ( .A(n683), .Z(n708) );
  XNOR2_X1 U557 ( .A(n574), .B(n573), .ZN(n581) );
  INV_X1 U558 ( .A(KEYINPUT60), .ZN(n629) );
  INV_X1 U559 ( .A(n618), .ZN(n617) );
  XOR2_X1 U560 ( .A(KEYINPUT28), .B(KEYINPUT109), .Z(n474) );
  XNOR2_X1 U561 ( .A(n742), .B(n475), .ZN(n441) );
  XNOR2_X1 U562 ( .A(n441), .B(n440), .ZN(n448) );
  XOR2_X1 U563 ( .A(KEYINPUT78), .B(KEYINPUT8), .Z(n443) );
  NAND2_X1 U564 ( .A1(G234), .A2(n744), .ZN(n442) );
  XNOR2_X1 U565 ( .A(n443), .B(n442), .ZN(n514) );
  NAND2_X1 U566 ( .A1(G221), .A2(n514), .ZN(n446) );
  XOR2_X1 U567 ( .A(KEYINPUT92), .B(KEYINPUT24), .Z(n445) );
  XNOR2_X1 U568 ( .A(G128), .B(KEYINPUT23), .ZN(n444) );
  NAND2_X1 U569 ( .A1(G234), .A2(n617), .ZN(n449) );
  XNOR2_X1 U570 ( .A(KEYINPUT20), .B(n449), .ZN(n451) );
  NAND2_X1 U571 ( .A1(n451), .A2(G217), .ZN(n450) );
  NAND2_X1 U572 ( .A1(n451), .A2(G221), .ZN(n452) );
  XNOR2_X1 U573 ( .A(n452), .B(KEYINPUT21), .ZN(n570) );
  NOR2_X1 U574 ( .A1(n685), .A2(n570), .ZN(n458) );
  XNOR2_X1 U575 ( .A(n453), .B(KEYINPUT14), .ZN(n455) );
  NAND2_X1 U576 ( .A1(G902), .A2(n455), .ZN(n562) );
  NOR2_X1 U577 ( .A1(G900), .A2(n562), .ZN(n454) );
  NAND2_X1 U578 ( .A1(G953), .A2(n454), .ZN(n457) );
  NAND2_X1 U579 ( .A1(G952), .A2(n455), .ZN(n456) );
  XOR2_X1 U580 ( .A(KEYINPUT88), .B(n456), .Z(n702) );
  NAND2_X1 U581 ( .A1(n744), .A2(n702), .ZN(n565) );
  NAND2_X1 U582 ( .A1(n457), .A2(n565), .ZN(n522) );
  AND2_X1 U583 ( .A1(n458), .A2(n522), .ZN(n529) );
  XNOR2_X2 U584 ( .A(G143), .B(G128), .ZN(n511) );
  INV_X1 U585 ( .A(n459), .ZN(n460) );
  XNOR2_X1 U586 ( .A(KEYINPUT68), .B(n460), .ZN(n461) );
  XNOR2_X1 U587 ( .A(n490), .B(G146), .ZN(n462) );
  XNOR2_X1 U588 ( .A(G119), .B(G113), .ZN(n468) );
  INV_X1 U589 ( .A(KEYINPUT86), .ZN(n463) );
  NAND2_X1 U590 ( .A1(KEYINPUT69), .A2(n463), .ZN(n466) );
  INV_X1 U591 ( .A(KEYINPUT69), .ZN(n464) );
  NAND2_X1 U592 ( .A1(n464), .A2(KEYINPUT86), .ZN(n465) );
  NAND2_X1 U593 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U594 ( .A(n468), .B(n467), .ZN(n469) );
  NOR2_X1 U595 ( .A1(n638), .A2(G902), .ZN(n472) );
  XNOR2_X1 U596 ( .A(G472), .B(KEYINPUT93), .ZN(n471) );
  NAND2_X1 U597 ( .A1(n529), .A2(n688), .ZN(n473) );
  XNOR2_X1 U598 ( .A(n474), .B(n473), .ZN(n483) );
  XNOR2_X1 U599 ( .A(KEYINPUT90), .B(n475), .ZN(n739) );
  XNOR2_X1 U600 ( .A(n478), .B(n477), .ZN(n479) );
  NAND2_X1 U601 ( .A1(G227), .A2(n744), .ZN(n480) );
  NOR2_X1 U602 ( .A1(n483), .A2(n532), .ZN(n541) );
  XOR2_X1 U603 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n488) );
  NAND2_X1 U604 ( .A1(G224), .A2(n744), .ZN(n487) );
  XNOR2_X1 U605 ( .A(n488), .B(n487), .ZN(n489) );
  NAND2_X1 U606 ( .A1(G210), .A2(n494), .ZN(n492) );
  NAND2_X1 U607 ( .A1(G214), .A2(n494), .ZN(n672) );
  NAND2_X1 U608 ( .A1(n541), .A2(n568), .ZN(n552) );
  INV_X1 U609 ( .A(n552), .ZN(n656) );
  XOR2_X1 U610 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n497) );
  XNOR2_X1 U611 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n496) );
  XNOR2_X1 U612 ( .A(n497), .B(n496), .ZN(n498) );
  NAND2_X1 U613 ( .A1(G214), .A2(n499), .ZN(n500) );
  XNOR2_X1 U614 ( .A(G131), .B(n501), .ZN(n505) );
  XNOR2_X1 U615 ( .A(n503), .B(n502), .ZN(n504) );
  NOR2_X1 U616 ( .A1(n624), .A2(G902), .ZN(n509) );
  XOR2_X1 U617 ( .A(G475), .B(KEYINPUT13), .Z(n508) );
  XNOR2_X1 U618 ( .A(n510), .B(G134), .ZN(n513) );
  XNOR2_X1 U619 ( .A(n513), .B(n512), .ZN(n518) );
  XOR2_X1 U620 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n516) );
  NAND2_X1 U621 ( .A1(G217), .A2(n514), .ZN(n515) );
  XNOR2_X1 U622 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U623 ( .A(n518), .B(n517), .ZN(n721) );
  NOR2_X1 U624 ( .A1(G902), .A2(n721), .ZN(n519) );
  NOR2_X1 U625 ( .A1(n520), .A2(n538), .ZN(n649) );
  INV_X1 U626 ( .A(n528), .ZN(n547) );
  NOR2_X1 U627 ( .A1(n649), .A2(n547), .ZN(n677) );
  INV_X1 U628 ( .A(n677), .ZN(n598) );
  NAND2_X1 U629 ( .A1(n656), .A2(n598), .ZN(n521) );
  NAND2_X1 U630 ( .A1(KEYINPUT47), .A2(n521), .ZN(n527) );
  INV_X1 U631 ( .A(n570), .ZN(n684) );
  NAND2_X1 U632 ( .A1(n685), .A2(n684), .ZN(n690) );
  NOR2_X1 U633 ( .A1(n532), .A2(n690), .ZN(n596) );
  NOR2_X1 U634 ( .A1(n537), .A2(n538), .ZN(n585) );
  NAND2_X1 U635 ( .A1(n545), .A2(n585), .ZN(n525) );
  XNOR2_X1 U636 ( .A(KEYINPUT77), .B(n653), .ZN(n526) );
  NAND2_X1 U637 ( .A1(n527), .A2(n526), .ZN(n534) );
  INV_X1 U638 ( .A(n659), .ZN(n655) );
  AND2_X1 U639 ( .A1(n529), .A2(n600), .ZN(n530) );
  NAND2_X1 U640 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U641 ( .A(n539), .B(KEYINPUT102), .ZN(n675) );
  XNOR2_X1 U642 ( .A(n540), .B(KEYINPUT41), .ZN(n683) );
  INV_X1 U643 ( .A(n541), .ZN(n542) );
  NOR2_X1 U644 ( .A1(n683), .A2(n542), .ZN(n544) );
  XNOR2_X1 U645 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n543) );
  XOR2_X1 U646 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n548) );
  NAND2_X1 U647 ( .A1(n545), .A2(n673), .ZN(n546) );
  XOR2_X1 U648 ( .A(KEYINPUT47), .B(KEYINPUT67), .Z(n549) );
  NOR2_X1 U649 ( .A1(n677), .A2(n549), .ZN(n550) );
  XNOR2_X1 U650 ( .A(n550), .B(KEYINPUT71), .ZN(n551) );
  NOR2_X1 U651 ( .A1(n554), .A2(n533), .ZN(n555) );
  NAND2_X1 U652 ( .A1(n555), .A2(n672), .ZN(n556) );
  XNOR2_X1 U653 ( .A(n556), .B(KEYINPUT43), .ZN(n557) );
  XNOR2_X1 U654 ( .A(KEYINPUT108), .B(n558), .ZN(n759) );
  XNOR2_X1 U655 ( .A(n559), .B(KEYINPUT81), .ZN(n561) );
  NAND2_X1 U656 ( .A1(n560), .A2(n649), .ZN(n670) );
  INV_X1 U657 ( .A(n562), .ZN(n563) );
  NOR2_X1 U658 ( .A1(G898), .A2(n744), .ZN(n734) );
  NAND2_X1 U659 ( .A1(n563), .A2(n734), .ZN(n564) );
  NAND2_X1 U660 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U661 ( .A(KEYINPUT89), .B(n566), .Z(n567) );
  NAND2_X1 U662 ( .A1(n568), .A2(n567), .ZN(n569) );
  INV_X1 U663 ( .A(n594), .ZN(n572) );
  NOR2_X1 U664 ( .A1(n570), .A2(n675), .ZN(n571) );
  NAND2_X1 U665 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U666 ( .A1(n575), .A2(n439), .ZN(n577) );
  INV_X1 U667 ( .A(KEYINPUT106), .ZN(n576) );
  NOR2_X1 U668 ( .A1(n600), .A2(n578), .ZN(n579) );
  XNOR2_X1 U669 ( .A(n579), .B(KEYINPUT75), .ZN(n580) );
  NOR2_X1 U670 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U671 ( .A(n582), .B(KEYINPUT74), .ZN(n583) );
  XNOR2_X1 U672 ( .A(n583), .B(KEYINPUT32), .ZN(n756) );
  NOR2_X1 U673 ( .A1(n691), .A2(n690), .ZN(n593) );
  NOR2_X1 U674 ( .A1(KEYINPUT83), .A2(n755), .ZN(n588) );
  INV_X1 U675 ( .A(KEYINPUT66), .ZN(n587) );
  NOR2_X1 U676 ( .A1(n588), .A2(n587), .ZN(n589) );
  INV_X1 U677 ( .A(KEYINPUT44), .ZN(n591) );
  NAND2_X1 U678 ( .A1(n688), .A2(n593), .ZN(n695) );
  NOR2_X1 U679 ( .A1(n688), .A2(n594), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U681 ( .A(KEYINPUT94), .B(n597), .ZN(n645) );
  NAND2_X1 U682 ( .A1(n663), .A2(n645), .ZN(n599) );
  NAND2_X1 U683 ( .A1(n599), .A2(n598), .ZN(n604) );
  INV_X1 U684 ( .A(n382), .ZN(n601) );
  OR2_X1 U685 ( .A1(n601), .A2(n600), .ZN(n602) );
  OR2_X1 U686 ( .A1(n603), .A2(n602), .ZN(n643) );
  NAND2_X1 U687 ( .A1(n604), .A2(n643), .ZN(n605) );
  XNOR2_X1 U688 ( .A(KEYINPUT103), .B(n605), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n606), .A2(KEYINPUT44), .ZN(n607) );
  NAND2_X1 U690 ( .A1(n607), .A2(KEYINPUT83), .ZN(n608) );
  AND2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n611), .A2(n610), .ZN(n612) );
  INV_X1 U693 ( .A(n729), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n618), .B(KEYINPUT80), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n619), .A2(KEYINPUT2), .ZN(n620) );
  NAND2_X1 U696 ( .A1(KEYINPUT2), .A2(n621), .ZN(n622) );
  AND2_X2 U697 ( .A1(n623), .A2(n622), .ZN(n714) );
  NAND2_X1 U698 ( .A1(G475), .A2(n714), .ZN(n626) );
  XNOR2_X1 U699 ( .A(n624), .B(KEYINPUT59), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n626), .B(n625), .ZN(n628) );
  NOR2_X1 U701 ( .A1(G952), .A2(n744), .ZN(n627) );
  XNOR2_X1 U702 ( .A(KEYINPUT85), .B(n627), .ZN(n713) );
  NAND2_X1 U703 ( .A1(n628), .A2(n713), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n630), .B(n629), .ZN(G60) );
  NAND2_X1 U705 ( .A1(G210), .A2(n714), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n631), .B(KEYINPUT55), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n635), .A2(n713), .ZN(n637) );
  INV_X1 U709 ( .A(KEYINPUT56), .ZN(n636) );
  XNOR2_X1 U710 ( .A(n637), .B(n636), .ZN(G51) );
  NAND2_X1 U711 ( .A1(n714), .A2(G472), .ZN(n640) );
  XOR2_X1 U712 ( .A(n638), .B(KEYINPUT62), .Z(n639) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(n641) );
  NAND2_X1 U714 ( .A1(n641), .A2(n713), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n642), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U716 ( .A(G101), .B(n643), .ZN(G3) );
  NOR2_X1 U717 ( .A1(n645), .A2(n659), .ZN(n644) );
  XOR2_X1 U718 ( .A(G104), .B(n644), .Z(G6) );
  INV_X1 U719 ( .A(n649), .ZN(n664) );
  NOR2_X1 U720 ( .A1(n645), .A2(n664), .ZN(n647) );
  XNOR2_X1 U721 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U723 ( .A(G107), .B(n648), .ZN(G9) );
  XOR2_X1 U724 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n651) );
  NAND2_X1 U725 ( .A1(n656), .A2(n649), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U727 ( .A(G128), .B(n652), .ZN(G30) );
  XNOR2_X1 U728 ( .A(G143), .B(n653), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(KEYINPUT115), .ZN(G45) );
  NAND2_X1 U730 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n657), .B(KEYINPUT116), .ZN(n658) );
  XNOR2_X1 U732 ( .A(G146), .B(n658), .ZN(G48) );
  NOR2_X1 U733 ( .A1(n659), .A2(n663), .ZN(n661) );
  XNOR2_X1 U734 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U736 ( .A(G113), .B(n662), .ZN(G15) );
  NOR2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U738 ( .A(G116), .B(n665), .Z(G18) );
  XOR2_X1 U739 ( .A(KEYINPUT37), .B(KEYINPUT119), .Z(n669) );
  INV_X1 U740 ( .A(n666), .ZN(n667) );
  XNOR2_X1 U741 ( .A(G125), .B(n667), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n669), .B(n668), .ZN(G27) );
  XNOR2_X1 U743 ( .A(G134), .B(n670), .ZN(G36) );
  XNOR2_X1 U744 ( .A(n671), .B(KEYINPUT2), .ZN(n707) );
  NOR2_X1 U745 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U749 ( .A(KEYINPUT121), .B(n680), .Z(n681) );
  NOR2_X1 U750 ( .A1(n709), .A2(n681), .ZN(n682) );
  XNOR2_X1 U751 ( .A(n682), .B(KEYINPUT122), .ZN(n700) );
  NOR2_X1 U752 ( .A1(n382), .A2(n684), .ZN(n686) );
  XOR2_X1 U753 ( .A(KEYINPUT49), .B(n686), .Z(n687) );
  NOR2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U755 ( .A(n689), .B(KEYINPUT120), .ZN(n694) );
  NAND2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U757 ( .A(KEYINPUT50), .B(n692), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U760 ( .A(KEYINPUT51), .B(n697), .ZN(n698) );
  NOR2_X1 U761 ( .A1(n708), .A2(n698), .ZN(n699) );
  NOR2_X1 U762 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U763 ( .A(KEYINPUT52), .B(n701), .Z(n703) );
  NAND2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U765 ( .A(KEYINPUT123), .B(n704), .ZN(n705) );
  NOR2_X1 U766 ( .A1(G953), .A2(n705), .ZN(n706) );
  NAND2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n711) );
  NOR2_X1 U768 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U770 ( .A(KEYINPUT53), .B(n712), .ZN(G75) );
  INV_X1 U771 ( .A(n713), .ZN(n726) );
  BUF_X2 U772 ( .A(n714), .Z(n723) );
  NAND2_X1 U773 ( .A1(n723), .A2(G469), .ZN(n718) );
  XOR2_X1 U774 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n715) );
  XNOR2_X1 U775 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U776 ( .A1(n726), .A2(n719), .ZN(G54) );
  NAND2_X1 U777 ( .A1(G478), .A2(n723), .ZN(n720) );
  XNOR2_X1 U778 ( .A(n720), .B(n721), .ZN(n722) );
  NOR2_X1 U779 ( .A1(n726), .A2(n722), .ZN(G63) );
  NAND2_X1 U780 ( .A1(G217), .A2(n723), .ZN(n724) );
  NAND2_X1 U781 ( .A1(G953), .A2(G224), .ZN(n727) );
  XNOR2_X1 U782 ( .A(KEYINPUT61), .B(n727), .ZN(n728) );
  AND2_X1 U783 ( .A1(n728), .A2(G898), .ZN(n731) );
  NOR2_X1 U784 ( .A1(n729), .A2(G953), .ZN(n730) );
  NOR2_X1 U785 ( .A1(n731), .A2(n730), .ZN(n737) );
  XOR2_X1 U786 ( .A(n732), .B(G101), .Z(n733) );
  NOR2_X1 U787 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U788 ( .A(KEYINPUT124), .B(n735), .Z(n736) );
  XNOR2_X1 U789 ( .A(n737), .B(n736), .ZN(G69) );
  XNOR2_X1 U790 ( .A(KEYINPUT125), .B(n738), .ZN(n743) );
  XOR2_X1 U791 ( .A(n740), .B(n739), .Z(n741) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(n747) );
  XNOR2_X1 U793 ( .A(n743), .B(n747), .ZN(n745) );
  NAND2_X1 U794 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U795 ( .A(n746), .B(KEYINPUT126), .ZN(n752) );
  XNOR2_X1 U796 ( .A(KEYINPUT127), .B(n747), .ZN(n748) );
  XNOR2_X1 U797 ( .A(G227), .B(n748), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n749), .A2(G900), .ZN(n750) );
  NAND2_X1 U799 ( .A1(n750), .A2(G953), .ZN(n751) );
  NAND2_X1 U800 ( .A1(n752), .A2(n751), .ZN(G72) );
  XOR2_X1 U801 ( .A(G137), .B(n753), .Z(G39) );
  XOR2_X1 U802 ( .A(n754), .B(G131), .Z(G33) );
  XNOR2_X1 U803 ( .A(n755), .B(G122), .ZN(G24) );
  XOR2_X1 U804 ( .A(G119), .B(n756), .Z(G21) );
  XNOR2_X1 U805 ( .A(G110), .B(KEYINPUT113), .ZN(n758) );
  XNOR2_X1 U806 ( .A(n758), .B(n757), .ZN(G12) );
  XNOR2_X1 U807 ( .A(G140), .B(n759), .ZN(G42) );
endmodule

