

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U321 ( .A(KEYINPUT116), .B(n461), .ZN(n542) );
  NOR2_X1 U322 ( .A1(n508), .A2(n460), .ZN(n461) );
  XNOR2_X1 U323 ( .A(n289), .B(KEYINPUT115), .ZN(n460) );
  NOR2_X1 U324 ( .A1(n563), .A2(n412), .ZN(n413) );
  XNOR2_X1 U325 ( .A(n387), .B(n290), .ZN(n389) );
  NOR2_X1 U326 ( .A1(n557), .A2(n512), .ZN(n409) );
  XNOR2_X1 U327 ( .A(KEYINPUT112), .B(KEYINPUT45), .ZN(n290) );
  XNOR2_X1 U328 ( .A(n386), .B(n423), .ZN(n480) );
  XOR2_X1 U329 ( .A(n384), .B(n383), .Z(n386) );
  XOR2_X1 U330 ( .A(n406), .B(n405), .Z(n571) );
  XOR2_X1 U331 ( .A(n369), .B(n368), .Z(n481) );
  XNOR2_X1 U332 ( .A(G15GAT), .B(G1GAT), .ZN(n371) );
  INV_X2 U333 ( .A(n559), .ZN(n562) );
  AND2_X1 U334 ( .A1(n545), .A2(n505), .ZN(n289) );
  NAND2_X1 U335 ( .A1(n566), .A2(n433), .ZN(n434) );
  XNOR2_X1 U336 ( .A(n432), .B(KEYINPUT54), .ZN(n566) );
  XNOR2_X1 U337 ( .A(n394), .B(n359), .ZN(n367) );
  XOR2_X1 U338 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n353) );
  BUF_X1 U339 ( .A(n580), .Z(n291) );
  XNOR2_X1 U340 ( .A(n563), .B(KEYINPUT36), .ZN(n580) );
  XNOR2_X1 U341 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n417) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G190GAT), .ZN(n355) );
  XNOR2_X1 U343 ( .A(n309), .B(n308), .ZN(n576) );
  XNOR2_X1 U344 ( .A(n292), .B(n307), .ZN(n308) );
  XOR2_X1 U345 ( .A(KEYINPUT41), .B(n576), .Z(n551) );
  XNOR2_X1 U346 ( .A(n355), .B(KEYINPUT79), .ZN(n419) );
  XOR2_X1 U347 ( .A(n299), .B(n298), .Z(n292) );
  XNOR2_X1 U348 ( .A(n420), .B(n306), .ZN(n307) );
  INV_X1 U349 ( .A(G134GAT), .ZN(n462) );
  XNOR2_X1 U350 ( .A(n454), .B(G176GAT), .ZN(n455) );
  XNOR2_X1 U351 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U352 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  XOR2_X1 U353 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n294) );
  XNOR2_X1 U354 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n293) );
  XOR2_X1 U355 ( .A(n294), .B(n293), .Z(n309) );
  XOR2_X1 U356 ( .A(KEYINPUT71), .B(KEYINPUT75), .Z(n296) );
  XNOR2_X1 U357 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n295) );
  XNOR2_X1 U358 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U359 ( .A(G99GAT), .B(G85GAT), .Z(n356) );
  XNOR2_X1 U360 ( .A(n297), .B(n356), .ZN(n299) );
  AND2_X1 U361 ( .A1(G230GAT), .A2(G233GAT), .ZN(n298) );
  XOR2_X1 U362 ( .A(KEYINPUT73), .B(G64GAT), .Z(n301) );
  XNOR2_X1 U363 ( .A(G176GAT), .B(G92GAT), .ZN(n300) );
  XNOR2_X1 U364 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U365 ( .A(G204GAT), .B(n302), .Z(n420) );
  XNOR2_X1 U366 ( .A(G106GAT), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U367 ( .A(n303), .B(G148GAT), .ZN(n332) );
  XOR2_X1 U368 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n305) );
  XNOR2_X1 U369 ( .A(G71GAT), .B(G57GAT), .ZN(n304) );
  XNOR2_X1 U370 ( .A(n305), .B(n304), .ZN(n384) );
  XNOR2_X1 U371 ( .A(n332), .B(n384), .ZN(n306) );
  INV_X1 U372 ( .A(n551), .ZN(n512) );
  XOR2_X1 U373 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n435) );
  XOR2_X1 U374 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n311) );
  XNOR2_X1 U375 ( .A(G141GAT), .B(KEYINPUT91), .ZN(n310) );
  XNOR2_X1 U376 ( .A(n311), .B(n310), .ZN(n341) );
  XOR2_X1 U377 ( .A(G85GAT), .B(n341), .Z(n313) );
  NAND2_X1 U378 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U379 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U380 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n315) );
  XNOR2_X1 U381 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n314) );
  XNOR2_X1 U382 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U383 ( .A(n317), .B(n316), .Z(n323) );
  XNOR2_X1 U384 ( .A(G127GAT), .B(G134GAT), .ZN(n318) );
  XNOR2_X1 U385 ( .A(n318), .B(KEYINPUT0), .ZN(n319) );
  XOR2_X1 U386 ( .A(n319), .B(KEYINPUT83), .Z(n321) );
  XNOR2_X1 U387 ( .A(G113GAT), .B(G120GAT), .ZN(n320) );
  XNOR2_X1 U388 ( .A(n321), .B(n320), .ZN(n440) );
  XNOR2_X1 U389 ( .A(G29GAT), .B(n440), .ZN(n322) );
  XNOR2_X1 U390 ( .A(n323), .B(n322), .ZN(n331) );
  XOR2_X1 U391 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n325) );
  XNOR2_X1 U392 ( .A(G1GAT), .B(KEYINPUT95), .ZN(n324) );
  XNOR2_X1 U393 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U394 ( .A(G57GAT), .B(G155GAT), .Z(n327) );
  XNOR2_X1 U395 ( .A(G162GAT), .B(G148GAT), .ZN(n326) );
  XNOR2_X1 U396 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U397 ( .A(n329), .B(n328), .Z(n330) );
  XOR2_X1 U398 ( .A(n331), .B(n330), .Z(n567) );
  XOR2_X1 U399 ( .A(G50GAT), .B(G162GAT), .Z(n363) );
  XOR2_X1 U400 ( .A(n363), .B(n332), .Z(n334) );
  NAND2_X1 U401 ( .A1(G228GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U402 ( .A(n334), .B(n333), .ZN(n345) );
  XOR2_X1 U403 ( .A(G204GAT), .B(G211GAT), .Z(n336) );
  XNOR2_X1 U404 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n335) );
  XNOR2_X1 U405 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U406 ( .A(n337), .B(KEYINPUT92), .Z(n339) );
  XOR2_X1 U407 ( .A(G22GAT), .B(G155GAT), .Z(n370) );
  XNOR2_X1 U408 ( .A(n370), .B(KEYINPUT24), .ZN(n338) );
  XNOR2_X1 U409 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U410 ( .A(n340), .B(KEYINPUT94), .Z(n343) );
  XNOR2_X1 U411 ( .A(n341), .B(KEYINPUT22), .ZN(n342) );
  XNOR2_X1 U412 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U413 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U414 ( .A(KEYINPUT21), .B(G218GAT), .Z(n347) );
  XNOR2_X1 U415 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n346) );
  XNOR2_X1 U416 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U417 ( .A(G197GAT), .B(n348), .Z(n428) );
  XOR2_X1 U418 ( .A(n349), .B(n428), .Z(n468) );
  AND2_X1 U419 ( .A1(n567), .A2(n468), .ZN(n433) );
  XOR2_X1 U420 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n351) );
  XNOR2_X1 U421 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n350) );
  XNOR2_X1 U422 ( .A(n351), .B(n350), .ZN(n369) );
  XNOR2_X1 U423 ( .A(G43GAT), .B(G29GAT), .ZN(n352) );
  XNOR2_X1 U424 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U425 ( .A(KEYINPUT68), .B(n354), .Z(n394) );
  XOR2_X1 U426 ( .A(n356), .B(n419), .Z(n358) );
  NAND2_X1 U427 ( .A1(G232GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U429 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n361) );
  XNOR2_X1 U430 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n360) );
  XNOR2_X1 U431 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U432 ( .A(n362), .B(G106GAT), .Z(n365) );
  XNOR2_X1 U433 ( .A(G218GAT), .B(n363), .ZN(n364) );
  XNOR2_X1 U434 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n368) );
  INV_X1 U436 ( .A(n481), .ZN(n563) );
  XOR2_X1 U437 ( .A(n370), .B(G78GAT), .Z(n373) );
  XNOR2_X1 U438 ( .A(n371), .B(KEYINPUT69), .ZN(n393) );
  XNOR2_X1 U439 ( .A(n393), .B(G127GAT), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n372), .B(n373), .ZN(n377) );
  XOR2_X1 U441 ( .A(KEYINPUT14), .B(G64GAT), .Z(n375) );
  NAND2_X1 U442 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U444 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U445 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n379) );
  XNOR2_X1 U446 ( .A(KEYINPUT82), .B(KEYINPUT15), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U448 ( .A(n380), .B(KEYINPUT81), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U450 ( .A(G8GAT), .B(G183GAT), .Z(n385) );
  XOR2_X1 U451 ( .A(G211GAT), .B(n385), .Z(n423) );
  NAND2_X1 U452 ( .A1(n580), .A2(n480), .ZN(n387) );
  NOR2_X1 U453 ( .A1(n389), .A2(n576), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n390), .B(KEYINPUT113), .ZN(n407) );
  XOR2_X1 U455 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n392) );
  XNOR2_X1 U456 ( .A(G197GAT), .B(G8GAT), .ZN(n391) );
  XNOR2_X1 U457 ( .A(n392), .B(n391), .ZN(n398) );
  XOR2_X1 U458 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n396) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n406) );
  NAND2_X1 U462 ( .A1(G229GAT), .A2(G233GAT), .ZN(n404) );
  XOR2_X1 U463 ( .A(G22GAT), .B(G141GAT), .Z(n400) );
  XNOR2_X1 U464 ( .A(G169GAT), .B(G113GAT), .ZN(n399) );
  XNOR2_X1 U465 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U466 ( .A(G36GAT), .B(G50GAT), .Z(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U468 ( .A(n404), .B(n403), .ZN(n405) );
  NOR2_X1 U469 ( .A1(n407), .A2(n571), .ZN(n408) );
  XNOR2_X1 U470 ( .A(KEYINPUT114), .B(n408), .ZN(n416) );
  INV_X1 U471 ( .A(KEYINPUT47), .ZN(n414) );
  XNOR2_X1 U472 ( .A(KEYINPUT110), .B(n480), .ZN(n560) );
  INV_X1 U473 ( .A(n571), .ZN(n557) );
  XNOR2_X1 U474 ( .A(n409), .B(KEYINPUT46), .ZN(n410) );
  NOR2_X1 U475 ( .A1(n560), .A2(n410), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n411), .B(KEYINPUT111), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n415) );
  NOR2_X1 U478 ( .A1(n416), .A2(n415), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n458) );
  XOR2_X1 U480 ( .A(n419), .B(n420), .Z(n422) );
  NAND2_X1 U481 ( .A1(G226GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n424) );
  XOR2_X1 U483 ( .A(n424), .B(n423), .Z(n431) );
  XOR2_X1 U484 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n426) );
  XNOR2_X1 U485 ( .A(KEYINPUT88), .B(KEYINPUT18), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U487 ( .A(G169GAT), .B(n427), .Z(n450) );
  INV_X1 U488 ( .A(n428), .ZN(n429) );
  XOR2_X1 U489 ( .A(n450), .B(n429), .Z(n430) );
  XOR2_X1 U490 ( .A(n431), .B(n430), .Z(n502) );
  INV_X1 U491 ( .A(n502), .ZN(n528) );
  NOR2_X1 U492 ( .A1(n458), .A2(n528), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n436), .B(KEYINPUT55), .ZN(n453) );
  XOR2_X1 U495 ( .A(G99GAT), .B(G190GAT), .Z(n438) );
  XNOR2_X1 U496 ( .A(G183GAT), .B(G71GAT), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U498 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U501 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n444) );
  XNOR2_X1 U502 ( .A(G43GAT), .B(G176GAT), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U504 ( .A(n446), .B(n445), .Z(n452) );
  XOR2_X1 U505 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n448) );
  XNOR2_X1 U506 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U509 ( .A(n452), .B(n451), .Z(n530) );
  INV_X1 U510 ( .A(n530), .ZN(n505) );
  NAND2_X1 U511 ( .A1(n453), .A2(n505), .ZN(n559) );
  NOR2_X1 U512 ( .A1(n512), .A2(n559), .ZN(n456) );
  XNOR2_X1 U513 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n454) );
  XNOR2_X1 U514 ( .A(KEYINPUT28), .B(KEYINPUT65), .ZN(n457) );
  XOR2_X1 U515 ( .A(n457), .B(n468), .Z(n533) );
  INV_X1 U516 ( .A(n533), .ZN(n508) );
  XNOR2_X1 U517 ( .A(n502), .B(KEYINPUT27), .ZN(n472) );
  INV_X1 U518 ( .A(n567), .ZN(n499) );
  NAND2_X1 U519 ( .A1(n472), .A2(n499), .ZN(n476) );
  NOR2_X1 U520 ( .A1(n458), .A2(n476), .ZN(n545) );
  NAND2_X1 U521 ( .A1(n542), .A2(n563), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n463) );
  XNOR2_X1 U523 ( .A(n465), .B(n464), .ZN(G1343GAT) );
  XOR2_X1 U524 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n486) );
  NOR2_X1 U525 ( .A1(n576), .A2(n557), .ZN(n497) );
  NAND2_X1 U526 ( .A1(n505), .A2(n502), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n468), .A2(n466), .ZN(n467) );
  XOR2_X1 U528 ( .A(KEYINPUT25), .B(n467), .Z(n474) );
  NOR2_X1 U529 ( .A1(n505), .A2(n468), .ZN(n470) );
  XNOR2_X1 U530 ( .A(KEYINPUT99), .B(KEYINPUT26), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U532 ( .A(KEYINPUT98), .B(n471), .Z(n568) );
  NAND2_X1 U533 ( .A1(n472), .A2(n568), .ZN(n473) );
  NAND2_X1 U534 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n567), .A2(n475), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n508), .A2(n476), .ZN(n477) );
  NAND2_X1 U537 ( .A1(n477), .A2(n530), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n479), .A2(n478), .ZN(n493) );
  NAND2_X1 U539 ( .A1(n481), .A2(n480), .ZN(n482) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(n482), .Z(n483) );
  AND2_X1 U541 ( .A1(n493), .A2(n483), .ZN(n513) );
  NAND2_X1 U542 ( .A1(n497), .A2(n513), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT100), .B(n484), .Z(n491) );
  NAND2_X1 U544 ( .A1(n491), .A2(n499), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NAND2_X1 U547 ( .A1(n491), .A2(n502), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U550 ( .A1(n505), .A2(n491), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NAND2_X1 U552 ( .A1(n491), .A2(n508), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .Z(n501) );
  NAND2_X1 U555 ( .A1(n291), .A2(n493), .ZN(n494) );
  NOR2_X1 U556 ( .A1(n480), .A2(n494), .ZN(n496) );
  XOR2_X1 U557 ( .A(KEYINPUT37), .B(KEYINPUT102), .Z(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n525) );
  NAND2_X1 U559 ( .A1(n525), .A2(n497), .ZN(n498) );
  XOR2_X1 U560 ( .A(KEYINPUT38), .B(n498), .Z(n509) );
  NAND2_X1 U561 ( .A1(n509), .A2(n499), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  XOR2_X1 U563 ( .A(G36GAT), .B(KEYINPUT103), .Z(n504) );
  NAND2_X1 U564 ( .A1(n509), .A2(n502), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n509), .A2(n505), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n506), .B(KEYINPUT40), .ZN(n507) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NAND2_X1 U569 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U570 ( .A(n510), .B(KEYINPUT104), .ZN(n511) );
  XNOR2_X1 U571 ( .A(G50GAT), .B(n511), .ZN(G1331GAT) );
  NOR2_X1 U572 ( .A1(n571), .A2(n512), .ZN(n526) );
  NAND2_X1 U573 ( .A1(n526), .A2(n513), .ZN(n514) );
  XOR2_X1 U574 ( .A(KEYINPUT105), .B(n514), .Z(n521) );
  NOR2_X1 U575 ( .A1(n567), .A2(n521), .ZN(n516) );
  XNOR2_X1 U576 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n515) );
  XNOR2_X1 U577 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n517), .Z(G1332GAT) );
  NOR2_X1 U579 ( .A1(n528), .A2(n521), .ZN(n519) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n519), .B(n518), .ZN(G1333GAT) );
  NOR2_X1 U582 ( .A1(n530), .A2(n521), .ZN(n520) );
  XOR2_X1 U583 ( .A(G71GAT), .B(n520), .Z(G1334GAT) );
  NOR2_X1 U584 ( .A1(n533), .A2(n521), .ZN(n523) );
  XNOR2_X1 U585 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G78GAT), .B(n524), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n532) );
  NOR2_X1 U589 ( .A1(n567), .A2(n532), .ZN(n527) );
  XOR2_X1 U590 ( .A(G85GAT), .B(n527), .Z(G1336GAT) );
  NOR2_X1 U591 ( .A1(n528), .A2(n532), .ZN(n529) );
  XOR2_X1 U592 ( .A(G92GAT), .B(n529), .Z(G1337GAT) );
  NOR2_X1 U593 ( .A1(n530), .A2(n532), .ZN(n531) );
  XOR2_X1 U594 ( .A(G99GAT), .B(n531), .Z(G1338GAT) );
  NOR2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n535) );
  XNOR2_X1 U596 ( .A(KEYINPUT109), .B(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  NAND2_X1 U599 ( .A1(n571), .A2(n542), .ZN(n537) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT118), .Z(n539) );
  NAND2_X1 U602 ( .A1(n551), .A2(n542), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U604 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U606 ( .A1(n542), .A2(n560), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n543), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  NAND2_X1 U609 ( .A1(n568), .A2(n545), .ZN(n546) );
  XOR2_X1 U610 ( .A(KEYINPUT120), .B(n546), .Z(n555) );
  NAND2_X1 U611 ( .A1(n571), .A2(n555), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n549) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U616 ( .A(KEYINPUT121), .B(n550), .Z(n553) );
  NAND2_X1 U617 ( .A1(n551), .A2(n555), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n555), .A2(n480), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n563), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n559), .ZN(n558) );
  XOR2_X1 U624 ( .A(G169GAT), .B(n558), .Z(G1348GAT) );
  NAND2_X1 U625 ( .A1(n562), .A2(n560), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n564), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(G190GAT), .ZN(G1351GAT) );
  AND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U632 ( .A(KEYINPUT125), .B(n570), .ZN(n581) );
  AND2_X1 U633 ( .A1(n571), .A2(n581), .ZN(n575) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(KEYINPUT60), .ZN(n573) );
  XNOR2_X1 U636 ( .A(KEYINPUT126), .B(n573), .ZN(n574) );
  XNOR2_X1 U637 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U639 ( .A1(n581), .A2(n576), .ZN(n577) );
  XNOR2_X1 U640 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n480), .A2(n581), .ZN(n579) );
  XNOR2_X1 U642 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U643 ( .A1(n581), .A2(n291), .ZN(n582) );
  XNOR2_X1 U644 ( .A(n582), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

