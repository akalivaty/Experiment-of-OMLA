//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1124,
    new_n1125, new_n1126, new_n1127;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT64), .Z(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n464), .B1(new_n463), .B2(new_n465), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n460), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n461), .ZN(new_n473));
  NAND3_X1  g048(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n475), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n476));
  OR2_X1    g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  XOR2_X1   g054(.A(new_n475), .B(KEYINPUT67), .Z(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(new_n483), .B2(G112), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n482), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  AND3_X1   g066(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT69), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n495), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n498));
  XOR2_X1   g073(.A(KEYINPUT70), .B(KEYINPUT4), .Z(new_n499));
  OAI211_X1 g074(.A(new_n491), .B(new_n499), .C1(new_n466), .C2(new_n467), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(new_n483), .B2(G114), .ZN(new_n502));
  INV_X1    g077(.A(G102), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(new_n483), .ZN(new_n504));
  OAI211_X1 g079(.A(G126), .B(G2105), .C1(new_n492), .C2(new_n493), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT68), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n475), .A2(new_n507), .A3(G126), .A4(G2105), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n501), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT71), .B1(new_n512), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT6), .B(G651), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n523), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n519), .A2(new_n523), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n522), .A2(new_n528), .ZN(G166));
  AND2_X1   g104(.A1(new_n519), .A2(new_n523), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n524), .A2(G51), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n531), .A2(new_n533), .A3(new_n534), .A4(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  AOI22_X1  g112(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n521), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n530), .A2(G90), .B1(G52), .B2(new_n524), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n521), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n524), .A2(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n526), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n524), .A2(G53), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(KEYINPUT72), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n555), .B(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G91), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OAI221_X1 g135(.A(new_n558), .B1(new_n559), .B2(new_n526), .C1(new_n521), .C2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND2_X1  g137(.A1(new_n530), .A2(G87), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n524), .A2(G49), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  AOI22_X1  g141(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  OR3_X1    g142(.A1(new_n567), .A2(KEYINPUT73), .A3(new_n521), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n530), .A2(G86), .B1(G48), .B2(new_n524), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT73), .B1(new_n567), .B2(new_n521), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G305));
  AOI22_X1  g146(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n530), .A2(G85), .B1(G47), .B2(new_n524), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(G301), .A2(G868), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n519), .A2(G66), .ZN(new_n578));
  NAND2_X1  g153(.A1(G79), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G54), .B2(new_n524), .ZN(new_n581));
  XOR2_X1   g156(.A(KEYINPUT75), .B(KEYINPUT10), .Z(new_n582));
  NAND3_X1  g157(.A1(new_n530), .A2(G92), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n582), .ZN(new_n584));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n526), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n581), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT76), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n577), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n577), .B1(new_n593), .B2(G868), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G299), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n481), .A2(G123), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n484), .A2(G135), .ZN(new_n607));
  NOR2_X1   g182(.A1(G99), .A2(G2105), .ZN(new_n608));
  OAI21_X1  g183(.A(G2104), .B1(new_n483), .B2(G111), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n606), .B(new_n607), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G2096), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n466), .A2(new_n467), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n462), .A2(G2105), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n615), .B(new_n616), .Z(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT13), .B(G2100), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n612), .A2(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2435), .ZN(new_n622));
  XOR2_X1   g197(.A(G2427), .B(G2438), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XOR2_X1   g200(.A(G2451), .B(G2454), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2443), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT78), .B(KEYINPUT79), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2446), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n631), .B(new_n633), .Z(new_n634));
  AND2_X1   g209(.A1(new_n634), .A2(G14), .ZN(G401));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT80), .ZN(new_n637));
  XOR2_X1   g212(.A(G2084), .B(G2090), .Z(new_n638));
  XNOR2_X1  g213(.A(G2072), .B(G2078), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n637), .B(KEYINPUT82), .ZN(new_n643));
  INV_X1    g218(.A(new_n638), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT17), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(new_n639), .Z(new_n647));
  NOR2_X1   g222(.A1(new_n643), .A2(new_n644), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n642), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(new_n611), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(G227));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1961), .B(G1966), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT83), .ZN(new_n654));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n652), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n654), .A2(new_n655), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n661), .A2(new_n658), .A3(new_n656), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n656), .A2(new_n652), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n663), .A2(new_n660), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n659), .B(new_n662), .C1(new_n664), .C2(new_n658), .ZN(new_n665));
  XOR2_X1   g240(.A(G1991), .B(G1996), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G229));
  NOR2_X1   g246(.A1(G5), .A2(G16), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(G171), .B2(G16), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G1961), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT97), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT31), .B(G11), .ZN(new_n676));
  OR2_X1    g251(.A1(G16), .A2(G21), .ZN(new_n677));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(G286), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(G1966), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT96), .ZN(new_n682));
  INV_X1    g257(.A(G29), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n610), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  INV_X1    g260(.A(G28), .ZN(new_n686));
  AOI21_X1  g261(.A(G29), .B1(new_n686), .B2(KEYINPUT30), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(KEYINPUT30), .B2(new_n686), .ZN(new_n688));
  AND3_X1   g263(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n675), .A2(new_n676), .A3(new_n682), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT98), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT99), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n678), .A2(G20), .ZN(new_n693));
  OAI211_X1 g268(.A(KEYINPUT23), .B(new_n693), .C1(new_n597), .C2(new_n678), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(KEYINPUT23), .B2(new_n693), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G1956), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(G1956), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n683), .A2(G35), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G162), .B2(new_n683), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT29), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n696), .A2(new_n697), .B1(G2090), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n691), .B1(new_n692), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n548), .A2(new_n678), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n678), .B2(G19), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(G1341), .ZN(new_n706));
  NOR2_X1   g281(.A1(G29), .A2(G32), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n481), .A2(G129), .B1(G105), .B2(new_n614), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT26), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n484), .A2(G141), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n707), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT27), .B(G1996), .Z(new_n715));
  AOI22_X1  g290(.A1(new_n714), .A2(new_n715), .B1(new_n705), .B2(G1341), .ZN(new_n716));
  OAI221_X1 g291(.A(new_n716), .B1(new_n714), .B2(new_n715), .C1(new_n700), .C2(G2090), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n484), .A2(G139), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n614), .A2(G103), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  AOI22_X1  g295(.A1(new_n613), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n718), .B(new_n720), .C1(new_n483), .C2(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G33), .B(new_n722), .S(G29), .Z(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G2072), .Z(new_n724));
  NOR2_X1   g299(.A1(KEYINPUT24), .A2(G34), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  AOI21_X1  g302(.A(G29), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI22_X1  g303(.A1(G160), .A2(G29), .B1(KEYINPUT95), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(KEYINPUT95), .B2(new_n728), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2084), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n673), .A2(G1961), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n683), .A2(G27), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G164), .B2(new_n683), .ZN(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n724), .A2(new_n731), .A3(new_n732), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n678), .A2(G4), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n593), .B2(new_n678), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1348), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n717), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n701), .A2(new_n692), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n702), .A2(new_n706), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n678), .A2(G23), .ZN(new_n744));
  INV_X1    g319(.A(G288), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n678), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT88), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT33), .B(G1976), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  MUX2_X1   g324(.A(G6), .B(G305), .S(G16), .Z(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT32), .B(G1981), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n678), .A2(G22), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G166), .B2(new_n678), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1971), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n749), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT34), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n678), .A2(G24), .ZN(new_n765));
  INV_X1    g340(.A(G290), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(new_n678), .ZN(new_n767));
  INV_X1    g342(.A(G1986), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT84), .ZN(new_n770));
  INV_X1    g345(.A(G25), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G29), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(G29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n481), .A2(G119), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT85), .ZN(new_n775));
  OR2_X1    g350(.A1(G95), .A2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n776), .B(G2104), .C1(G107), .C2(new_n483), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n484), .A2(G131), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n773), .B1(new_n779), .B2(G29), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n772), .B1(new_n780), .B2(new_n770), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(KEYINPUT87), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT35), .B(G1991), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT86), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT87), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(new_n772), .C1(new_n780), .C2(new_n770), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n782), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n785), .B1(new_n782), .B2(new_n787), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n788), .A2(new_n789), .A3(KEYINPUT90), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n760), .A2(KEYINPUT34), .A3(new_n761), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n764), .A2(new_n769), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n743), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n791), .A2(new_n790), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n795), .A2(KEYINPUT36), .A3(new_n769), .A4(new_n764), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n683), .A2(G26), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT93), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT28), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n484), .A2(G140), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT91), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n484), .A2(KEYINPUT91), .A3(G140), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(G104), .A2(G2105), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n805), .B(G2104), .C1(G116), .C2(new_n483), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n481), .A2(G128), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G29), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n809), .A2(KEYINPUT92), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(KEYINPUT92), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n799), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT94), .B(G2067), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  AND3_X1   g389(.A1(new_n794), .A2(new_n796), .A3(new_n814), .ZN(G311));
  NAND3_X1  g390(.A1(new_n794), .A2(new_n814), .A3(new_n796), .ZN(G150));
  AOI22_X1  g391(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(new_n521), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n524), .A2(G55), .ZN(new_n819));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n526), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NOR2_X1   g400(.A1(new_n592), .A2(new_n600), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT39), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n548), .B(new_n822), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(G860), .ZN(G145));
  XNOR2_X1  g407(.A(new_n610), .B(G160), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G162), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n712), .B(new_n510), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(new_n617), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n617), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n779), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n837), .A2(new_n779), .A3(new_n838), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n722), .A2(KEYINPUT101), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n808), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n808), .A2(new_n842), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n481), .A2(G130), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n484), .A2(G142), .ZN(new_n846));
  OR2_X1    g421(.A1(G106), .A2(G2105), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n847), .B(G2104), .C1(G118), .C2(new_n483), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n843), .A2(new_n844), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n843), .A2(new_n844), .ZN(new_n851));
  INV_X1    g426(.A(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n840), .A2(new_n841), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n841), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n850), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n855), .A2(new_n856), .A3(new_n839), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n835), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n840), .A2(new_n850), .A3(new_n853), .A4(new_n841), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n856), .B1(new_n855), .B2(new_n839), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n861), .A3(new_n834), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT102), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n858), .A2(new_n865), .A3(new_n859), .A4(new_n862), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n864), .A2(KEYINPUT40), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT40), .B1(new_n864), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(G395));
  INV_X1    g444(.A(G868), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n823), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n602), .B(new_n830), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n597), .A2(new_n587), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n588), .A2(G299), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(KEYINPUT41), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n873), .B2(new_n874), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n876), .B1(new_n872), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT42), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n766), .A2(G288), .ZN(new_n884));
  XNOR2_X1  g459(.A(G305), .B(G303), .ZN(new_n885));
  NOR2_X1   g460(.A1(G290), .A2(new_n745), .ZN(new_n886));
  OR4_X1    g461(.A1(new_n883), .A2(new_n884), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G290), .B(G288), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT103), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n885), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n882), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n871), .B1(new_n893), .B2(new_n870), .ZN(G295));
  OAI21_X1  g469(.A(new_n871), .B1(new_n893), .B2(new_n870), .ZN(G331));
  XNOR2_X1  g470(.A(G301), .B(G286), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n830), .A3(KEYINPUT104), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n896), .A2(new_n830), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n830), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n880), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n900), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n903), .A2(new_n875), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n892), .A2(KEYINPUT105), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n902), .A2(new_n904), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(KEYINPUT105), .A3(new_n892), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n859), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n880), .A2(new_n903), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT106), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n880), .A2(new_n915), .A3(new_n903), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n875), .B1(new_n901), .B2(new_n897), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n892), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n908), .A2(new_n892), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n919), .A2(KEYINPUT43), .A3(new_n859), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n912), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT44), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n919), .A2(new_n911), .A3(new_n859), .A4(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n923), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n927), .B1(new_n912), .B2(new_n921), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT44), .B1(new_n924), .B2(new_n925), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT107), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(G397));
  INV_X1    g509(.A(G2067), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n808), .B(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n471), .A2(G40), .A3(new_n477), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G1384), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n510), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OR3_X1    g517(.A1(new_n938), .A2(new_n942), .A3(KEYINPUT108), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT108), .B1(new_n938), .B2(new_n942), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n936), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT109), .ZN(new_n948));
  INV_X1    g523(.A(G1996), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n712), .B(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n779), .B(new_n784), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n945), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(G290), .B(G1986), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n945), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT123), .ZN(new_n958));
  INV_X1    g533(.A(G8), .ZN(new_n959));
  AOI211_X1 g534(.A(new_n941), .B(G1384), .C1(new_n501), .C2(new_n509), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT45), .B1(new_n510), .B2(new_n939), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n942), .A2(KEYINPUT110), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n937), .ZN(new_n965));
  INV_X1    g540(.A(G1971), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT50), .B1(new_n510), .B2(new_n939), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  AOI211_X1 g544(.A(new_n969), .B(G1384), .C1(new_n501), .C2(new_n509), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n937), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n971), .A2(G2090), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n959), .B1(new_n973), .B2(KEYINPUT114), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(KEYINPUT114), .B2(new_n973), .ZN(new_n975));
  NAND2_X1  g550(.A1(G303), .A2(G8), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT55), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(KEYINPUT115), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n569), .B1(new_n521), .B2(new_n567), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(G1981), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(G305), .B2(G1981), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT112), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n982), .A2(KEYINPUT49), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n501), .B2(new_n509), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n937), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G8), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(KEYINPUT49), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n983), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n986), .B1(G1976), .B2(new_n745), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT111), .B(G1976), .Z(new_n993));
  OAI211_X1 g568(.A(new_n990), .B(new_n991), .C1(new_n745), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n989), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n978), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n959), .B1(new_n967), .B2(new_n972), .ZN(new_n998));
  INV_X1    g573(.A(new_n977), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n975), .A2(new_n977), .B1(KEYINPUT115), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n958), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n975), .A2(new_n977), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(KEYINPUT115), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1005), .A2(KEYINPUT123), .A3(new_n996), .A4(new_n978), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT121), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n942), .A2(new_n937), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n680), .ZN(new_n1012));
  INV_X1    g587(.A(G2084), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1013), .B(new_n937), .C1(new_n968), .C2(new_n970), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n959), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1009), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n961), .A2(new_n960), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1966), .B1(new_n1018), .B2(new_n937), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1014), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1016), .B(G8), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G286), .A2(G8), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT119), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1008), .B1(new_n1017), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(G8), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT51), .B1(new_n1027), .B2(KEYINPUT120), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1023), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(KEYINPUT121), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT51), .B1(new_n1015), .B2(new_n1023), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT62), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1023), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(KEYINPUT122), .A2(KEYINPUT53), .ZN(new_n1036));
  OR2_X1    g611(.A1(KEYINPUT122), .A2(KEYINPUT53), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1036), .B(new_n1037), .C1(new_n965), .C2(G2078), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n735), .A2(KEYINPUT53), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n971), .A2(KEYINPUT117), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(new_n937), .C1(new_n968), .C2(new_n970), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  OAI221_X1 g618(.A(new_n1038), .B1(new_n1011), .B2(new_n1039), .C1(new_n1043), .C2(G1961), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1044), .A2(G171), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1035), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT125), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(KEYINPUT62), .ZN(new_n1049));
  AOI211_X1 g624(.A(KEYINPUT125), .B(new_n1033), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1348), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n985), .A2(G2067), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(new_n592), .ZN(new_n1055));
  XNOR2_X1  g630(.A(G299), .B(KEYINPUT57), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT56), .B(G2072), .Z(new_n1057));
  INV_X1    g632(.A(new_n971), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n965), .A2(new_n1057), .B1(new_n1058), .B2(G1956), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1055), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1056), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1059), .A2(new_n1056), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(KEYINPUT61), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1054), .A2(new_n1064), .A3(new_n593), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1052), .A2(new_n593), .A3(new_n1053), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT60), .B1(new_n1055), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n1069));
  INV_X1    g644(.A(new_n985), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT58), .B(G1341), .ZN(new_n1071));
  OAI22_X1  g646(.A1(new_n965), .A2(G1996), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n548), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1073), .B1(new_n1072), .B2(new_n548), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1069), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1076), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(KEYINPUT59), .A3(new_n1074), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1060), .B(new_n1061), .C1(new_n1068), .C2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT54), .B1(G301), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(KEYINPUT54), .B2(G301), .ZN(new_n1084));
  XOR2_X1   g659(.A(new_n1044), .B(new_n1084), .Z(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(new_n1048), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1007), .B1(new_n1051), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1976), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n989), .A2(new_n1088), .A3(new_n745), .ZN(new_n1089));
  OR2_X1    g664(.A1(G305), .A2(G1981), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n986), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n995), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n989), .A2(KEYINPUT113), .A3(new_n992), .A4(new_n994), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n977), .A2(KEYINPUT116), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n998), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1015), .A2(G168), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n998), .B2(new_n1095), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1091), .B1(new_n1099), .B2(KEYINPUT63), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1097), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1005), .A2(new_n996), .A3(new_n1102), .A4(new_n978), .ZN(new_n1103));
  OAI221_X1 g678(.A(new_n1100), .B1(new_n1101), .B2(new_n1000), .C1(KEYINPUT63), .C2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n957), .B1(new_n1087), .B2(new_n1104), .ZN(new_n1105));
  NOR4_X1   g680(.A1(new_n948), .A2(new_n784), .A3(new_n779), .A4(new_n951), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n808), .A2(G2067), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n945), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n945), .A2(new_n768), .A3(new_n766), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT48), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n952), .A2(new_n954), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT46), .B1(new_n945), .B2(new_n949), .ZN(new_n1112));
  XOR2_X1   g687(.A(new_n1112), .B(KEYINPUT126), .Z(new_n1113));
  NAND3_X1  g688(.A1(new_n945), .A2(KEYINPUT46), .A3(new_n949), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1114), .B(KEYINPUT127), .Z(new_n1115));
  AND2_X1   g690(.A1(new_n936), .A2(new_n713), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1113), .B(new_n1115), .C1(new_n946), .C2(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1117), .A2(KEYINPUT47), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(KEYINPUT47), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1108), .B(new_n1111), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1105), .A2(new_n1121), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g697(.A(G319), .ZN(new_n1124));
  AOI211_X1 g698(.A(new_n1124), .B(G229), .C1(new_n924), .C2(new_n925), .ZN(new_n1125));
  NAND2_X1  g699(.A1(new_n864), .A2(new_n866), .ZN(new_n1126));
  NOR2_X1   g700(.A1(G227), .A2(G401), .ZN(new_n1127));
  AND3_X1   g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(G308));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(G225));
endmodule


