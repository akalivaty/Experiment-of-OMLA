//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n834, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G141gat), .B(G148gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n202), .B(new_n205), .C1(new_n206), .C2(KEYINPUT2), .ZN(new_n207));
  AND2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT75), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT75), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n205), .A2(new_n211), .A3(new_n202), .ZN(new_n212));
  AND2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n202), .A2(KEYINPUT76), .A3(KEYINPUT2), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT76), .B1(new_n202), .B2(KEYINPUT2), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n207), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT77), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n207), .B(new_n224), .C1(new_n216), .C2(new_n219), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n226));
  INV_X1    g025(.A(G113gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G120gat), .ZN(new_n228));
  INV_X1    g027(.A(G120gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G113gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n227), .A2(G120gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT67), .B1(new_n227), .B2(G120gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n237), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n232), .A2(new_n226), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n234), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n225), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n220), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n223), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT78), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT78), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n223), .A2(new_n242), .A3(new_n246), .A4(new_n243), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT4), .B1(new_n241), .B2(new_n220), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n250), .A2(KEYINPUT79), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n241), .A2(new_n220), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(KEYINPUT79), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n248), .A2(new_n249), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n249), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n241), .A2(new_n220), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(new_n252), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT5), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n260), .B2(KEYINPUT5), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT81), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n254), .A2(new_n250), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n269));
  AND4_X1   g068(.A1(new_n266), .A2(new_n248), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n267), .B1(new_n245), .B2(new_n247), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n266), .B1(new_n271), .B2(new_n269), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n265), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G1gat), .B(G29gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT0), .ZN(new_n275));
  XNOR2_X1  g074(.A(G57gat), .B(G85gat), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n275), .B(new_n276), .Z(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n277), .B(new_n265), .C1(new_n270), .C2(new_n272), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n273), .A2(KEYINPUT6), .A3(new_n278), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G8gat), .B(G36gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G226gat), .ZN(new_n289));
  INV_X1    g088(.A(G233gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G169gat), .ZN(new_n298));
  INV_X1    g097(.A(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(KEYINPUT26), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n293), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT27), .B(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n303), .A2(KEYINPUT28), .A3(new_n304), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n299), .A2(KEYINPUT64), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G176gat), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT23), .A4(new_n298), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n296), .A2(KEYINPUT23), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n300), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n317), .A2(new_n293), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT24), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n293), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n314), .B(new_n316), .C1(new_n318), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT65), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n293), .A2(new_n322), .A3(new_n319), .ZN(new_n323));
  OAI211_X1 g122(.A(G183gat), .B(G190gat), .C1(KEYINPUT65), .C2(KEYINPUT24), .ZN(new_n324));
  OR2_X1    g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n310), .B1(new_n294), .B2(KEYINPUT23), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n316), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT66), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n310), .A2(new_n321), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n326), .A2(KEYINPUT66), .A3(new_n316), .A4(new_n327), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n309), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n292), .B1(new_n332), .B2(KEYINPUT29), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n332), .B2(new_n292), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT22), .ZN(new_n336));
  XOR2_X1   g135(.A(KEYINPUT72), .B(G211gat), .Z(new_n337));
  INV_X1    g136(.A(G218gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G197gat), .B(G204gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G211gat), .B(G218gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n309), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n321), .A2(new_n310), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n329), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n331), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT73), .A3(new_n291), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n333), .A2(new_n335), .A3(new_n346), .A4(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n346), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n291), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n332), .A2(new_n292), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n288), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n353), .A2(new_n358), .A3(new_n288), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(KEYINPUT30), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n353), .A2(new_n358), .A3(new_n288), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n362), .A2(KEYINPUT74), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT74), .B1(new_n362), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT89), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT89), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n361), .B(new_n368), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n284), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT92), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT92), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n284), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G78gat), .B(G106gat), .ZN(new_n375));
  INV_X1    g174(.A(G50gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(KEYINPUT83), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n377), .B(new_n379), .Z(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n225), .A2(new_n355), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n354), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n345), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n342), .B1(new_n339), .B2(new_n340), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n355), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n346), .A2(KEYINPUT84), .A3(new_n355), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT3), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n220), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n383), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n346), .A2(new_n355), .A3(new_n220), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n220), .B2(KEYINPUT3), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT85), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n397), .B1(new_n398), .B2(new_n354), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n382), .A2(KEYINPUT85), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n225), .B2(new_n355), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n397), .B(new_n354), .C1(new_n400), .C2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n395), .B(new_n396), .C1(new_n399), .C2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT87), .B(G22gat), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n394), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n394), .B2(new_n405), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n381), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n405), .A3(new_n406), .ZN(new_n410));
  INV_X1    g209(.A(G22gat), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n411), .B1(new_n394), .B2(new_n405), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT88), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n410), .B(new_n380), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n405), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n413), .A3(G22gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n409), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n241), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n351), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n332), .A2(new_n241), .ZN(new_n421));
  NAND2_X1  g220(.A1(G227gat), .A2(G233gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT68), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(KEYINPUT68), .A3(new_n425), .ZN(new_n429));
  XNOR2_X1  g228(.A(G15gat), .B(G43gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT69), .ZN(new_n431));
  XNOR2_X1  g230(.A(G71gat), .B(G99gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n424), .B2(KEYINPUT32), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n433), .B(KEYINPUT70), .Z(new_n436));
  OAI211_X1 g235(.A(KEYINPUT32), .B(new_n424), .C1(new_n436), .C2(new_n425), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n423), .B1(new_n420), .B2(new_n421), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT34), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n439), .A2(KEYINPUT71), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n421), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(new_n440), .A3(new_n422), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT71), .B1(new_n439), .B2(new_n440), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n438), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n435), .A2(new_n445), .A3(new_n437), .A4(new_n446), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT35), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n418), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n372), .A2(new_n374), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n366), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n284), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n418), .A2(new_n451), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT35), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n353), .A2(new_n358), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n333), .A2(new_n335), .A3(new_n354), .A4(new_n352), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n346), .B1(new_n356), .B2(new_n357), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT37), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT38), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n461), .A2(new_n464), .A3(new_n465), .A4(new_n287), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n362), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n353), .A2(new_n358), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT37), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n287), .A3(new_n461), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n467), .B1(new_n470), .B2(KEYINPUT38), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n282), .A3(new_n283), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT39), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n248), .A2(new_n268), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n474), .B1(new_n475), .B2(new_n258), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n271), .A2(KEYINPUT90), .A3(new_n249), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n474), .A3(new_n258), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT90), .B1(new_n271), .B2(new_n249), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n259), .A2(new_n252), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n473), .B1(new_n481), .B2(new_n249), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n478), .A2(KEYINPUT40), .A3(new_n277), .A4(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n478), .A2(new_n277), .A3(new_n483), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT40), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n489), .A2(new_n367), .A3(new_n279), .A4(new_n369), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n418), .B(new_n472), .C1(new_n486), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n450), .A2(KEYINPUT36), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n448), .A2(new_n493), .A3(new_n449), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n418), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(new_n457), .B2(new_n496), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n455), .A2(new_n459), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G15gat), .B(G22gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT16), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(G1gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(KEYINPUT96), .A2(G8gat), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n501), .B(new_n502), .C1(G1gat), .C2(new_n499), .ZN(new_n503));
  NOR2_X1   g302(.A1(KEYINPUT96), .A2(G8gat), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n504), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT97), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT97), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n505), .A2(new_n509), .A3(new_n506), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(G57gat), .A2(G64gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(G57gat), .A2(G64gat), .ZN(new_n513));
  AND2_X1   g312(.A1(G71gat), .A2(G78gat), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(KEYINPUT9), .ZN(new_n515));
  NOR2_X1   g314(.A1(G71gat), .A2(G78gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n515), .A2(new_n517), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT99), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT99), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n515), .A2(new_n521), .A3(new_n517), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n518), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n511), .A2(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n527));
  NOR2_X1   g326(.A1(new_n524), .A2(KEYINPUT21), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT100), .ZN(new_n529));
  AND2_X1   g328(.A1(G231gat), .A2(G233gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n530), .ZN(new_n533));
  XNOR2_X1  g332(.A(G127gat), .B(G155gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n534), .B1(new_n532), .B2(new_n533), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n527), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  INV_X1    g338(.A(new_n527), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n526), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n538), .A2(new_n541), .A3(new_n526), .ZN(new_n544));
  XOR2_X1   g343(.A(G183gat), .B(G211gat), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n544), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n545), .B1(new_n548), .B2(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OR3_X1    g350(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT93), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT93), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G29gat), .ZN(new_n558));
  INV_X1    g357(.A(G36gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n376), .A2(G43gat), .ZN(new_n562));
  INV_X1    g361(.A(G43gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G50gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n562), .A2(new_n564), .A3(KEYINPUT15), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT95), .B1(new_n376), .B2(G43gat), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n563), .B2(G50gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n376), .A2(KEYINPUT95), .A3(G43gat), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT15), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n565), .A2(KEYINPUT94), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(KEYINPUT94), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n560), .B1(new_n552), .B2(new_n555), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI22_X1  g372(.A1(new_n561), .A2(new_n565), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT17), .ZN(new_n575));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  INV_X1    g375(.A(G85gat), .ZN(new_n577));
  INV_X1    g376(.A(G92gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(KEYINPUT8), .A2(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT7), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n577), .B2(new_n578), .ZN(new_n581));
  NAND3_X1  g380(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G99gat), .B(G106gat), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n583), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n575), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n574), .B2(new_n586), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT101), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT102), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n591), .A2(new_n593), .ZN(new_n597));
  OR3_X1    g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  OAI21_X1  g400(.A(new_n596), .B1(new_n595), .B2(new_n597), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n601), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n596), .B(new_n604), .C1(new_n595), .C2(new_n597), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G113gat), .B(G141gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT11), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n298), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G197gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT13), .Z(new_n614));
  AOI21_X1  g413(.A(new_n574), .B1(new_n508), .B2(new_n510), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n508), .A2(new_n510), .A3(new_n574), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n616), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n614), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n575), .A2(new_n507), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(new_n613), .A3(new_n617), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n622), .A2(KEYINPUT18), .A3(new_n613), .A4(new_n617), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n612), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n621), .A2(new_n625), .A3(new_n627), .A4(new_n612), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n524), .B(new_n586), .C1(KEYINPUT103), .C2(new_n585), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT10), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n585), .A2(KEYINPUT103), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n587), .B1(new_n523), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n524), .A2(KEYINPUT10), .A3(new_n586), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n633), .A2(new_n636), .ZN(new_n642));
  INV_X1    g441(.A(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(G120gat), .B(G148gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT104), .ZN(new_n646));
  XOR2_X1   g445(.A(G176gat), .B(G204gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n641), .A2(new_n644), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n641), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n639), .A2(KEYINPUT106), .A3(new_n640), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n644), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n648), .B(KEYINPUT105), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n651), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n632), .A2(new_n658), .ZN(new_n659));
  NOR4_X1   g458(.A1(new_n498), .A2(new_n551), .A3(new_n607), .A4(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n284), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT107), .B(G1gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1324gat));
  INV_X1    g463(.A(new_n370), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  NAND3_X1  g465(.A1(new_n660), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  OR3_X1    g467(.A1(new_n667), .A2(KEYINPUT108), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT108), .B1(new_n667), .B2(new_n668), .ZN(new_n670));
  INV_X1    g469(.A(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n660), .A2(new_n665), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n668), .B1(new_n672), .B2(G8gat), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n669), .B(new_n670), .C1(new_n671), .C2(new_n673), .ZN(G1325gat));
  INV_X1    g473(.A(G15gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n675), .A3(new_n451), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n660), .A2(new_n495), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(new_n675), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n496), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  NOR2_X1   g480(.A1(new_n498), .A2(new_n606), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n550), .A2(new_n659), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n661), .A2(new_n558), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT109), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n687), .A2(KEYINPUT45), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n498), .B2(new_n606), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n415), .A2(G22gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT88), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n692), .A2(new_n410), .A3(new_n380), .A4(new_n416), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n450), .B1(new_n693), .B2(new_n409), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n366), .B1(new_n282), .B2(new_n283), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n452), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n283), .A2(new_n282), .B1(new_n367), .B2(new_n369), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n453), .B1(new_n373), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n698), .B2(new_n372), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n448), .A2(new_n493), .A3(new_n449), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n493), .B1(new_n448), .B2(new_n449), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n695), .B2(new_n418), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n484), .B(KEYINPUT91), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n704), .A2(new_n279), .A3(new_n665), .A4(new_n489), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n472), .A2(new_n418), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI211_X1 g506(.A(KEYINPUT44), .B(new_n607), .C1(new_n699), .C2(new_n707), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n690), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n683), .ZN(new_n710));
  OAI21_X1  g509(.A(G29gat), .B1(new_n710), .B2(new_n284), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n687), .A2(KEYINPUT45), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n688), .A2(new_n711), .A3(new_n712), .ZN(G1328gat));
  NAND4_X1  g512(.A1(new_n682), .A2(new_n559), .A3(new_n665), .A4(new_n683), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT46), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT110), .ZN(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n710), .B2(new_n370), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n716), .B(new_n717), .C1(KEYINPUT46), .C2(new_n714), .ZN(G1329gat));
  NAND4_X1  g517(.A1(new_n690), .A2(new_n495), .A3(new_n683), .A4(new_n708), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G43gat), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n450), .A2(G43gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n682), .A2(new_n683), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(new_n722), .A3(KEYINPUT47), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n724));
  INV_X1    g523(.A(new_n722), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n720), .B2(KEYINPUT111), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n719), .A2(new_n727), .A3(G43gat), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n724), .B(KEYINPUT47), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n720), .A2(KEYINPUT111), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n728), .A3(new_n722), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT112), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n723), .B1(new_n729), .B2(new_n733), .ZN(G1330gat));
  OAI21_X1  g533(.A(new_n376), .B1(new_n684), .B2(new_n418), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n496), .A2(G50gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n710), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g537(.A1(new_n550), .A2(new_n606), .A3(new_n631), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n739), .A2(new_n498), .A3(new_n658), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n661), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n665), .ZN(new_n743));
  NOR2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  AND2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n744), .B2(new_n743), .ZN(G1333gat));
  NAND2_X1  g546(.A1(new_n740), .A2(new_n495), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n450), .A2(G71gat), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n748), .A2(G71gat), .B1(new_n740), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n740), .A2(new_n496), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT113), .B(G78gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n550), .A2(new_n632), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n682), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n658), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n758), .A2(new_n577), .A3(new_n661), .A4(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n550), .A2(new_n632), .A3(new_n658), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n709), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G85gat), .B1(new_n762), .B2(new_n284), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(G1336gat));
  NOR3_X1   g563(.A1(new_n370), .A2(new_n658), .A3(G92gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n758), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n690), .A2(new_n665), .A3(new_n708), .A4(new_n761), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n756), .A2(KEYINPUT114), .A3(new_n757), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n757), .A2(KEYINPUT114), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n682), .A2(new_n755), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT115), .B1(new_n774), .B2(new_n765), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776));
  INV_X1    g575(.A(new_n765), .ZN(new_n777));
  AOI211_X1 g576(.A(new_n776), .B(new_n777), .C1(new_n771), .C2(new_n773), .ZN(new_n778));
  INV_X1    g577(.A(new_n769), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n775), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n770), .B1(new_n780), .B2(new_n767), .ZN(G1337gat));
  NOR3_X1   g580(.A1(new_n658), .A2(G99gat), .A3(new_n450), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n758), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G99gat), .B1(new_n762), .B2(new_n702), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1338gat));
  NAND3_X1  g584(.A1(new_n709), .A2(new_n496), .A3(new_n761), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n418), .A2(new_n658), .A3(G106gat), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n774), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n758), .A2(new_n788), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n790), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n789), .A2(new_n790), .B1(new_n792), .B2(new_n787), .ZN(G1339gat));
  NAND4_X1  g592(.A1(new_n550), .A2(new_n606), .A3(new_n631), .A4(new_n658), .ZN(new_n794));
  XNOR2_X1  g593(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n653), .A2(new_n654), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n639), .B2(new_n640), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n637), .A2(new_n643), .A3(new_n638), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n649), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n796), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n650), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT55), .B1(new_n796), .B2(new_n800), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT117), .B1(new_n802), .B2(new_n805), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n632), .A3(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n618), .A2(new_n620), .A3(new_n614), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n613), .B1(new_n622), .B2(new_n617), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n611), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n629), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n658), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n607), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n813), .B(new_n817), .ZN(new_n818));
  AND4_X1   g617(.A1(new_n607), .A2(new_n818), .A3(new_n807), .A4(new_n808), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n794), .B1(new_n820), .B2(new_n550), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n665), .A2(new_n284), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n694), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n632), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g625(.A1(new_n759), .A2(new_n229), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT120), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n759), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n830), .A2(KEYINPUT119), .A3(G120gat), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT119), .B1(new_n830), .B2(G120gat), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(G1341gat));
  NAND2_X1  g632(.A1(new_n824), .A2(new_n550), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(G127gat), .ZN(G1342gat));
  AOI21_X1  g634(.A(new_n606), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n823), .A2(new_n694), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n837), .B(new_n838), .Z(G1343gat));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n495), .A2(new_n665), .A3(new_n284), .ZN(new_n841));
  INV_X1    g640(.A(G141gat), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n631), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n821), .B2(new_n496), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n496), .A2(KEYINPUT57), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n814), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n796), .A2(new_n800), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n796), .A2(KEYINPUT122), .A3(new_n800), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n632), .B(new_n803), .C1(new_n852), .C2(KEYINPUT55), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n607), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n551), .B1(new_n854), .B2(new_n819), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n845), .B1(new_n855), .B2(new_n794), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n841), .B(new_n843), .C1(new_n844), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n495), .A2(new_n418), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n821), .A2(new_n632), .A3(new_n822), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n842), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n840), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT123), .B(KEYINPUT58), .C1(new_n857), .C2(new_n860), .ZN(new_n864));
  OAI22_X1  g663(.A1(new_n863), .A2(new_n864), .B1(new_n862), .B2(new_n861), .ZN(G1344gat));
  AND2_X1   g664(.A1(new_n823), .A2(new_n858), .ZN(new_n866));
  INV_X1    g665(.A(G148gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n759), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n841), .B1(new_n844), .B2(new_n856), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n658), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(KEYINPUT59), .A3(new_n867), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n821), .A2(new_n496), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n418), .A2(KEYINPUT57), .ZN(new_n875));
  INV_X1    g674(.A(new_n854), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n607), .A2(new_n818), .A3(new_n803), .A4(new_n806), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n550), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n794), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n875), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n874), .A2(new_n759), .A3(new_n880), .A4(new_n841), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n872), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n868), .B1(new_n871), .B2(new_n882), .ZN(G1345gat));
  OAI21_X1  g682(.A(G155gat), .B1(new_n869), .B2(new_n551), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n203), .A3(new_n550), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1346gat));
  OAI21_X1  g685(.A(G162gat), .B1(new_n869), .B2(new_n606), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n823), .A2(new_n204), .A3(new_n607), .A4(new_n858), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(KEYINPUT124), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n661), .A2(new_n370), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n821), .A2(new_n694), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(G169gat), .B1(new_n895), .B2(new_n632), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n894), .B(KEYINPUT125), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n458), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n821), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n631), .A2(new_n298), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(G1348gat));
  AOI21_X1  g700(.A(G176gat), .B1(new_n895), .B2(new_n759), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n658), .B1(new_n311), .B2(new_n313), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n899), .B2(new_n903), .ZN(G1349gat));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n550), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G183gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n895), .A2(new_n303), .A3(new_n550), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(KEYINPUT126), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n908), .B(new_n910), .ZN(G1350gat));
  AOI21_X1  g710(.A(new_n304), .B1(new_n899), .B2(new_n607), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT61), .Z(new_n913));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n304), .A3(new_n607), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1351gat));
  AND2_X1   g714(.A1(new_n821), .A2(new_n894), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n858), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n631), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n897), .A2(new_n495), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n874), .A2(new_n880), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n632), .A2(G197gat), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n918), .A2(G197gat), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(G1352gat));
  NAND3_X1  g722(.A1(new_n874), .A2(new_n759), .A3(new_n880), .ZN(new_n924));
  INV_X1    g723(.A(new_n919), .ZN(new_n925));
  OAI21_X1  g724(.A(G204gat), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n658), .A2(G204gat), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n927), .B1(new_n917), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n916), .A2(KEYINPUT127), .A3(new_n858), .A4(new_n928), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n930), .A2(KEYINPUT62), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT62), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n926), .B1(new_n932), .B2(new_n933), .ZN(G1353gat));
  INV_X1    g733(.A(new_n917), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n337), .A3(new_n550), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n874), .A2(new_n550), .A3(new_n880), .A4(new_n919), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT63), .B1(new_n937), .B2(G211gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(G1354gat));
  OAI21_X1  g740(.A(G218gat), .B1(new_n920), .B2(new_n606), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n935), .A2(new_n338), .A3(new_n607), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1355gat));
endmodule


