

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U551 ( .A(KEYINPUT30), .ZN(n722) );
  XNOR2_X1 U552 ( .A(n722), .B(KEYINPUT103), .ZN(n723) );
  XNOR2_X1 U553 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U554 ( .A(KEYINPUT32), .B(KEYINPUT104), .ZN(n739) );
  XNOR2_X1 U555 ( .A(n740), .B(n739), .ZN(n760) );
  NAND2_X1 U556 ( .A1(n688), .A2(n687), .ZN(n732) );
  XNOR2_X1 U557 ( .A(KEYINPUT68), .B(n517), .ZN(n883) );
  NOR2_X1 U558 ( .A1(n614), .A2(G651), .ZN(n641) );
  AND2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n879) );
  NAND2_X1 U560 ( .A1(n879), .A2(G113), .ZN(n519) );
  NOR2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n516) );
  XOR2_X1 U562 ( .A(KEYINPUT17), .B(n516), .Z(n517) );
  NAND2_X1 U563 ( .A1(G137), .A2(n883), .ZN(n518) );
  AND2_X1 U564 ( .A1(n519), .A2(n518), .ZN(n682) );
  INV_X1 U565 ( .A(G2104), .ZN(n523) );
  NOR2_X1 U566 ( .A1(n523), .A2(G2105), .ZN(n520) );
  XNOR2_X2 U567 ( .A(n520), .B(KEYINPUT66), .ZN(n886) );
  NAND2_X1 U568 ( .A1(G101), .A2(n886), .ZN(n522) );
  INV_X1 U569 ( .A(KEYINPUT23), .ZN(n521) );
  XNOR2_X1 U570 ( .A(n522), .B(n521), .ZN(n526) );
  NAND2_X1 U571 ( .A1(n523), .A2(G2105), .ZN(n524) );
  XNOR2_X1 U572 ( .A(n524), .B(KEYINPUT65), .ZN(n878) );
  NAND2_X1 U573 ( .A1(n878), .A2(G125), .ZN(n525) );
  NAND2_X1 U574 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U575 ( .A(n527), .B(KEYINPUT67), .ZN(n683) );
  AND2_X1 U576 ( .A1(n682), .A2(n683), .ZN(G160) );
  XOR2_X1 U577 ( .A(KEYINPUT0), .B(G543), .Z(n614) );
  NAND2_X1 U578 ( .A1(G52), .A2(n641), .ZN(n528) );
  XOR2_X1 U579 ( .A(KEYINPUT70), .B(n528), .Z(n539) );
  INV_X1 U580 ( .A(G651), .ZN(n533) );
  NOR2_X1 U581 ( .A1(n614), .A2(n533), .ZN(n635) );
  NAND2_X1 U582 ( .A1(n635), .A2(G77), .ZN(n531) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n529) );
  XNOR2_X1 U584 ( .A(n529), .B(KEYINPUT64), .ZN(n636) );
  NAND2_X1 U585 ( .A1(G90), .A2(n636), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U587 ( .A(n532), .B(KEYINPUT9), .ZN(n537) );
  NOR2_X1 U588 ( .A1(G543), .A2(n533), .ZN(n535) );
  XNOR2_X1 U589 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n534) );
  XNOR2_X1 U590 ( .A(n535), .B(n534), .ZN(n640) );
  NAND2_X1 U591 ( .A1(G64), .A2(n640), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U593 ( .A1(n539), .A2(n538), .ZN(G171) );
  INV_X1 U594 ( .A(G171), .ZN(G301) );
  XOR2_X1 U595 ( .A(KEYINPUT79), .B(KEYINPUT18), .Z(n541) );
  NAND2_X1 U596 ( .A1(G123), .A2(n878), .ZN(n540) );
  XNOR2_X1 U597 ( .A(n541), .B(n540), .ZN(n548) );
  NAND2_X1 U598 ( .A1(n879), .A2(G111), .ZN(n543) );
  NAND2_X1 U599 ( .A1(G99), .A2(n886), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n883), .A2(G135), .ZN(n544) );
  XOR2_X1 U602 ( .A(KEYINPUT80), .B(n544), .Z(n545) );
  NOR2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n923) );
  XNOR2_X1 U605 ( .A(G2096), .B(n923), .ZN(n549) );
  OR2_X1 U606 ( .A1(G2100), .A2(n549), .ZN(G156) );
  INV_X1 U607 ( .A(G69), .ZN(G235) );
  NAND2_X1 U608 ( .A1(G94), .A2(G452), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n550), .B(KEYINPUT71), .ZN(G173) );
  XOR2_X1 U610 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n552) );
  NAND2_X1 U611 ( .A1(G7), .A2(G661), .ZN(n551) );
  XNOR2_X1 U612 ( .A(n552), .B(n551), .ZN(G223) );
  XOR2_X1 U613 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n554) );
  INV_X1 U614 ( .A(G223), .ZN(n830) );
  NAND2_X1 U615 ( .A1(G567), .A2(n830), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n554), .B(n553), .ZN(G234) );
  NAND2_X1 U617 ( .A1(G56), .A2(n640), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT14), .B(n555), .Z(n561) );
  NAND2_X1 U619 ( .A1(G81), .A2(n636), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n556), .B(KEYINPUT12), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G68), .A2(n635), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U623 ( .A(KEYINPUT13), .B(n559), .Z(n560) );
  NOR2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n641), .A2(G43), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n998) );
  INV_X1 U627 ( .A(G860), .ZN(n596) );
  OR2_X1 U628 ( .A1(n998), .A2(n596), .ZN(G153) );
  NAND2_X1 U629 ( .A1(G868), .A2(G301), .ZN(n572) );
  NAND2_X1 U630 ( .A1(G66), .A2(n640), .ZN(n565) );
  NAND2_X1 U631 ( .A1(G92), .A2(n636), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G79), .A2(n635), .ZN(n567) );
  NAND2_X1 U634 ( .A1(G54), .A2(n641), .ZN(n566) );
  NAND2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT15), .B(n570), .Z(n993) );
  OR2_X1 U638 ( .A1(n993), .A2(G868), .ZN(n571) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(G284) );
  NAND2_X1 U640 ( .A1(G65), .A2(n640), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G53), .A2(n641), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT72), .B(n575), .Z(n579) );
  NAND2_X1 U644 ( .A1(n636), .A2(G91), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n635), .A2(G78), .ZN(n576) );
  AND2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(G299) );
  NAND2_X1 U648 ( .A1(G89), .A2(n636), .ZN(n580) );
  XNOR2_X1 U649 ( .A(KEYINPUT4), .B(n580), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n635), .A2(G76), .ZN(n581) );
  XOR2_X1 U651 ( .A(KEYINPUT75), .B(n581), .Z(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U653 ( .A(n584), .B(KEYINPUT5), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G63), .A2(n640), .ZN(n586) );
  NAND2_X1 U655 ( .A1(G51), .A2(n641), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U657 ( .A(KEYINPUT6), .B(n587), .Z(n588) );
  NAND2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U659 ( .A(n590), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U660 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U661 ( .A1(G868), .A2(G299), .ZN(n591) );
  XOR2_X1 U662 ( .A(KEYINPUT77), .B(n591), .Z(n595) );
  INV_X1 U663 ( .A(G868), .ZN(n592) );
  NOR2_X1 U664 ( .A1(G286), .A2(n592), .ZN(n593) );
  XNOR2_X1 U665 ( .A(KEYINPUT76), .B(n593), .ZN(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U667 ( .A1(G559), .A2(n596), .ZN(n597) );
  XNOR2_X1 U668 ( .A(KEYINPUT78), .B(n597), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n598), .A2(n993), .ZN(n599) );
  XNOR2_X1 U670 ( .A(KEYINPUT16), .B(n599), .ZN(G148) );
  NOR2_X1 U671 ( .A1(G868), .A2(n998), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G868), .A2(n993), .ZN(n600) );
  NOR2_X1 U673 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U674 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U675 ( .A1(n993), .A2(G559), .ZN(n654) );
  XNOR2_X1 U676 ( .A(n998), .B(n654), .ZN(n603) );
  NOR2_X1 U677 ( .A1(n603), .A2(G860), .ZN(n611) );
  NAND2_X1 U678 ( .A1(n635), .A2(G80), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G93), .A2(n636), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n610) );
  NAND2_X1 U681 ( .A1(G67), .A2(n640), .ZN(n607) );
  NAND2_X1 U682 ( .A1(G55), .A2(n641), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U684 ( .A(KEYINPUT81), .B(n608), .Z(n609) );
  NOR2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n656) );
  XNOR2_X1 U686 ( .A(n611), .B(n656), .ZN(G145) );
  NAND2_X1 U687 ( .A1(G74), .A2(G651), .ZN(n612) );
  XNOR2_X1 U688 ( .A(KEYINPUT83), .B(n612), .ZN(n613) );
  NOR2_X1 U689 ( .A1(n640), .A2(n613), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n614), .A2(G87), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n641), .A2(G49), .ZN(n617) );
  XOR2_X1 U693 ( .A(KEYINPUT82), .B(n617), .Z(n618) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U695 ( .A(KEYINPUT84), .B(n620), .Z(G288) );
  NAND2_X1 U696 ( .A1(n641), .A2(G48), .ZN(n627) );
  NAND2_X1 U697 ( .A1(G61), .A2(n640), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G86), .A2(n636), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n635), .A2(G73), .ZN(n623) );
  XOR2_X1 U701 ( .A(KEYINPUT2), .B(n623), .Z(n624) );
  NOR2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U704 ( .A(KEYINPUT85), .B(n628), .Z(G305) );
  AND2_X1 U705 ( .A1(n640), .A2(G60), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n635), .A2(G72), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G85), .A2(n636), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n641), .A2(G47), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(G290) );
  NAND2_X1 U712 ( .A1(n635), .A2(G75), .ZN(n638) );
  NAND2_X1 U713 ( .A1(G88), .A2(n636), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U715 ( .A(KEYINPUT86), .B(n639), .Z(n645) );
  NAND2_X1 U716 ( .A1(G62), .A2(n640), .ZN(n643) );
  NAND2_X1 U717 ( .A1(G50), .A2(n641), .ZN(n642) );
  AND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n645), .A2(n644), .ZN(G303) );
  INV_X1 U720 ( .A(G303), .ZN(G166) );
  INV_X1 U721 ( .A(G299), .ZN(n984) );
  XNOR2_X1 U722 ( .A(n984), .B(n656), .ZN(n652) );
  XNOR2_X1 U723 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n647) );
  XNOR2_X1 U724 ( .A(G305), .B(KEYINPUT19), .ZN(n646) );
  XNOR2_X1 U725 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U726 ( .A(G288), .B(n648), .ZN(n650) );
  XNOR2_X1 U727 ( .A(G290), .B(G166), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U729 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(n998), .ZN(n900) );
  XOR2_X1 U731 ( .A(n900), .B(n654), .Z(n655) );
  NAND2_X1 U732 ( .A1(G868), .A2(n655), .ZN(n658) );
  OR2_X1 U733 ( .A1(n656), .A2(G868), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n658), .A2(n657), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2078), .A2(G2084), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n659), .B(KEYINPUT20), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n660), .B(KEYINPUT89), .ZN(n661) );
  NAND2_X1 U738 ( .A1(n661), .A2(G2090), .ZN(n662) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U741 ( .A(KEYINPUT90), .B(G44), .ZN(n664) );
  XNOR2_X1 U742 ( .A(n664), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U743 ( .A1(G120), .A2(G108), .ZN(n665) );
  NOR2_X1 U744 ( .A1(G235), .A2(n665), .ZN(n666) );
  NAND2_X1 U745 ( .A1(G57), .A2(n666), .ZN(n836) );
  NAND2_X1 U746 ( .A1(G567), .A2(n836), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n667), .B(KEYINPUT92), .ZN(n673) );
  XOR2_X1 U748 ( .A(KEYINPUT91), .B(KEYINPUT22), .Z(n669) );
  NAND2_X1 U749 ( .A1(G132), .A2(G82), .ZN(n668) );
  XNOR2_X1 U750 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X1 U751 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U752 ( .A1(G96), .A2(n671), .ZN(n837) );
  NAND2_X1 U753 ( .A1(G2106), .A2(n837), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n673), .A2(n672), .ZN(n857) );
  NAND2_X1 U755 ( .A1(G661), .A2(G483), .ZN(n674) );
  XOR2_X1 U756 ( .A(KEYINPUT93), .B(n674), .Z(n675) );
  NOR2_X1 U757 ( .A1(n857), .A2(n675), .ZN(n835) );
  NAND2_X1 U758 ( .A1(n835), .A2(G36), .ZN(G176) );
  NAND2_X1 U759 ( .A1(G102), .A2(n886), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G138), .A2(n883), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n681) );
  NAND2_X1 U762 ( .A1(G126), .A2(n878), .ZN(n679) );
  NAND2_X1 U763 ( .A1(G114), .A2(n879), .ZN(n678) );
  NAND2_X1 U764 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U765 ( .A1(n681), .A2(n680), .ZN(G164) );
  XNOR2_X1 U766 ( .A(G1986), .B(G290), .ZN(n990) );
  AND2_X1 U767 ( .A1(n682), .A2(G40), .ZN(n684) );
  NAND2_X1 U768 ( .A1(n684), .A2(n683), .ZN(n686) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n688) );
  NOR2_X1 U770 ( .A1(n686), .A2(n688), .ZN(n685) );
  XNOR2_X1 U771 ( .A(n685), .B(KEYINPUT94), .ZN(n815) );
  NAND2_X1 U772 ( .A1(n990), .A2(n815), .ZN(n805) );
  INV_X1 U773 ( .A(n686), .ZN(n687) );
  NAND2_X1 U774 ( .A1(G8), .A2(n732), .ZN(n765) );
  NOR2_X1 U775 ( .A1(G1981), .A2(G305), .ZN(n689) );
  XOR2_X1 U776 ( .A(n689), .B(KEYINPUT24), .Z(n690) );
  NOR2_X1 U777 ( .A1(n765), .A2(n690), .ZN(n770) );
  INV_X1 U778 ( .A(n732), .ZN(n715) );
  AND2_X1 U779 ( .A1(n715), .A2(G1996), .ZN(n691) );
  XOR2_X1 U780 ( .A(n691), .B(KEYINPUT26), .Z(n693) );
  NAND2_X1 U781 ( .A1(n732), .A2(G1341), .ZN(n692) );
  NAND2_X1 U782 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U783 ( .A1(n998), .A2(n694), .ZN(n695) );
  OR2_X1 U784 ( .A1(n993), .A2(n695), .ZN(n702) );
  NAND2_X1 U785 ( .A1(n993), .A2(n695), .ZN(n700) );
  INV_X1 U786 ( .A(G2067), .ZN(n964) );
  NOR2_X1 U787 ( .A1(n732), .A2(n964), .ZN(n696) );
  XOR2_X1 U788 ( .A(n696), .B(KEYINPUT102), .Z(n698) );
  NAND2_X1 U789 ( .A1(n732), .A2(G1348), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n702), .A2(n701), .ZN(n708) );
  NAND2_X1 U793 ( .A1(G2072), .A2(n715), .ZN(n703) );
  XNOR2_X1 U794 ( .A(n703), .B(KEYINPUT100), .ZN(n704) );
  XNOR2_X1 U795 ( .A(KEYINPUT27), .B(n704), .ZN(n706) );
  AND2_X1 U796 ( .A1(n732), .A2(G1956), .ZN(n705) );
  NOR2_X1 U797 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U798 ( .A1(n984), .A2(n709), .ZN(n707) );
  NAND2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n713) );
  NOR2_X1 U800 ( .A1(n984), .A2(n709), .ZN(n711) );
  XNOR2_X1 U801 ( .A(KEYINPUT101), .B(KEYINPUT28), .ZN(n710) );
  XNOR2_X1 U802 ( .A(n711), .B(n710), .ZN(n712) );
  NAND2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U804 ( .A(n714), .B(KEYINPUT29), .ZN(n719) );
  XOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .Z(n968) );
  NOR2_X1 U806 ( .A1(n968), .A2(n732), .ZN(n717) );
  NOR2_X1 U807 ( .A1(n715), .A2(G1961), .ZN(n716) );
  NOR2_X1 U808 ( .A1(n717), .A2(n716), .ZN(n720) );
  NOR2_X1 U809 ( .A1(G301), .A2(n720), .ZN(n718) );
  NOR2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n730) );
  AND2_X1 U811 ( .A1(G301), .A2(n720), .ZN(n727) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n765), .ZN(n743) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n732), .ZN(n741) );
  NOR2_X1 U814 ( .A1(n743), .A2(n741), .ZN(n721) );
  NAND2_X1 U815 ( .A1(G8), .A2(n721), .ZN(n724) );
  NOR2_X1 U816 ( .A1(G168), .A2(n725), .ZN(n726) );
  NOR2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U818 ( .A(n728), .B(KEYINPUT31), .ZN(n729) );
  NOR2_X1 U819 ( .A1(n730), .A2(n729), .ZN(n742) );
  INV_X1 U820 ( .A(n742), .ZN(n731) );
  NAND2_X1 U821 ( .A1(G286), .A2(n731), .ZN(n737) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n765), .ZN(n734) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U825 ( .A1(n735), .A2(G303), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U827 ( .A1(n738), .A2(G8), .ZN(n740) );
  NAND2_X1 U828 ( .A1(n741), .A2(G8), .ZN(n745) );
  NOR2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n761) );
  NAND2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n994) );
  INV_X1 U832 ( .A(n994), .ZN(n746) );
  OR2_X1 U833 ( .A1(n746), .A2(n765), .ZN(n750) );
  INV_X1 U834 ( .A(n750), .ZN(n747) );
  AND2_X1 U835 ( .A1(n761), .A2(n747), .ZN(n748) );
  AND2_X1 U836 ( .A1(n760), .A2(n748), .ZN(n754) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n755) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U839 ( .A1(n755), .A2(n749), .ZN(n985) );
  OR2_X1 U840 ( .A1(n750), .A2(n985), .ZN(n752) );
  INV_X1 U841 ( .A(KEYINPUT33), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n759) );
  NAND2_X1 U844 ( .A1(n755), .A2(KEYINPUT33), .ZN(n756) );
  OR2_X1 U845 ( .A1(n765), .A2(n756), .ZN(n757) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n999) );
  NAND2_X1 U847 ( .A1(n757), .A2(n999), .ZN(n758) );
  OR2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n768) );
  NAND2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n764) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U851 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U855 ( .A1(n770), .A2(n769), .ZN(n803) );
  XNOR2_X1 U856 ( .A(KEYINPUT37), .B(G2067), .ZN(n813) );
  NAND2_X1 U857 ( .A1(G104), .A2(n886), .ZN(n771) );
  XOR2_X1 U858 ( .A(KEYINPUT95), .B(n771), .Z(n773) );
  NAND2_X1 U859 ( .A1(G140), .A2(n883), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U861 ( .A(KEYINPUT34), .B(n774), .ZN(n781) );
  NAND2_X1 U862 ( .A1(n879), .A2(G116), .ZN(n775) );
  XNOR2_X1 U863 ( .A(KEYINPUT97), .B(n775), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n878), .A2(G128), .ZN(n776) );
  XOR2_X1 U865 ( .A(KEYINPUT96), .B(n776), .Z(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U867 ( .A(n779), .B(KEYINPUT35), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U869 ( .A(KEYINPUT36), .B(n782), .ZN(n896) );
  NOR2_X1 U870 ( .A1(n813), .A2(n896), .ZN(n935) );
  NAND2_X1 U871 ( .A1(n935), .A2(n815), .ZN(n811) );
  INV_X1 U872 ( .A(n815), .ZN(n800) );
  NAND2_X1 U873 ( .A1(n879), .A2(G117), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G141), .A2(n883), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n886), .A2(G105), .ZN(n785) );
  XOR2_X1 U877 ( .A(KEYINPUT38), .B(n785), .Z(n786) );
  NOR2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n878), .A2(G129), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n876) );
  NAND2_X1 U881 ( .A1(n876), .A2(G1996), .ZN(n798) );
  NAND2_X1 U882 ( .A1(n879), .A2(G107), .ZN(n791) );
  NAND2_X1 U883 ( .A1(G131), .A2(n883), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n878), .A2(G119), .ZN(n792) );
  XOR2_X1 U886 ( .A(KEYINPUT98), .B(n792), .Z(n793) );
  NOR2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G95), .A2(n886), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n874) );
  NAND2_X1 U890 ( .A1(G1991), .A2(n874), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U892 ( .A(n799), .B(KEYINPUT99), .ZN(n932) );
  NOR2_X1 U893 ( .A1(n800), .A2(n932), .ZN(n808) );
  INV_X1 U894 ( .A(n808), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n811), .A2(n801), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n818) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n876), .ZN(n921) );
  NOR2_X1 U899 ( .A1(G1991), .A2(n874), .ZN(n925) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n925), .A2(n806), .ZN(n807) );
  NOR2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n921), .A2(n809), .ZN(n810) );
  XNOR2_X1 U904 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n813), .A2(n896), .ZN(n918) );
  NAND2_X1 U907 ( .A1(n814), .A2(n918), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n819), .ZN(G329) );
  XOR2_X1 U911 ( .A(G2454), .B(G2435), .Z(n821) );
  XNOR2_X1 U912 ( .A(G2438), .B(G2427), .ZN(n820) );
  XNOR2_X1 U913 ( .A(n821), .B(n820), .ZN(n828) );
  XOR2_X1 U914 ( .A(KEYINPUT105), .B(G2446), .Z(n823) );
  XNOR2_X1 U915 ( .A(G2443), .B(G2430), .ZN(n822) );
  XNOR2_X1 U916 ( .A(n823), .B(n822), .ZN(n824) );
  XOR2_X1 U917 ( .A(n824), .B(G2451), .Z(n826) );
  XNOR2_X1 U918 ( .A(G1348), .B(G1341), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n826), .B(n825), .ZN(n827) );
  XNOR2_X1 U920 ( .A(n828), .B(n827), .ZN(n829) );
  NAND2_X1 U921 ( .A1(n829), .A2(G14), .ZN(n907) );
  XOR2_X1 U922 ( .A(KEYINPUT106), .B(n907), .Z(G401) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n830), .ZN(G217) );
  NAND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n832) );
  INV_X1 U925 ( .A(G661), .ZN(n831) );
  NOR2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U927 ( .A(n833), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(G188) );
  XOR2_X1 U930 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  XOR2_X1 U931 ( .A(G108), .B(KEYINPUT118), .Z(G238) );
  INV_X1 U933 ( .A(G132), .ZN(G219) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  INV_X1 U935 ( .A(G82), .ZN(G220) );
  NOR2_X1 U936 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XOR2_X1 U938 ( .A(KEYINPUT110), .B(G1976), .Z(n839) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1961), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n840), .B(KEYINPUT41), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U944 ( .A(G1981), .B(G1966), .Z(n844) );
  XNOR2_X1 U945 ( .A(G1971), .B(G1956), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U947 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U948 ( .A(G2474), .B(KEYINPUT111), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(G229) );
  XOR2_X1 U950 ( .A(G2100), .B(G2096), .Z(n850) );
  XNOR2_X1 U951 ( .A(KEYINPUT42), .B(G2678), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U953 ( .A(KEYINPUT43), .B(G2072), .Z(n852) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U956 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U957 ( .A(G2078), .B(G2084), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(G227) );
  XNOR2_X1 U959 ( .A(KEYINPUT109), .B(n857), .ZN(G319) );
  NAND2_X1 U960 ( .A1(G124), .A2(n878), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n858), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G100), .A2(n886), .ZN(n860) );
  NAND2_X1 U963 ( .A1(G136), .A2(n883), .ZN(n859) );
  NAND2_X1 U964 ( .A1(n860), .A2(n859), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n879), .A2(G112), .ZN(n861) );
  XOR2_X1 U966 ( .A(KEYINPUT112), .B(n861), .Z(n862) );
  NOR2_X1 U967 ( .A1(n863), .A2(n862), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U969 ( .A(KEYINPUT113), .B(n866), .ZN(G162) );
  NAND2_X1 U970 ( .A1(G130), .A2(n878), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G118), .A2(n879), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G106), .A2(n886), .ZN(n870) );
  NAND2_X1 U974 ( .A1(G142), .A2(n883), .ZN(n869) );
  NAND2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U976 ( .A(n871), .B(KEYINPUT45), .Z(n872) );
  NOR2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n875) );
  XNOR2_X1 U978 ( .A(n875), .B(n874), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n877), .B(n876), .ZN(n892) );
  NAND2_X1 U980 ( .A1(G127), .A2(n878), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G115), .A2(n879), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n882), .B(KEYINPUT47), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G139), .A2(n883), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n889) );
  NAND2_X1 U986 ( .A1(n886), .A2(G103), .ZN(n887) );
  XOR2_X1 U987 ( .A(KEYINPUT114), .B(n887), .Z(n888) );
  NOR2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n913) );
  XNOR2_X1 U989 ( .A(G160), .B(n913), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n890), .B(n923), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n898) );
  XOR2_X1 U992 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n894) );
  XNOR2_X1 U993 ( .A(G164), .B(G162), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U997 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U998 ( .A(G286), .B(n993), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1000 ( .A(G301), .B(n902), .Z(n903) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n903), .ZN(n904) );
  XOR2_X1 U1002 ( .A(KEYINPUT115), .B(n904), .Z(G397) );
  XNOR2_X1 U1003 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G229), .A2(G227), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n907), .ZN(n908) );
  NOR2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1008 ( .A(KEYINPUT117), .B(n910), .Z(n912) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G57), .ZN(G237) );
  INV_X1 U1013 ( .A(G29), .ZN(n940) );
  XNOR2_X1 U1014 ( .A(KEYINPUT121), .B(KEYINPUT52), .ZN(n937) );
  XOR2_X1 U1015 ( .A(G2072), .B(n913), .Z(n915) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n914) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1018 ( .A(KEYINPUT120), .B(n916), .ZN(n917) );
  XNOR2_X1 U1019 ( .A(n917), .B(KEYINPUT50), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n931) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n920) );
  NOR2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1023 ( .A(KEYINPUT51), .B(n922), .Z(n929) );
  XNOR2_X1 U1024 ( .A(G160), .B(G2084), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1027 ( .A(KEYINPUT119), .B(n927), .Z(n928) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(n937), .B(n936), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n981) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n981), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n1018) );
  XNOR2_X1 U1036 ( .A(G1971), .B(G22), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(G1976), .B(G23), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1039 ( .A(KEYINPUT126), .B(n943), .Z(n945) );
  XNOR2_X1 U1040 ( .A(G1986), .B(G24), .ZN(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT58), .B(n946), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(G1961), .B(G5), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G1966), .B(G21), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n961) );
  XNOR2_X1 U1047 ( .A(G1956), .B(G20), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(G1341), .B(G19), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(G1981), .B(G6), .ZN(n951) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(KEYINPUT125), .B(n953), .ZN(n954) );
  NOR2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G1348), .B(KEYINPUT59), .ZN(n956) );
  XNOR2_X1 U1054 ( .A(n956), .B(G4), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(KEYINPUT60), .B(n959), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1058 ( .A(KEYINPUT61), .B(n962), .Z(n963) );
  NOR2_X1 U1059 ( .A1(G16), .A2(n963), .ZN(n1015) );
  XNOR2_X1 U1060 ( .A(G26), .B(n964), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n965), .A2(G28), .ZN(n974) );
  XNOR2_X1 U1062 ( .A(G1996), .B(G32), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(G33), .B(G2072), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(G1991), .B(G25), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(G27), .B(n968), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1070 ( .A(KEYINPUT53), .B(n975), .Z(n978) );
  XOR2_X1 U1071 ( .A(G34), .B(KEYINPUT54), .Z(n976) );
  XNOR2_X1 U1072 ( .A(G2084), .B(n976), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(G35), .B(G2090), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n982) );
  XOR2_X1 U1076 ( .A(n982), .B(n981), .Z(n983) );
  NOR2_X1 U1077 ( .A1(G29), .A2(n983), .ZN(n1012) );
  XOR2_X1 U1078 ( .A(KEYINPUT56), .B(G16), .Z(n1010) );
  XNOR2_X1 U1079 ( .A(n984), .B(G1956), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n1008) );
  XNOR2_X1 U1081 ( .A(G1961), .B(G171), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(n987), .B(KEYINPUT124), .ZN(n992) );
  INV_X1 U1083 ( .A(G1971), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(G166), .A2(n988), .ZN(n989) );
  NOR2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(G1348), .B(n993), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(n998), .B(G1341), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G168), .B(G1966), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n1001), .B(KEYINPUT57), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(KEYINPUT123), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(G11), .A2(n1013), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(n1016), .B(KEYINPUT127), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1019), .ZN(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

