

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814;

  AND2_X1 U374 ( .A1(n734), .A2(n369), .ZN(n603) );
  NOR2_X1 U375 ( .A1(n598), .A2(n760), .ZN(n384) );
  BUF_X1 U376 ( .A(n659), .Z(n354) );
  XNOR2_X1 U377 ( .A(n532), .B(KEYINPUT67), .ZN(n533) );
  INV_X1 U378 ( .A(n750), .ZN(n595) );
  NAND2_X2 U379 ( .A1(n626), .A2(n754), .ZN(n750) );
  XNOR2_X1 U380 ( .A(n537), .B(KEYINPUT16), .ZN(n357) );
  NAND2_X2 U381 ( .A1(n678), .A2(G953), .ZN(n714) );
  XNOR2_X2 U382 ( .A(n612), .B(KEYINPUT79), .ZN(n427) );
  XNOR2_X2 U383 ( .A(n555), .B(KEYINPUT70), .ZN(n556) );
  XNOR2_X2 U384 ( .A(n622), .B(n621), .ZN(n687) );
  XNOR2_X2 U385 ( .A(n536), .B(n789), .ZN(n490) );
  NAND2_X1 U386 ( .A1(n387), .A2(n467), .ZN(n386) );
  NOR2_X1 U387 ( .A1(n589), .A2(KEYINPUT91), .ZN(n582) );
  XNOR2_X2 U388 ( .A(n490), .B(n489), .ZN(n709) );
  XNOR2_X1 U389 ( .A(n636), .B(KEYINPUT19), .ZN(n623) );
  NOR2_X2 U390 ( .A1(n623), .A2(n366), .ZN(n423) );
  XOR2_X2 U391 ( .A(KEYINPUT62), .B(n688), .Z(n689) );
  XNOR2_X2 U392 ( .A(n554), .B(n477), .ZN(n702) );
  XOR2_X2 U393 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n374) );
  NAND2_X2 U394 ( .A1(n386), .A2(n389), .ZN(n422) );
  OR2_X2 U395 ( .A1(n688), .A2(G902), .ZN(n546) );
  XNOR2_X2 U396 ( .A(n711), .B(n710), .ZN(n712) );
  AND2_X4 U397 ( .A1(n394), .A2(n665), .ZN(n801) );
  XOR2_X2 U398 ( .A(n663), .B(KEYINPUT38), .Z(n363) );
  XNOR2_X1 U399 ( .A(n355), .B(KEYINPUT102), .ZN(n390) );
  NOR2_X2 U400 ( .A1(n608), .A2(n682), .ZN(n355) );
  NAND2_X1 U401 ( .A1(n356), .A2(KEYINPUT77), .ZN(n419) );
  NAND2_X1 U402 ( .A1(n438), .A2(n421), .ZN(n356) );
  XNOR2_X2 U403 ( .A(n357), .B(n481), .ZN(n789) );
  INV_X2 U404 ( .A(G953), .ZN(n808) );
  XNOR2_X2 U405 ( .A(n757), .B(n548), .ZN(n659) );
  NAND2_X2 U406 ( .A1(n427), .A2(n616), .ZN(n617) );
  INV_X1 U407 ( .A(n629), .ZN(n440) );
  NOR2_X2 U408 ( .A1(n673), .A2(n672), .ZN(n385) );
  AND2_X1 U409 ( .A1(n392), .A2(n390), .ZN(n389) );
  NOR2_X1 U410 ( .A1(n687), .A2(n439), .ZN(n437) );
  NAND2_X1 U411 ( .A1(n443), .A2(n441), .ZN(n383) );
  XNOR2_X1 U412 ( .A(n585), .B(KEYINPUT33), .ZN(n746) );
  NAND2_X1 U413 ( .A1(n671), .A2(KEYINPUT2), .ZN(n673) );
  BUF_X1 U414 ( .A(n378), .Z(n358) );
  NOR2_X2 U415 ( .A1(n674), .A2(n385), .ZN(n378) );
  NOR2_X2 U416 ( .A1(n674), .A2(n385), .ZN(n379) );
  XNOR2_X2 U417 ( .A(n395), .B(n654), .ZN(n394) );
  XNOR2_X2 U418 ( .A(n798), .B(G146), .ZN(n554) );
  XNOR2_X2 U419 ( .A(n536), .B(n535), .ZN(n798) );
  INV_X1 U420 ( .A(KEYINPUT66), .ZN(n476) );
  XNOR2_X1 U421 ( .A(n633), .B(n632), .ZN(n635) );
  INV_X1 U422 ( .A(G237), .ZN(n491) );
  NAND2_X1 U423 ( .A1(n419), .A2(n418), .ZN(n414) );
  NAND2_X1 U424 ( .A1(n416), .A2(n413), .ZN(n399) );
  AND2_X1 U425 ( .A1(n415), .A2(n812), .ZN(n413) );
  NOR2_X1 U426 ( .A1(n426), .A2(KEYINPUT77), .ZN(n417) );
  NAND2_X1 U427 ( .A1(n455), .A2(KEYINPUT92), .ZN(n447) );
  NOR2_X1 U428 ( .A1(G953), .A2(G237), .ZN(n538) );
  INV_X1 U429 ( .A(n683), .ZN(n467) );
  INV_X1 U430 ( .A(G104), .ZN(n479) );
  INV_X1 U431 ( .A(KEYINPUT78), .ZN(n433) );
  XOR2_X1 U432 ( .A(G122), .B(G116), .Z(n505) );
  XNOR2_X1 U433 ( .A(G134), .B(G107), .ZN(n504) );
  OR2_X1 U434 ( .A1(n579), .A2(n476), .ZN(n471) );
  AND2_X1 U435 ( .A1(n579), .A2(n476), .ZN(n472) );
  XOR2_X1 U436 ( .A(n675), .B(KEYINPUT59), .Z(n676) );
  AND2_X1 U437 ( .A1(n406), .A2(n360), .ZN(n403) );
  NAND2_X1 U438 ( .A1(n359), .A2(n407), .ZN(n406) );
  AND2_X1 U439 ( .A1(n635), .A2(n434), .ZN(n436) );
  NOR2_X1 U440 ( .A1(n435), .A2(KEYINPUT82), .ZN(n434) );
  INV_X1 U441 ( .A(n634), .ZN(n435) );
  INV_X1 U442 ( .A(KEYINPUT65), .ZN(n464) );
  NAND2_X1 U443 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U444 ( .A1(n383), .A2(n611), .ZN(n612) );
  NAND2_X1 U445 ( .A1(n397), .A2(n396), .ZN(n395) );
  NAND2_X1 U446 ( .A1(n400), .A2(n399), .ZN(n396) );
  NAND2_X1 U447 ( .A1(n373), .A2(n463), .ZN(n462) );
  NAND2_X1 U448 ( .A1(n669), .A2(n464), .ZN(n463) );
  OR2_X1 U449 ( .A1(n373), .A2(KEYINPUT65), .ZN(n465) );
  XNOR2_X1 U450 ( .A(G134), .B(G131), .ZN(n535) );
  XNOR2_X1 U451 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n484) );
  NAND2_X1 U452 ( .A1(n412), .A2(n411), .ZN(n585) );
  NOR2_X1 U453 ( .A1(n659), .A2(n750), .ZN(n412) );
  NAND2_X1 U454 ( .A1(n492), .A2(n459), .ZN(n454) );
  NAND2_X1 U455 ( .A1(n453), .A2(n669), .ZN(n452) );
  INV_X1 U456 ( .A(n492), .ZN(n453) );
  INV_X1 U457 ( .A(G902), .ZN(n570) );
  XNOR2_X1 U458 ( .A(G101), .B(G113), .ZN(n539) );
  XNOR2_X1 U459 ( .A(n483), .B(G101), .ZN(n790) );
  XNOR2_X1 U460 ( .A(G110), .B(G107), .ZN(n483) );
  XOR2_X1 U461 ( .A(G119), .B(KEYINPUT84), .Z(n562) );
  XNOR2_X1 U462 ( .A(G140), .B(G137), .ZN(n566) );
  XNOR2_X1 U463 ( .A(G104), .B(KEYINPUT80), .ZN(n550) );
  NAND2_X1 U464 ( .A1(G237), .A2(G234), .ZN(n494) );
  XNOR2_X1 U465 ( .A(n647), .B(n646), .ZN(n656) );
  XNOR2_X1 U466 ( .A(n510), .B(n509), .ZN(n698) );
  NAND2_X1 U467 ( .A1(n656), .A2(n730), .ZN(n428) );
  INV_X1 U468 ( .A(n619), .ZN(n456) );
  INV_X1 U469 ( .A(KEYINPUT32), .ZN(n474) );
  AND2_X1 U470 ( .A1(n471), .A2(n580), .ZN(n470) );
  INV_X1 U471 ( .A(KEYINPUT60), .ZN(n430) );
  NOR2_X1 U472 ( .A1(n767), .A2(KEYINPUT47), .ZN(n359) );
  OR2_X1 U473 ( .A1(n634), .A2(n439), .ZN(n360) );
  AND2_X1 U474 ( .A1(n665), .A2(n371), .ZN(n361) );
  AND2_X1 U475 ( .A1(n454), .A2(n450), .ZN(n362) );
  XNOR2_X1 U476 ( .A(G902), .B(KEYINPUT15), .ZN(n669) );
  INV_X1 U477 ( .A(n584), .ZN(n411) );
  NOR2_X1 U478 ( .A1(n618), .A2(n619), .ZN(n364) );
  OR2_X1 U479 ( .A1(n455), .A2(KEYINPUT92), .ZN(n365) );
  NAND2_X1 U480 ( .A1(n610), .A2(n499), .ZN(n366) );
  AND2_X1 U481 ( .A1(n451), .A2(n454), .ZN(n367) );
  XNOR2_X1 U482 ( .A(n500), .B(KEYINPUT0), .ZN(n368) );
  OR2_X1 U483 ( .A1(n598), .A2(n597), .ZN(n369) );
  XOR2_X1 U484 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n370) );
  INV_X1 U485 ( .A(KEYINPUT82), .ZN(n439) );
  AND2_X1 U486 ( .A1(n459), .A2(KEYINPUT65), .ZN(n371) );
  XOR2_X1 U487 ( .A(KEYINPUT87), .B(KEYINPUT45), .Z(n372) );
  AND2_X1 U488 ( .A1(n466), .A2(n670), .ZN(n373) );
  AND2_X1 U489 ( .A1(KEYINPUT2), .A2(KEYINPUT86), .ZN(n375) );
  AND2_X1 U490 ( .A1(n373), .A2(n464), .ZN(n376) );
  NAND2_X1 U491 ( .A1(n465), .A2(n462), .ZN(n377) );
  BUF_X1 U492 ( .A(n428), .Z(n380) );
  NOR2_X1 U493 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X2 U494 ( .A1(n607), .A2(n606), .ZN(n682) );
  XNOR2_X1 U495 ( .A(n617), .B(n433), .ZN(n381) );
  XNOR2_X1 U496 ( .A(n617), .B(n433), .ZN(n620) );
  NAND2_X1 U497 ( .A1(n425), .A2(n424), .ZN(n388) );
  NOR2_X1 U498 ( .A1(n757), .A2(n637), .ZN(n409) );
  XNOR2_X1 U499 ( .A(n380), .B(n374), .ZN(n382) );
  XNOR2_X1 U500 ( .A(n428), .B(n374), .ZN(n410) );
  XNOR2_X1 U501 ( .A(n398), .B(n653), .ZN(n397) );
  AND2_X1 U502 ( .A1(n402), .A2(n377), .ZN(n461) );
  NAND2_X1 U503 ( .A1(n383), .A2(n757), .ZN(n597) );
  XNOR2_X1 U504 ( .A(n384), .B(KEYINPUT31), .ZN(n734) );
  NOR2_X1 U505 ( .A1(n739), .A2(n385), .ZN(n745) );
  NAND2_X1 U506 ( .A1(n388), .A2(KEYINPUT90), .ZN(n387) );
  NAND2_X1 U507 ( .A1(n393), .A2(n593), .ZN(n392) );
  NAND2_X1 U508 ( .A1(n589), .A2(n591), .ZN(n393) );
  AND2_X1 U509 ( .A1(n394), .A2(n361), .ZN(n401) );
  NAND2_X1 U510 ( .A1(n410), .A2(n652), .ZN(n398) );
  NAND2_X1 U511 ( .A1(n414), .A2(n812), .ZN(n400) );
  NAND2_X1 U512 ( .A1(n671), .A2(n801), .ZN(n666) );
  NAND2_X1 U513 ( .A1(n671), .A2(n401), .ZN(n402) );
  XNOR2_X2 U514 ( .A(n422), .B(n372), .ZN(n671) );
  NAND2_X1 U515 ( .A1(n404), .A2(n403), .ZN(n426) );
  NAND2_X1 U516 ( .A1(n405), .A2(KEYINPUT82), .ZN(n404) );
  INV_X1 U517 ( .A(n635), .ZN(n405) );
  INV_X1 U518 ( .A(n729), .ZN(n407) );
  NAND2_X1 U519 ( .A1(n408), .A2(n440), .ZN(n650) );
  XNOR2_X1 U520 ( .A(n409), .B(n628), .ZN(n408) );
  XNOR2_X1 U521 ( .A(n382), .B(G131), .ZN(G33) );
  NAND2_X1 U522 ( .A1(n577), .A2(n604), .ZN(n475) );
  XNOR2_X2 U523 ( .A(n534), .B(n533), .ZN(n604) );
  NAND2_X1 U524 ( .A1(n589), .A2(n581), .ZN(n424) );
  XNOR2_X1 U525 ( .A(n629), .B(n558), .ZN(n584) );
  XNOR2_X2 U526 ( .A(n557), .B(n556), .ZN(n629) );
  INV_X1 U527 ( .A(n437), .ZN(n415) );
  AND2_X1 U528 ( .A1(n438), .A2(n417), .ZN(n416) );
  NAND2_X1 U529 ( .A1(n437), .A2(KEYINPUT77), .ZN(n418) );
  INV_X1 U530 ( .A(n426), .ZN(n421) );
  XNOR2_X2 U531 ( .A(n423), .B(n368), .ZN(n583) );
  INV_X1 U532 ( .A(n582), .ZN(n425) );
  XNOR2_X1 U533 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U534 ( .A1(n620), .A2(n363), .ZN(n647) );
  NOR2_X2 U535 ( .A1(n686), .A2(n684), .ZN(n589) );
  XNOR2_X2 U536 ( .A(n475), .B(n474), .ZN(n686) );
  NAND2_X1 U537 ( .A1(n381), .A2(n364), .ZN(n622) );
  NAND2_X1 U538 ( .A1(n429), .A2(n596), .ZN(n443) );
  NAND2_X1 U539 ( .A1(n440), .A2(n595), .ZN(n429) );
  NOR2_X2 U540 ( .A1(n473), .A2(n469), .ZN(n684) );
  XNOR2_X1 U541 ( .A(n431), .B(n430), .ZN(G60) );
  NAND2_X1 U542 ( .A1(n679), .A2(n714), .ZN(n431) );
  XNOR2_X1 U543 ( .A(n565), .B(n564), .ZN(n569) );
  NAND2_X1 U544 ( .A1(n631), .A2(n630), .ZN(n729) );
  NAND2_X1 U545 ( .A1(n627), .A2(n754), .ZN(n637) );
  OR2_X2 U546 ( .A1(n702), .A2(G902), .ZN(n557) );
  XNOR2_X2 U547 ( .A(n432), .B(G143), .ZN(n506) );
  XNOR2_X2 U548 ( .A(G128), .B(KEYINPUT64), .ZN(n432) );
  NAND2_X1 U549 ( .A1(n436), .A2(n687), .ZN(n438) );
  NAND2_X1 U550 ( .A1(n595), .A2(n442), .ZN(n441) );
  NOR2_X1 U551 ( .A1(n629), .A2(n596), .ZN(n442) );
  NAND2_X1 U552 ( .A1(n444), .A2(n365), .ZN(n636) );
  NAND2_X1 U553 ( .A1(n446), .A2(n445), .ZN(n444) );
  NAND2_X1 U554 ( .A1(n449), .A2(KEYINPUT92), .ZN(n445) );
  NAND2_X1 U555 ( .A1(n448), .A2(n447), .ZN(n446) );
  INV_X1 U556 ( .A(n449), .ZN(n448) );
  NAND2_X1 U557 ( .A1(n709), .A2(n492), .ZN(n455) );
  NAND2_X1 U558 ( .A1(n367), .A2(n455), .ZN(n618) );
  NAND2_X1 U559 ( .A1(n451), .A2(n362), .ZN(n449) );
  INV_X1 U560 ( .A(n648), .ZN(n450) );
  OR2_X2 U561 ( .A1(n709), .A2(n452), .ZN(n451) );
  NAND2_X1 U562 ( .A1(n457), .A2(n456), .ZN(n588) );
  XNOR2_X1 U563 ( .A(n458), .B(n370), .ZN(n457) );
  NAND2_X1 U564 ( .A1(n746), .A2(n583), .ZN(n458) );
  NAND2_X1 U565 ( .A1(n461), .A2(n460), .ZN(n674) );
  INV_X1 U566 ( .A(n669), .ZN(n459) );
  NAND2_X1 U567 ( .A1(n666), .A2(n376), .ZN(n460) );
  NAND2_X1 U568 ( .A1(n459), .A2(n375), .ZN(n466) );
  NAND2_X1 U569 ( .A1(n468), .A2(n470), .ZN(n469) );
  NAND2_X1 U570 ( .A1(n604), .A2(n472), .ZN(n468) );
  NOR2_X1 U571 ( .A1(n604), .A2(n476), .ZN(n473) );
  XOR2_X1 U572 ( .A(n553), .B(n552), .Z(n477) );
  NAND2_X1 U573 ( .A1(n729), .A2(KEYINPUT47), .ZN(n633) );
  XNOR2_X2 U574 ( .A(G119), .B(KEYINPUT3), .ZN(n478) );
  XNOR2_X2 U575 ( .A(n478), .B(G116), .ZN(n537) );
  XNOR2_X1 U576 ( .A(G113), .B(G122), .ZN(n480) );
  XNOR2_X1 U577 ( .A(n480), .B(n479), .ZN(n520) );
  INV_X1 U578 ( .A(n520), .ZN(n481) );
  XNOR2_X2 U579 ( .A(n506), .B(KEYINPUT4), .ZN(n536) );
  XNOR2_X1 U580 ( .A(n790), .B(KEYINPUT72), .ZN(n553) );
  XNOR2_X1 U581 ( .A(G146), .B(G125), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n519), .B(n484), .ZN(n487) );
  NAND2_X1 U583 ( .A1(n808), .A2(G224), .ZN(n485) );
  XNOR2_X1 U584 ( .A(n485), .B(KEYINPUT94), .ZN(n486) );
  XNOR2_X1 U585 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U586 ( .A(n553), .B(n488), .ZN(n489) );
  NAND2_X1 U587 ( .A1(n491), .A2(n570), .ZN(n493) );
  NAND2_X1 U588 ( .A1(n493), .A2(G210), .ZN(n492) );
  AND2_X1 U589 ( .A1(n493), .A2(G214), .ZN(n648) );
  XNOR2_X1 U590 ( .A(n494), .B(KEYINPUT14), .ZN(n779) );
  INV_X1 U591 ( .A(G952), .ZN(n678) );
  NAND2_X1 U592 ( .A1(n808), .A2(n678), .ZN(n496) );
  OR2_X1 U593 ( .A1(n808), .A2(G902), .ZN(n495) );
  AND2_X1 U594 ( .A1(n496), .A2(n495), .ZN(n497) );
  AND2_X1 U595 ( .A1(n779), .A2(n497), .ZN(n610) );
  INV_X1 U596 ( .A(KEYINPUT95), .ZN(n498) );
  XNOR2_X1 U597 ( .A(n498), .B(G898), .ZN(n792) );
  NAND2_X1 U598 ( .A1(n792), .A2(G953), .ZN(n499) );
  INV_X1 U599 ( .A(KEYINPUT69), .ZN(n500) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n503) );
  NAND2_X1 U601 ( .A1(G234), .A2(n808), .ZN(n501) );
  XOR2_X1 U602 ( .A(KEYINPUT8), .B(n501), .Z(n559) );
  NAND2_X1 U603 ( .A1(G217), .A2(n559), .ZN(n502) );
  XNOR2_X1 U604 ( .A(n503), .B(n502), .ZN(n510) );
  XNOR2_X1 U605 ( .A(n505), .B(n504), .ZN(n508) );
  INV_X1 U606 ( .A(n506), .ZN(n507) );
  XNOR2_X1 U607 ( .A(n508), .B(n507), .ZN(n509) );
  NAND2_X1 U608 ( .A1(n698), .A2(n570), .ZN(n512) );
  XNOR2_X1 U609 ( .A(KEYINPUT98), .B(G478), .ZN(n511) );
  XNOR2_X1 U610 ( .A(n512), .B(n511), .ZN(n602) );
  INV_X1 U611 ( .A(n602), .ZN(n525) );
  XOR2_X1 U612 ( .A(KEYINPUT97), .B(G140), .Z(n514) );
  XNOR2_X1 U613 ( .A(G143), .B(G131), .ZN(n513) );
  XNOR2_X1 U614 ( .A(n514), .B(n513), .ZN(n518) );
  XOR2_X1 U615 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n516) );
  NAND2_X1 U616 ( .A1(n538), .A2(G214), .ZN(n515) );
  XNOR2_X1 U617 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U618 ( .A(n518), .B(n517), .ZN(n522) );
  XNOR2_X1 U619 ( .A(n519), .B(KEYINPUT10), .ZN(n568) );
  XNOR2_X1 U620 ( .A(n568), .B(n520), .ZN(n521) );
  XNOR2_X1 U621 ( .A(n522), .B(n521), .ZN(n675) );
  NAND2_X1 U622 ( .A1(n675), .A2(n570), .ZN(n524) );
  XNOR2_X1 U623 ( .A(KEYINPUT13), .B(G475), .ZN(n523) );
  XNOR2_X1 U624 ( .A(n524), .B(n523), .ZN(n601) );
  NAND2_X1 U625 ( .A1(n525), .A2(n601), .ZN(n770) );
  NAND2_X1 U626 ( .A1(G234), .A2(n669), .ZN(n526) );
  XNOR2_X1 U627 ( .A(KEYINPUT20), .B(n526), .ZN(n571) );
  NAND2_X1 U628 ( .A1(n571), .A2(G221), .ZN(n528) );
  INV_X1 U629 ( .A(KEYINPUT21), .ZN(n527) );
  XNOR2_X1 U630 ( .A(n528), .B(n527), .ZN(n754) );
  INV_X1 U631 ( .A(n754), .ZN(n529) );
  OR2_X1 U632 ( .A1(n770), .A2(n529), .ZN(n530) );
  XNOR2_X1 U633 ( .A(n530), .B(KEYINPUT101), .ZN(n531) );
  NAND2_X1 U634 ( .A1(n583), .A2(n531), .ZN(n534) );
  XNOR2_X1 U635 ( .A(KEYINPUT76), .B(KEYINPUT22), .ZN(n532) );
  NAND2_X1 U636 ( .A1(n538), .A2(G210), .ZN(n540) );
  XNOR2_X1 U637 ( .A(n540), .B(n539), .ZN(n542) );
  XNOR2_X1 U638 ( .A(G137), .B(KEYINPUT5), .ZN(n541) );
  XNOR2_X1 U639 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U640 ( .A(n537), .B(n543), .ZN(n544) );
  XNOR2_X1 U641 ( .A(n554), .B(n544), .ZN(n688) );
  XNOR2_X1 U642 ( .A(G472), .B(KEYINPUT75), .ZN(n545) );
  XNOR2_X2 U643 ( .A(n546), .B(n545), .ZN(n757) );
  INV_X1 U644 ( .A(KEYINPUT100), .ZN(n547) );
  XNOR2_X1 U645 ( .A(n547), .B(KEYINPUT6), .ZN(n548) );
  NAND2_X1 U646 ( .A1(n808), .A2(G227), .ZN(n549) );
  XNOR2_X1 U647 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U648 ( .A(n551), .B(n566), .ZN(n552) );
  XNOR2_X1 U649 ( .A(KEYINPUT71), .B(G469), .ZN(n555) );
  XNOR2_X1 U650 ( .A(KEYINPUT68), .B(KEYINPUT1), .ZN(n558) );
  BUF_X1 U651 ( .A(n584), .Z(n751) );
  XNOR2_X1 U652 ( .A(n751), .B(KEYINPUT93), .ZN(n643) );
  NAND2_X1 U653 ( .A1(G221), .A2(n559), .ZN(n565) );
  XOR2_X1 U654 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n561) );
  XNOR2_X1 U655 ( .A(G128), .B(G110), .ZN(n560) );
  XNOR2_X1 U656 ( .A(n561), .B(n560), .ZN(n563) );
  INV_X1 U657 ( .A(n566), .ZN(n567) );
  XNOR2_X1 U658 ( .A(n568), .B(n567), .ZN(n799) );
  XNOR2_X1 U659 ( .A(n569), .B(n799), .ZN(n693) );
  NAND2_X1 U660 ( .A1(n693), .A2(n570), .ZN(n575) );
  NAND2_X1 U661 ( .A1(n571), .A2(G217), .ZN(n573) );
  INV_X1 U662 ( .A(KEYINPUT25), .ZN(n572) );
  XNOR2_X1 U663 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X2 U664 ( .A(n575), .B(n574), .ZN(n626) );
  INV_X1 U665 ( .A(n626), .ZN(n580) );
  AND2_X1 U666 ( .A1(n643), .A2(n580), .ZN(n576) );
  AND2_X1 U667 ( .A1(n354), .A2(n576), .ZN(n577) );
  INV_X1 U668 ( .A(n757), .ZN(n578) );
  NOR2_X1 U669 ( .A1(n411), .A2(n578), .ZN(n579) );
  OR2_X1 U670 ( .A1(KEYINPUT44), .A2(KEYINPUT91), .ZN(n581) );
  INV_X1 U671 ( .A(n601), .ZN(n586) );
  NAND2_X1 U672 ( .A1(n586), .A2(n602), .ZN(n619) );
  XNOR2_X1 U673 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n587) );
  XNOR2_X2 U674 ( .A(n588), .B(n587), .ZN(n683) );
  NAND2_X1 U675 ( .A1(n683), .A2(KEYINPUT90), .ZN(n590) );
  AND2_X1 U676 ( .A1(n590), .A2(KEYINPUT44), .ZN(n591) );
  INV_X1 U677 ( .A(KEYINPUT44), .ZN(n592) );
  NAND2_X1 U678 ( .A1(n592), .A2(KEYINPUT90), .ZN(n593) );
  INV_X1 U679 ( .A(n583), .ZN(n598) );
  OR2_X1 U680 ( .A1(n757), .A2(n750), .ZN(n594) );
  OR2_X1 U681 ( .A1(n751), .A2(n594), .ZN(n760) );
  INV_X1 U682 ( .A(KEYINPUT96), .ZN(n596) );
  NAND2_X1 U683 ( .A1(n602), .A2(n601), .ZN(n600) );
  INV_X1 U684 ( .A(KEYINPUT99), .ZN(n599) );
  XNOR2_X1 U685 ( .A(n600), .B(n599), .ZN(n735) );
  OR2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n732) );
  AND2_X1 U687 ( .A1(n735), .A2(n732), .ZN(n767) );
  NOR2_X1 U688 ( .A1(n603), .A2(n767), .ZN(n608) );
  BUF_X1 U689 ( .A(n604), .Z(n605) );
  NAND2_X1 U690 ( .A1(n605), .A2(n354), .ZN(n607) );
  NAND2_X1 U691 ( .A1(n751), .A2(n626), .ZN(n606) );
  NAND2_X1 U692 ( .A1(G953), .A2(G900), .ZN(n609) );
  NAND2_X1 U693 ( .A1(n610), .A2(n609), .ZN(n625) );
  INV_X1 U694 ( .A(n625), .ZN(n611) );
  OR2_X1 U695 ( .A1(n757), .A2(n648), .ZN(n615) );
  INV_X1 U696 ( .A(KEYINPUT104), .ZN(n613) );
  XNOR2_X1 U697 ( .A(n613), .B(KEYINPUT30), .ZN(n614) );
  XNOR2_X1 U698 ( .A(n615), .B(n614), .ZN(n616) );
  INV_X1 U699 ( .A(KEYINPUT105), .ZN(n621) );
  BUF_X1 U700 ( .A(n623), .Z(n624) );
  INV_X1 U701 ( .A(n624), .ZN(n631) );
  XNOR2_X1 U702 ( .A(KEYINPUT28), .B(KEYINPUT106), .ZN(n628) );
  INV_X1 U703 ( .A(n650), .ZN(n630) );
  INV_X1 U704 ( .A(KEYINPUT83), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n767), .A2(KEYINPUT47), .ZN(n634) );
  BUF_X1 U706 ( .A(n636), .Z(n638) );
  NOR2_X1 U707 ( .A1(n732), .A2(n637), .ZN(n657) );
  NAND2_X1 U708 ( .A1(n638), .A2(n657), .ZN(n639) );
  OR2_X1 U709 ( .A1(n354), .A2(n639), .ZN(n641) );
  INV_X1 U710 ( .A(KEYINPUT36), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U712 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U713 ( .A(n644), .B(KEYINPUT108), .ZN(n812) );
  INV_X1 U714 ( .A(n618), .ZN(n663) );
  INV_X1 U715 ( .A(KEYINPUT73), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n645), .B(KEYINPUT39), .ZN(n646) );
  INV_X1 U717 ( .A(n732), .ZN(n730) );
  NAND2_X1 U718 ( .A1(n363), .A2(n450), .ZN(n766) );
  NOR2_X1 U719 ( .A1(n766), .A2(n770), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n649), .B(KEYINPUT41), .ZN(n764) );
  NOR2_X1 U721 ( .A1(n764), .A2(n650), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n651), .B(KEYINPUT42), .ZN(n814) );
  INV_X1 U723 ( .A(n814), .ZN(n652) );
  INV_X1 U724 ( .A(KEYINPUT46), .ZN(n653) );
  INV_X1 U725 ( .A(KEYINPUT48), .ZN(n654) );
  INV_X1 U726 ( .A(n735), .ZN(n655) );
  NAND2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n681) );
  AND2_X1 U728 ( .A1(n657), .A2(n450), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n751), .A2(n658), .ZN(n660) );
  OR2_X1 U730 ( .A1(n660), .A2(n354), .ZN(n662) );
  XNOR2_X1 U731 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n661) );
  XNOR2_X1 U732 ( .A(n662), .B(n661), .ZN(n664) );
  OR2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n680) );
  AND2_X1 U734 ( .A1(n681), .A2(n680), .ZN(n665) );
  INV_X1 U735 ( .A(KEYINPUT2), .ZN(n667) );
  NOR2_X1 U736 ( .A1(n667), .A2(KEYINPUT86), .ZN(n668) );
  INV_X1 U737 ( .A(n801), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n378), .A2(G475), .ZN(n677) );
  XNOR2_X1 U739 ( .A(n677), .B(n676), .ZN(n679) );
  XNOR2_X1 U740 ( .A(n680), .B(G140), .ZN(G42) );
  XNOR2_X1 U741 ( .A(n681), .B(G134), .ZN(G36) );
  XOR2_X1 U742 ( .A(G101), .B(n682), .Z(G3) );
  XOR2_X1 U743 ( .A(n683), .B(G122), .Z(G24) );
  BUF_X1 U744 ( .A(n684), .Z(n685) );
  XOR2_X1 U745 ( .A(n685), .B(G110), .Z(G12) );
  XOR2_X1 U746 ( .A(n686), .B(G119), .Z(G21) );
  XNOR2_X1 U747 ( .A(n687), .B(G143), .ZN(G45) );
  NAND2_X1 U748 ( .A1(n379), .A2(G472), .ZN(n690) );
  XNOR2_X1 U749 ( .A(n690), .B(n689), .ZN(n691) );
  NAND2_X1 U750 ( .A1(n691), .A2(n714), .ZN(n692) );
  XNOR2_X1 U751 ( .A(n692), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U752 ( .A1(n379), .A2(G217), .ZN(n695) );
  XNOR2_X1 U753 ( .A(n693), .B(KEYINPUT120), .ZN(n694) );
  XNOR2_X1 U754 ( .A(n695), .B(n694), .ZN(n696) );
  NAND2_X1 U755 ( .A1(n696), .A2(n714), .ZN(n697) );
  XNOR2_X1 U756 ( .A(n697), .B(KEYINPUT121), .ZN(G66) );
  NAND2_X1 U757 ( .A1(n378), .A2(G478), .ZN(n699) );
  XNOR2_X1 U758 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X1 U759 ( .A1(n700), .A2(n714), .ZN(n701) );
  XNOR2_X1 U760 ( .A(n701), .B(KEYINPUT119), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n358), .A2(G469), .ZN(n706) );
  XOR2_X1 U762 ( .A(KEYINPUT118), .B(KEYINPUT57), .Z(n703) );
  XNOR2_X1 U763 ( .A(n703), .B(KEYINPUT58), .ZN(n704) );
  XNOR2_X1 U764 ( .A(n702), .B(n704), .ZN(n705) );
  XNOR2_X1 U765 ( .A(n706), .B(n705), .ZN(n708) );
  INV_X1 U766 ( .A(n714), .ZN(n707) );
  NOR2_X1 U767 ( .A1(n708), .A2(n707), .ZN(G54) );
  NAND2_X1 U768 ( .A1(n379), .A2(G210), .ZN(n713) );
  BUF_X1 U769 ( .A(n709), .Z(n711) );
  XNOR2_X1 U770 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n710) );
  XNOR2_X1 U771 ( .A(n713), .B(n712), .ZN(n715) );
  NAND2_X1 U772 ( .A1(n715), .A2(n714), .ZN(n717) );
  XNOR2_X1 U773 ( .A(KEYINPUT89), .B(KEYINPUT56), .ZN(n716) );
  XNOR2_X1 U774 ( .A(n717), .B(n716), .ZN(G51) );
  NOR2_X1 U775 ( .A1(n369), .A2(n732), .ZN(n718) );
  XOR2_X1 U776 ( .A(G104), .B(n718), .Z(G6) );
  XOR2_X1 U777 ( .A(KEYINPUT111), .B(KEYINPUT27), .Z(n720) );
  XNOR2_X1 U778 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n719) );
  XNOR2_X1 U779 ( .A(n720), .B(n719), .ZN(n724) );
  NOR2_X1 U780 ( .A1(n369), .A2(n735), .ZN(n722) );
  XNOR2_X1 U781 ( .A(G107), .B(KEYINPUT26), .ZN(n721) );
  XNOR2_X1 U782 ( .A(n722), .B(n721), .ZN(n723) );
  XOR2_X1 U783 ( .A(n724), .B(n723), .Z(G9) );
  NOR2_X1 U784 ( .A1(n729), .A2(n735), .ZN(n728) );
  XOR2_X1 U785 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n726) );
  XNOR2_X1 U786 ( .A(G128), .B(KEYINPUT113), .ZN(n725) );
  XNOR2_X1 U787 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U788 ( .A(n728), .B(n727), .ZN(G30) );
  NAND2_X1 U789 ( .A1(n407), .A2(n730), .ZN(n731) );
  XNOR2_X1 U790 ( .A(n731), .B(G146), .ZN(G48) );
  NOR2_X1 U791 ( .A1(n732), .A2(n734), .ZN(n733) );
  XOR2_X1 U792 ( .A(G113), .B(n733), .Z(G15) );
  NOR2_X1 U793 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U794 ( .A(G116), .B(n736), .Z(G18) );
  XOR2_X1 U795 ( .A(KEYINPUT81), .B(KEYINPUT2), .Z(n742) );
  NOR2_X1 U796 ( .A1(n801), .A2(n742), .ZN(n738) );
  INV_X1 U797 ( .A(KEYINPUT85), .ZN(n737) );
  NOR2_X1 U798 ( .A1(n738), .A2(n737), .ZN(n739) );
  INV_X1 U799 ( .A(n671), .ZN(n741) );
  NOR2_X1 U800 ( .A1(n801), .A2(KEYINPUT85), .ZN(n740) );
  NOR2_X1 U801 ( .A1(n741), .A2(n740), .ZN(n743) );
  OR2_X1 U802 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U803 ( .A1(n745), .A2(n744), .ZN(n749) );
  INV_X1 U804 ( .A(n746), .ZN(n774) );
  NOR2_X1 U805 ( .A1(n764), .A2(n774), .ZN(n747) );
  NOR2_X1 U806 ( .A1(n747), .A2(G953), .ZN(n748) );
  NAND2_X1 U807 ( .A1(n749), .A2(n748), .ZN(n783) );
  NAND2_X1 U808 ( .A1(n751), .A2(n750), .ZN(n753) );
  XNOR2_X1 U809 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n752) );
  XNOR2_X1 U810 ( .A(n753), .B(n752), .ZN(n759) );
  NOR2_X1 U811 ( .A1(n754), .A2(n626), .ZN(n755) );
  XNOR2_X1 U812 ( .A(KEYINPUT49), .B(n755), .ZN(n756) );
  AND2_X1 U813 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U814 ( .A1(n759), .A2(n758), .ZN(n761) );
  NAND2_X1 U815 ( .A1(n761), .A2(n760), .ZN(n763) );
  XOR2_X1 U816 ( .A(KEYINPUT51), .B(KEYINPUT115), .Z(n762) );
  XNOR2_X1 U817 ( .A(n763), .B(n762), .ZN(n765) );
  NOR2_X1 U818 ( .A1(n765), .A2(n764), .ZN(n777) );
  NOR2_X1 U819 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U820 ( .A(KEYINPUT117), .B(n768), .Z(n773) );
  NOR2_X1 U821 ( .A1(n363), .A2(n450), .ZN(n769) );
  NOR2_X1 U822 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U823 ( .A(KEYINPUT116), .B(n771), .ZN(n772) );
  NOR2_X1 U824 ( .A1(n773), .A2(n772), .ZN(n775) );
  NOR2_X1 U825 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U826 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U827 ( .A(KEYINPUT52), .B(n778), .ZN(n781) );
  NAND2_X1 U828 ( .A1(n779), .A2(G952), .ZN(n780) );
  NOR2_X1 U829 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U830 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U831 ( .A(KEYINPUT53), .B(n784), .ZN(G75) );
  NAND2_X1 U832 ( .A1(n671), .A2(n808), .ZN(n788) );
  NAND2_X1 U833 ( .A1(G953), .A2(G224), .ZN(n785) );
  XNOR2_X1 U834 ( .A(KEYINPUT61), .B(n785), .ZN(n786) );
  NAND2_X1 U835 ( .A1(n786), .A2(n792), .ZN(n787) );
  NAND2_X1 U836 ( .A1(n788), .A2(n787), .ZN(n796) );
  XOR2_X1 U837 ( .A(KEYINPUT123), .B(n790), .Z(n791) );
  XNOR2_X1 U838 ( .A(n789), .B(n791), .ZN(n794) );
  NOR2_X1 U839 ( .A1(n792), .A2(n808), .ZN(n793) );
  NOR2_X1 U840 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U841 ( .A(n796), .B(n795), .ZN(n797) );
  XNOR2_X1 U842 ( .A(KEYINPUT122), .B(n797), .ZN(G69) );
  XNOR2_X1 U843 ( .A(n799), .B(KEYINPUT124), .ZN(n800) );
  XNOR2_X1 U844 ( .A(n798), .B(n800), .ZN(n804) );
  XNOR2_X1 U845 ( .A(n801), .B(n804), .ZN(n802) );
  NOR2_X1 U846 ( .A1(n802), .A2(G953), .ZN(n803) );
  XNOR2_X1 U847 ( .A(KEYINPUT125), .B(n803), .ZN(n811) );
  XNOR2_X1 U848 ( .A(G227), .B(n804), .ZN(n805) );
  NAND2_X1 U849 ( .A1(n805), .A2(G900), .ZN(n806) );
  XOR2_X1 U850 ( .A(KEYINPUT126), .B(n806), .Z(n807) );
  NOR2_X1 U851 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U852 ( .A(KEYINPUT127), .B(n809), .ZN(n810) );
  NAND2_X1 U853 ( .A1(n811), .A2(n810), .ZN(G72) );
  XOR2_X1 U854 ( .A(G125), .B(n812), .Z(n813) );
  XNOR2_X1 U855 ( .A(KEYINPUT37), .B(n813), .ZN(G27) );
  XOR2_X1 U856 ( .A(G137), .B(n814), .Z(G39) );
endmodule

