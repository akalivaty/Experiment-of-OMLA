//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(KEYINPUT90), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(KEYINPUT90), .ZN(new_n204));
  NOR2_X1   g003(.A1(KEYINPUT91), .A2(G36gat), .ZN(new_n205));
  AND2_X1   g004(.A1(KEYINPUT91), .A2(G36gat), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n203), .A2(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n202), .A2(new_n208), .A3(KEYINPUT14), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G50gat), .ZN(new_n214));
  INV_X1    g013(.A(G50gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G43gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT15), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n207), .A2(new_n212), .A3(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(KEYINPUT92), .A2(G50gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(KEYINPUT92), .A2(G50gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n213), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT93), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n223), .B(new_n213), .C1(new_n219), .C2(new_n220), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n216), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n218), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n217), .B1(new_n207), .B2(new_n212), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT94), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT94), .ZN(new_n230));
  INV_X1    g029(.A(new_n228), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n221), .A2(KEYINPUT93), .B1(G43gat), .B2(new_n215), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT15), .B1(new_n232), .B2(new_n224), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n230), .B(new_n231), .C1(new_n233), .C2(new_n218), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G1gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT16), .ZN(new_n237));
  INV_X1    g036(.A(G15gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G22gat), .ZN(new_n239));
  INV_X1    g038(.A(G22gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G15gat), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n237), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(G1gat), .B1(new_n239), .B2(new_n241), .ZN(new_n243));
  OAI21_X1  g042(.A(G8gat), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n237), .A2(new_n239), .A3(new_n241), .ZN(new_n245));
  INV_X1    g044(.A(G8gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(G15gat), .B(G22gat), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n245), .B(new_n246), .C1(G1gat), .C2(new_n247), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n244), .A2(new_n248), .A3(KEYINPUT95), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT95), .B1(new_n244), .B2(new_n248), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G229gat), .A2(G233gat), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT17), .B1(new_n229), .B2(new_n234), .ZN(new_n255));
  OAI211_X1 g054(.A(KEYINPUT17), .B(new_n231), .C1(new_n233), .C2(new_n218), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(new_n244), .A3(new_n248), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n253), .B(new_n254), .C1(new_n255), .C2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT18), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT96), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n251), .B1(new_n229), .B2(new_n234), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT17), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n235), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n257), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT96), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT18), .A4(new_n254), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n254), .B(KEYINPUT13), .Z(new_n269));
  AND3_X1   g068(.A1(new_n229), .A2(new_n251), .A3(new_n234), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n269), .B1(new_n270), .B2(new_n261), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT97), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(KEYINPUT97), .B(new_n269), .C1(new_n270), .C2(new_n261), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n273), .A2(new_n274), .B1(new_n259), .B2(new_n258), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G113gat), .B(G141gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT89), .B(G197gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(KEYINPUT11), .B(G169gat), .Z(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT12), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n276), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n275), .A3(new_n282), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G113gat), .B(G120gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n291));
  INV_X1    g090(.A(G113gat), .ZN(new_n292));
  INV_X1    g091(.A(G120gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G113gat), .A2(G120gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT70), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n290), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(KEYINPUT68), .B(G127gat), .Z(new_n298));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(G134gat), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G127gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT68), .B(G127gat), .ZN(new_n303));
  OAI211_X1 g102(.A(KEYINPUT69), .B(new_n302), .C1(new_n303), .C2(new_n301), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n297), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n291), .ZN(new_n306));
  INV_X1    g105(.A(G127gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(G134gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(new_n294), .A3(new_n295), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G141gat), .B(G148gat), .Z(new_n311));
  INV_X1    g110(.A(KEYINPUT2), .ZN(new_n312));
  INV_X1    g111(.A(G155gat), .ZN(new_n313));
  INV_X1    g112(.A(G162gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G141gat), .B(G148gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n321), .A2(new_n312), .B1(G155gat), .B2(G162gat), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n316), .A2(KEYINPUT75), .ZN(new_n324));
  INV_X1    g123(.A(new_n316), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT75), .B1(new_n313), .B2(new_n314), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n318), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT3), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n330), .B(new_n318), .C1(new_n323), .C2(new_n327), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n310), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  MUX2_X1   g131(.A(KEYINPUT75), .B(new_n326), .S(new_n316), .Z(new_n333));
  NAND2_X1  g132(.A1(new_n322), .A2(new_n320), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n311), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n333), .A2(new_n335), .B1(new_n317), .B2(new_n311), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(new_n305), .A3(new_n309), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n332), .A2(KEYINPUT4), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341));
  AND4_X1   g140(.A1(new_n341), .A2(new_n336), .A3(new_n305), .A4(new_n309), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AND4_X1   g142(.A1(KEYINPUT84), .A2(new_n338), .A3(new_n340), .A4(new_n343), .ZN(new_n344));
  AOI211_X1 g143(.A(new_n306), .B(new_n288), .C1(new_n307), .C2(G134gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n346), .B1(new_n298), .B2(G134gat), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n303), .A2(KEYINPUT69), .A3(new_n301), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n345), .B1(new_n349), .B2(new_n297), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n341), .B1(new_n350), .B2(new_n336), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n342), .B1(new_n351), .B2(new_n332), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT84), .B1(new_n352), .B2(new_n340), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n344), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n310), .A2(new_n328), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n337), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n354), .B(KEYINPUT39), .C1(new_n340), .C2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n343), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(new_n339), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(KEYINPUT84), .A3(new_n340), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT39), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n363));
  XOR2_X1   g162(.A(G1gat), .B(G29gat), .Z(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G57gat), .B(G85gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n362), .A2(new_n363), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT39), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n344), .B2(new_n353), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT85), .B1(new_n372), .B2(new_n368), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n357), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT40), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n357), .B(KEYINPUT40), .C1(new_n370), .C2(new_n373), .ZN(new_n377));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(KEYINPUT74), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  XNOR2_X1  g180(.A(G197gat), .B(G204gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n383));
  INV_X1    g182(.A(G211gat), .ZN(new_n384));
  INV_X1    g183(.A(G218gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G211gat), .B(G218gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n382), .A3(new_n386), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394));
  INV_X1    g193(.A(G183gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT27), .ZN(new_n396));
  AOI21_X1  g195(.A(G190gat), .B1(new_n396), .B2(KEYINPUT66), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT27), .B(G183gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n397), .B1(KEYINPUT66), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G190gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(KEYINPUT28), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n405), .B(KEYINPUT67), .Z(new_n406));
  NAND2_X1  g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT26), .ZN(new_n409));
  NOR2_X1   g208(.A1(G169gat), .A2(G176gat), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n406), .A2(new_n411), .B1(G183gat), .B2(G190gat), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G183gat), .A2(G190gat), .ZN(new_n414));
  OAI221_X1 g213(.A(new_n407), .B1(new_n414), .B2(KEYINPUT24), .C1(new_n410), .C2(KEYINPUT23), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n402), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n416), .A2(KEYINPUT24), .A3(new_n414), .ZN(new_n417));
  INV_X1    g216(.A(new_n410), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT23), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT25), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n415), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n415), .A2(new_n417), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT65), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT64), .B(G176gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n419), .A2(G169gat), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n423), .A3(new_n425), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT25), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n421), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n394), .B1(new_n413), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G226gat), .A2(G233gat), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT73), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(new_n430), .ZN(new_n435));
  INV_X1    g234(.A(new_n421), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n435), .A2(new_n436), .B1(new_n404), .B2(new_n412), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n434), .B1(new_n437), .B2(new_n433), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n404), .A2(new_n412), .ZN(new_n439));
  INV_X1    g238(.A(new_n428), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(new_n426), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT25), .B1(new_n441), .B2(new_n422), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n439), .B1(new_n442), .B2(new_n421), .ZN(new_n443));
  INV_X1    g242(.A(new_n433), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(KEYINPUT73), .A3(new_n444), .ZN(new_n445));
  AOI221_X4 g244(.A(new_n393), .B1(new_n432), .B2(new_n433), .C1(new_n438), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n432), .A2(new_n433), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n444), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n392), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n381), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n438), .A2(new_n445), .B1(new_n433), .B2(new_n432), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n392), .ZN(new_n452));
  INV_X1    g251(.A(new_n449), .ZN(new_n453));
  INV_X1    g252(.A(new_n381), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n455), .A3(KEYINPUT30), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n446), .A2(new_n449), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT30), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n454), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT77), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n356), .B2(new_n340), .ZN(new_n461));
  AOI211_X1 g260(.A(KEYINPUT77), .B(new_n339), .C1(new_n355), .C2(new_n337), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n359), .A2(new_n339), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n464), .A2(new_n466), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n369), .A3(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n456), .A2(new_n459), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n376), .A2(new_n377), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT86), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G78gat), .B(G106gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(KEYINPUT31), .B(G50gat), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n475), .B(new_n476), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT29), .B1(new_n390), .B2(new_n391), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n328), .B1(new_n479), .B2(KEYINPUT3), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n331), .A2(new_n394), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(new_n392), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT80), .B1(new_n481), .B2(new_n392), .ZN(new_n483));
  NAND2_X1  g282(.A1(G228gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  OAI221_X1 g285(.A(new_n480), .B1(KEYINPUT80), .B2(new_n484), .C1(new_n481), .C2(new_n392), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(G22gat), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(G22gat), .B1(new_n486), .B2(new_n487), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n478), .B(new_n488), .C1(new_n489), .C2(KEYINPUT82), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT83), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT83), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n488), .A2(new_n478), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n486), .A2(new_n487), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n240), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n488), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT81), .B1(new_n501), .B2(new_n477), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT81), .ZN(new_n503));
  AOI211_X1 g302(.A(new_n503), .B(new_n478), .C1(new_n500), .C2(new_n488), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n466), .B1(new_n463), .B2(new_n464), .ZN(new_n507));
  INV_X1    g306(.A(new_n469), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n368), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n470), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n468), .A2(KEYINPUT6), .A3(new_n369), .A4(new_n469), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n511), .A2(new_n512), .A3(new_n455), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT88), .B(KEYINPUT37), .ZN(new_n514));
  AOI211_X1 g313(.A(KEYINPUT38), .B(new_n454), .C1(new_n457), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n451), .A2(new_n393), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n447), .A2(new_n448), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n392), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT87), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT87), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n452), .A2(new_n453), .A3(new_n514), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n525), .B(new_n381), .C1(new_n457), .C2(new_n517), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n515), .A2(new_n524), .B1(new_n526), .B2(KEYINPUT38), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n506), .B1(new_n513), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n376), .A2(new_n471), .A3(KEYINPUT86), .A4(new_n377), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n474), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n511), .ZN(new_n531));
  INV_X1    g330(.A(new_n512), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n456), .A2(new_n459), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n506), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(G227gat), .A2(G233gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n350), .B1(new_n413), .B2(new_n431), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n439), .B(new_n310), .C1(new_n442), .C2(new_n421), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n537), .A3(new_n539), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT33), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G43gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(G71gat), .B(G99gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n542), .B(KEYINPUT32), .C1(new_n543), .C2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n542), .B2(KEYINPUT32), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n542), .A2(new_n543), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n549), .B1(new_n548), .B2(new_n550), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT34), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT34), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n542), .A2(KEYINPUT32), .ZN(new_n556));
  INV_X1    g355(.A(new_n546), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n550), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT71), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n555), .B1(new_n561), .B2(new_n547), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n541), .B1(new_n554), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n553), .A2(KEYINPUT34), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n561), .A2(new_n555), .A3(new_n547), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n567), .A3(new_n540), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n563), .A2(new_n564), .A3(new_n565), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n565), .ZN(new_n570));
  NAND2_X1  g369(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n566), .A2(new_n567), .A3(new_n540), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n540), .B1(new_n566), .B2(new_n567), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n530), .A2(new_n536), .A3(new_n569), .A4(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n572), .A2(new_n573), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT35), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n498), .A2(new_n505), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n511), .A2(new_n512), .B1(new_n456), .B2(new_n459), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n563), .A2(new_n578), .A3(new_n579), .A4(new_n568), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n287), .B1(new_n575), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(new_n313), .ZN(new_n586));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT98), .B1(new_n590), .B2(KEYINPUT9), .ZN(new_n591));
  XNOR2_X1  g390(.A(G71gat), .B(G78gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G57gat), .B(G64gat), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n591), .B(new_n592), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT98), .ZN(new_n596));
  NOR2_X1   g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  OAI22_X1  g396(.A1(new_n594), .A2(new_n596), .B1(new_n590), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G57gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G64gat), .ZN(new_n600));
  INV_X1    g399(.A(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G57gat), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n594), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(G127gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(G127gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT21), .ZN(new_n612));
  INV_X1    g411(.A(new_n605), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n251), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n611), .A2(new_n615), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n589), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(new_n616), .A3(new_n588), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n623));
  NAND2_X1  g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT8), .ZN(new_n625));
  NAND2_X1  g424(.A1(G85gat), .A2(G92gat), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT7), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G85gat), .ZN(new_n629));
  INV_X1    g428(.A(G92gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n625), .A2(new_n628), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G99gat), .B(G106gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g435(.A1(KEYINPUT8), .A2(new_n624), .B1(new_n629), .B2(new_n630), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n637), .A2(new_n634), .A3(new_n628), .A4(new_n632), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(KEYINPUT99), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n633), .A2(new_n640), .A3(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT100), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n644), .A3(new_n641), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT92), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n215), .ZN(new_n648));
  NAND2_X1  g447(.A1(KEYINPUT92), .A2(G50gat), .ZN(new_n649));
  AOI21_X1  g448(.A(G43gat), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n216), .B1(new_n650), .B2(new_n223), .ZN(new_n651));
  INV_X1    g450(.A(new_n224), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n226), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n218), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n230), .B1(new_n655), .B2(new_n231), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n227), .A2(KEYINPUT94), .A3(new_n228), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n646), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(G232gat), .A2(G233gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT41), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n256), .A3(new_n645), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n658), .B(new_n660), .C1(new_n255), .C2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G190gat), .B(G218gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n623), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n659), .A2(KEYINPUT41), .ZN(new_n665));
  XNOR2_X1  g464(.A(G134gat), .B(G162gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n235), .A2(new_n646), .B1(KEYINPUT41), .B2(new_n659), .ZN(new_n668));
  INV_X1    g467(.A(new_n663), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n668), .B(new_n669), .C1(new_n255), .C2(new_n661), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n658), .A2(new_n660), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n255), .A2(new_n661), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n663), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n664), .A2(new_n667), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n673), .A2(new_n670), .A3(KEYINPUT101), .A4(new_n667), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n605), .A2(KEYINPUT10), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n639), .A2(new_n644), .A3(new_n641), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n644), .B1(new_n639), .B2(new_n641), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT10), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n605), .B1(new_n639), .B2(new_n641), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n636), .A2(new_n638), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n605), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n683), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(G230gat), .A2(G233gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR3_X1    g489(.A1(new_n684), .A2(new_n686), .A3(new_n689), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(G120gat), .B(G148gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(G176gat), .B(G204gat), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n693), .B(new_n694), .Z(new_n695));
  OR2_X1    g494(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n690), .A2(new_n691), .A3(new_n695), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n622), .A2(new_n677), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n584), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n533), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(new_n236), .ZN(G1324gat));
  INV_X1    g504(.A(new_n702), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT102), .B(KEYINPUT16), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(new_n246), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n706), .A2(new_n535), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n246), .B1(new_n706), .B2(new_n535), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT42), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(KEYINPUT42), .B2(new_n709), .ZN(G1325gat));
  NAND2_X1  g511(.A1(new_n574), .A2(new_n569), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT104), .B1(new_n574), .B2(new_n569), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n706), .A2(G15gat), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n584), .A2(new_n576), .A3(new_n701), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n719), .A2(KEYINPUT103), .A3(new_n238), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT103), .B1(new_n719), .B2(new_n238), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1326gat));
  OR3_X1    g523(.A1(new_n702), .A2(KEYINPUT106), .A3(new_n578), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT106), .B1(new_n702), .B2(new_n578), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT43), .B(G22gat), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n727), .B(new_n728), .Z(G1327gat));
  XNOR2_X1  g528(.A(new_n622), .B(KEYINPUT108), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n731), .A2(new_n287), .A3(new_n698), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n474), .A2(new_n529), .A3(new_n528), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n574), .A2(new_n536), .A3(new_n569), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n583), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n677), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n674), .B2(new_n676), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n664), .A2(new_n667), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n673), .A2(new_n670), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(KEYINPUT109), .A3(new_n675), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n733), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n575), .B2(new_n583), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n732), .B1(new_n738), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(KEYINPUT110), .B(new_n732), .C1(new_n738), .C2(new_n748), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(new_n533), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n203), .B2(new_n204), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n622), .A2(new_n677), .A3(new_n698), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n584), .A2(new_n755), .ZN(new_n756));
  NOR4_X1   g555(.A1(new_n756), .A2(new_n703), .A3(new_n203), .A4(new_n204), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n754), .A2(new_n759), .ZN(G1328gat));
  INV_X1    g559(.A(new_n756), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n534), .A2(new_n205), .A3(new_n206), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT46), .Z(new_n764));
  NAND3_X1  g563(.A1(new_n751), .A2(new_n535), .A3(new_n752), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n205), .B2(new_n206), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1329gat));
  INV_X1    g566(.A(new_n576), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n756), .A2(G43gat), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n749), .B1(new_n569), .B2(new_n574), .ZN(new_n771));
  OAI211_X1 g570(.A(KEYINPUT47), .B(new_n770), .C1(new_n771), .C2(new_n213), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n751), .A2(new_n717), .A3(new_n752), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n769), .B1(new_n773), .B2(G43gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n774), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g574(.A1(new_n648), .A2(new_n649), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n756), .A2(new_n776), .A3(new_n578), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT48), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n506), .B(new_n732), .C1(new_n738), .C2(new_n748), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n751), .A2(new_n506), .A3(new_n752), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n777), .B1(new_n785), .B2(new_n776), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n786), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g586(.A(new_n622), .ZN(new_n788));
  NOR4_X1   g587(.A1(new_n286), .A2(new_n788), .A3(new_n737), .A4(new_n699), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n736), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n703), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(new_n599), .ZN(G1332gat));
  INV_X1    g591(.A(new_n790), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n534), .B(KEYINPUT112), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(G1333gat));
  INV_X1    g600(.A(new_n717), .ZN(new_n802));
  OAI21_X1  g601(.A(G71gat), .B1(new_n802), .B2(new_n790), .ZN(new_n803));
  INV_X1    g602(.A(G71gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n576), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n790), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g606(.A1(new_n790), .A2(new_n578), .ZN(new_n808));
  XOR2_X1   g607(.A(KEYINPUT114), .B(G78gat), .Z(new_n809));
  XNOR2_X1  g608(.A(new_n808), .B(new_n809), .ZN(G1335gat));
  NOR2_X1   g609(.A1(new_n286), .A2(new_n622), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n698), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n736), .A2(new_n737), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT44), .ZN(new_n814));
  INV_X1    g613(.A(new_n748), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(G85gat), .B1(new_n817), .B2(new_n703), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n677), .B1(new_n575), .B2(new_n583), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n811), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(KEYINPUT51), .A3(new_n811), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n820), .A2(KEYINPUT115), .A3(new_n821), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n698), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n533), .A2(new_n629), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n818), .B1(new_n827), .B2(new_n828), .ZN(G1336gat));
  AOI21_X1  g628(.A(new_n630), .B1(new_n816), .B2(new_n535), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n794), .A2(G92gat), .A3(new_n699), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n822), .B2(new_n824), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT52), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n794), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n630), .B1(new_n816), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n825), .A2(new_n826), .A3(new_n831), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(G1337gat));
  OAI21_X1  g638(.A(G99gat), .B1(new_n817), .B2(new_n802), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n768), .A2(G99gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n827), .B2(new_n841), .ZN(G1338gat));
  XOR2_X1   g641(.A(KEYINPUT116), .B(G106gat), .Z(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n816), .B2(new_n506), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n578), .A2(G106gat), .A3(new_n699), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n822), .B2(new_n824), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT53), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n845), .A2(KEYINPUT53), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n825), .A2(new_n826), .A3(new_n846), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(G1339gat));
  NOR2_X1   g651(.A1(new_n700), .A2(new_n286), .ZN(new_n853));
  INV_X1    g652(.A(new_n689), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n682), .A2(new_n687), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n690), .A2(KEYINPUT54), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n854), .B1(new_n682), .B2(new_n687), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n695), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n859), .A3(KEYINPUT55), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n697), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT55), .B1(new_n856), .B2(new_n859), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT117), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n856), .A2(new_n859), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n697), .A4(new_n860), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n265), .A2(new_n254), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n270), .A2(new_n261), .A3(new_n269), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n281), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n285), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n869), .A2(new_n744), .A3(new_n874), .A4(new_n740), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n285), .A2(new_n698), .A3(new_n872), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n876), .B1(new_n869), .B2(new_n286), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n877), .B2(new_n746), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n853), .B1(new_n878), .B2(new_n730), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(new_n506), .A3(new_n768), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n533), .A3(new_n794), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n287), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(new_n292), .ZN(G1340gat));
  NOR2_X1   g682(.A1(new_n881), .A2(new_n699), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(new_n293), .ZN(G1341gat));
  OAI21_X1  g684(.A(new_n303), .B1(new_n881), .B2(new_n730), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n622), .A2(new_n298), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n881), .B2(new_n887), .ZN(G1342gat));
  NOR2_X1   g687(.A1(new_n535), .A2(new_n677), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT118), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n880), .A2(new_n301), .A3(new_n533), .A4(new_n890), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT56), .Z(new_n892));
  OAI21_X1  g691(.A(G134gat), .B1(new_n881), .B2(new_n677), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1343gat));
  NOR3_X1   g693(.A1(new_n715), .A2(new_n703), .A3(new_n716), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n268), .A2(new_n275), .A3(new_n282), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n282), .B1(new_n268), .B2(new_n275), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n863), .B(new_n868), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n285), .A2(new_n698), .A3(new_n872), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n898), .A2(new_n899), .B1(new_n744), .B2(new_n740), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n863), .A2(new_n868), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n745), .A2(new_n901), .A3(new_n873), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n730), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n853), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n578), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n287), .A2(G141gat), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n895), .A2(new_n794), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT58), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT119), .B1(new_n905), .B2(KEYINPUT57), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n912), .B(new_n913), .C1(new_n879), .C2(new_n578), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n861), .A2(new_n862), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n286), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n737), .B1(new_n916), .B2(new_n899), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n622), .B1(new_n918), .B2(new_n875), .ZN(new_n919));
  OAI211_X1 g718(.A(KEYINPUT57), .B(new_n506), .C1(new_n919), .C2(new_n853), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n911), .A2(new_n914), .A3(new_n920), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n713), .A2(new_n703), .A3(new_n835), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n286), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G141gat), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n910), .B(new_n924), .C1(new_n909), .C2(new_n908), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n923), .A2(new_n926), .A3(G141gat), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n923), .B2(G141gat), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n927), .A2(new_n928), .A3(new_n908), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT58), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n925), .B1(new_n929), .B2(new_n930), .ZN(G1344gat));
  AND2_X1   g730(.A1(new_n895), .A2(new_n905), .ZN(new_n932));
  INV_X1    g731(.A(G148gat), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n932), .A2(new_n933), .A3(new_n698), .A4(new_n794), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n921), .A2(new_n922), .ZN(new_n935));
  AOI211_X1 g734(.A(KEYINPUT59), .B(new_n933), .C1(new_n935), .C2(new_n698), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT59), .ZN(new_n937));
  NOR4_X1   g736(.A1(new_n873), .A2(new_n677), .A3(new_n862), .A4(new_n861), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n788), .B1(new_n917), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n578), .B1(new_n939), .B2(new_n904), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n941));
  OR3_X1    g740(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT57), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n905), .A2(KEYINPUT57), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n940), .B2(KEYINPUT57), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n698), .A3(new_n922), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n937), .B1(new_n946), .B2(G148gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n934), .B1(new_n936), .B2(new_n947), .ZN(G1345gat));
  AOI21_X1  g747(.A(new_n313), .B1(new_n935), .B2(new_n731), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n950));
  AND4_X1   g749(.A1(new_n313), .A2(new_n932), .A3(new_n622), .A4(new_n794), .ZN(new_n951));
  OR3_X1    g750(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1346gat));
  NAND3_X1  g753(.A1(new_n932), .A2(new_n314), .A3(new_n890), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n935), .A2(new_n746), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n314), .ZN(G1347gat));
  NOR4_X1   g756(.A1(new_n879), .A2(new_n533), .A3(new_n506), .A4(new_n768), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(new_n835), .ZN(new_n959));
  AOI21_X1  g758(.A(G169gat), .B1(new_n959), .B2(new_n286), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n535), .ZN(new_n961));
  INV_X1    g760(.A(G169gat), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n961), .A2(new_n962), .A3(new_n287), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n960), .A2(new_n963), .ZN(G1348gat));
  AOI21_X1  g763(.A(G176gat), .B1(new_n959), .B2(new_n698), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n961), .A2(new_n424), .A3(new_n699), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(new_n966), .ZN(G1349gat));
  NAND3_X1  g766(.A1(new_n959), .A2(new_n398), .A3(new_n622), .ZN(new_n968));
  OAI21_X1  g767(.A(G183gat), .B1(new_n961), .B2(new_n730), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n970), .B(new_n971), .Z(G1350gat));
  NAND3_X1  g771(.A1(new_n959), .A2(new_n402), .A3(new_n746), .ZN(new_n973));
  OAI21_X1  g772(.A(G190gat), .B1(new_n961), .B2(new_n677), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n974), .A2(KEYINPUT61), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n974), .A2(KEYINPUT61), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1351gat));
  NAND2_X1  g776(.A1(new_n835), .A2(new_n506), .ZN(new_n978));
  NOR4_X1   g777(.A1(new_n717), .A2(new_n533), .A3(new_n879), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(G197gat), .B1(new_n979), .B2(new_n286), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n945), .A2(KEYINPUT125), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n942), .A2(new_n982), .A3(new_n943), .A4(new_n944), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n717), .A2(new_n533), .A3(new_n534), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n286), .A2(G197gat), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n980), .B1(new_n986), .B2(new_n987), .ZN(G1352gat));
  XNOR2_X1  g787(.A(KEYINPUT126), .B(G204gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n989), .B1(new_n985), .B2(new_n699), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n699), .A2(new_n989), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n979), .A2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n993), .A2(KEYINPUT127), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n993), .A2(KEYINPUT127), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n990), .A2(new_n995), .A3(new_n997), .ZN(G1353gat));
  NAND3_X1  g797(.A1(new_n979), .A2(new_n384), .A3(new_n622), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n945), .A2(new_n622), .A3(new_n984), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n1000), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1001));
  AOI21_X1  g800(.A(KEYINPUT63), .B1(new_n1000), .B2(G211gat), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(G1354gat));
  AOI21_X1  g802(.A(G218gat), .B1(new_n979), .B2(new_n746), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n677), .A2(new_n385), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1004), .B1(new_n986), .B2(new_n1005), .ZN(G1355gat));
endmodule


