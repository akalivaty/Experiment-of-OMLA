

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  OR2_X1 U324 ( .A1(n480), .A2(n413), .ZN(n414) );
  XOR2_X1 U325 ( .A(n323), .B(n322), .Z(n292) );
  NOR2_X1 U326 ( .A1(n348), .A2(n347), .ZN(n349) );
  OR2_X1 U327 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U328 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U329 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U330 ( .A(n318), .B(n317), .ZN(n321) );
  XNOR2_X1 U331 ( .A(n434), .B(n433), .ZN(n438) );
  XNOR2_X1 U332 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n466) );
  XNOR2_X1 U333 ( .A(n467), .B(n466), .ZN(n527) );
  XNOR2_X1 U334 ( .A(n345), .B(KEYINPUT26), .ZN(n542) );
  INV_X1 U335 ( .A(n542), .ZN(n544) );
  INV_X1 U336 ( .A(KEYINPUT59), .ZN(n474) );
  XNOR2_X1 U337 ( .A(n454), .B(KEYINPUT65), .ZN(n551) );
  XNOR2_X1 U338 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U339 ( .A(n447), .B(G36GAT), .ZN(n448) );
  XNOR2_X1 U340 ( .A(n477), .B(n476), .ZN(G1352GAT) );
  XNOR2_X1 U341 ( .A(n449), .B(n448), .ZN(G1329GAT) );
  XOR2_X1 U342 ( .A(G211GAT), .B(KEYINPUT21), .Z(n294) );
  XNOR2_X1 U343 ( .A(G197GAT), .B(G218GAT), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n319) );
  XOR2_X1 U345 ( .A(KEYINPUT91), .B(n319), .Z(n296) );
  NAND2_X1 U346 ( .A1(G226GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n299) );
  XOR2_X1 U348 ( .A(G64GAT), .B(G92GAT), .Z(n298) );
  XNOR2_X1 U349 ( .A(G176GAT), .B(G204GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n439) );
  XOR2_X1 U351 ( .A(n299), .B(n439), .Z(n305) );
  XNOR2_X1 U352 ( .A(G169GAT), .B(G36GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n300), .B(G8GAT), .ZN(n416) );
  XOR2_X1 U354 ( .A(KEYINPUT17), .B(G190GAT), .Z(n302) );
  XNOR2_X1 U355 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U357 ( .A(KEYINPUT19), .B(n303), .Z(n332) );
  XNOR2_X1 U358 ( .A(n416), .B(n332), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n517) );
  XOR2_X1 U360 ( .A(KEYINPUT100), .B(KEYINPUT37), .Z(n415) );
  INV_X1 U361 ( .A(KEYINPUT94), .ZN(n369) );
  XOR2_X1 U362 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n307) );
  XNOR2_X1 U363 ( .A(G141GAT), .B(G155GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n309) );
  XOR2_X1 U365 ( .A(G162GAT), .B(KEYINPUT3), .Z(n308) );
  XOR2_X1 U366 ( .A(n309), .B(n308), .Z(n364) );
  XOR2_X1 U367 ( .A(KEYINPUT83), .B(KEYINPUT85), .Z(n311) );
  XNOR2_X1 U368 ( .A(KEYINPUT22), .B(G204GAT), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n323) );
  XOR2_X1 U370 ( .A(G148GAT), .B(G78GAT), .Z(n430) );
  XOR2_X1 U371 ( .A(G106GAT), .B(KEYINPUT73), .Z(n313) );
  XNOR2_X1 U372 ( .A(G50GAT), .B(G22GAT), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U374 ( .A(n430), .B(n314), .Z(n318) );
  NAND2_X1 U375 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  INV_X1 U376 ( .A(KEYINPUT23), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n319), .B(KEYINPUT24), .ZN(n320) );
  XNOR2_X1 U378 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U379 ( .A(n364), .B(n292), .Z(n560) );
  XOR2_X1 U380 ( .A(G127GAT), .B(KEYINPUT77), .Z(n325) );
  XNOR2_X1 U381 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n354) );
  XOR2_X1 U383 ( .A(n354), .B(G99GAT), .Z(n327) );
  NAND2_X1 U384 ( .A1(G227GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U386 ( .A(G71GAT), .B(G176GAT), .Z(n329) );
  XNOR2_X1 U387 ( .A(G169GAT), .B(G15GAT), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U389 ( .A(n331), .B(n330), .Z(n334) );
  XNOR2_X1 U390 ( .A(G43GAT), .B(n332), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n342) );
  XOR2_X1 U392 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n336) );
  XNOR2_X1 U393 ( .A(KEYINPUT80), .B(G120GAT), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U395 ( .A(KEYINPUT20), .B(KEYINPUT78), .Z(n338) );
  XNOR2_X1 U396 ( .A(G113GAT), .B(KEYINPUT79), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U398 ( .A(n340), .B(n339), .Z(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n563) );
  NOR2_X1 U400 ( .A1(n517), .A2(n563), .ZN(n343) );
  NOR2_X1 U401 ( .A1(n560), .A2(n343), .ZN(n344) );
  XOR2_X1 U402 ( .A(KEYINPUT25), .B(n344), .Z(n348) );
  NAND2_X1 U403 ( .A1(n563), .A2(n560), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n517), .B(KEYINPUT27), .ZN(n371) );
  NOR2_X1 U405 ( .A1(n542), .A2(n371), .ZN(n346) );
  XNOR2_X1 U406 ( .A(KEYINPUT92), .B(n346), .ZN(n347) );
  XNOR2_X1 U407 ( .A(KEYINPUT93), .B(n349), .ZN(n367) );
  XNOR2_X1 U408 ( .A(G120GAT), .B(G85GAT), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n350), .B(G57GAT), .ZN(n440) );
  XOR2_X1 U410 ( .A(G113GAT), .B(G1GAT), .Z(n424) );
  XOR2_X1 U411 ( .A(n440), .B(n424), .Z(n352) );
  NAND2_X1 U412 ( .A1(G225GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U414 ( .A(n353), .B(KEYINPUT88), .Z(n356) );
  XNOR2_X1 U415 ( .A(n354), .B(KEYINPUT4), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U417 ( .A(KEYINPUT87), .B(KEYINPUT5), .Z(n358) );
  XNOR2_X1 U418 ( .A(G29GAT), .B(G148GAT), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U420 ( .A(n360), .B(n359), .Z(n366) );
  XOR2_X1 U421 ( .A(KEYINPUT6), .B(KEYINPUT86), .Z(n362) );
  XNOR2_X1 U422 ( .A(KEYINPUT89), .B(KEYINPUT1), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n370) );
  NAND2_X1 U426 ( .A1(n367), .A2(n370), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n375) );
  XOR2_X1 U428 ( .A(n560), .B(KEYINPUT28), .Z(n528) );
  INV_X1 U429 ( .A(n528), .ZN(n373) );
  XNOR2_X1 U430 ( .A(KEYINPUT90), .B(n370), .ZN(n514) );
  NOR2_X1 U431 ( .A1(n514), .A2(n371), .ZN(n525) );
  NAND2_X1 U432 ( .A1(n525), .A2(n563), .ZN(n372) );
  NOR2_X1 U433 ( .A1(n373), .A2(n372), .ZN(n374) );
  NOR2_X1 U434 ( .A1(n375), .A2(n374), .ZN(n480) );
  XOR2_X1 U435 ( .A(G43GAT), .B(G29GAT), .Z(n377) );
  XNOR2_X1 U436 ( .A(KEYINPUT7), .B(KEYINPUT68), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U438 ( .A(n378), .B(KEYINPUT67), .Z(n380) );
  XNOR2_X1 U439 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n428) );
  XOR2_X1 U441 ( .A(KEYINPUT9), .B(G92GAT), .Z(n382) );
  XNOR2_X1 U442 ( .A(G190GAT), .B(G134GAT), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n428), .B(n383), .ZN(n397) );
  XOR2_X1 U445 ( .A(KEYINPUT74), .B(KEYINPUT10), .Z(n385) );
  XNOR2_X1 U446 ( .A(KEYINPUT73), .B(G85GAT), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U448 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n387) );
  XNOR2_X1 U449 ( .A(G36GAT), .B(KEYINPUT11), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U451 ( .A(n389), .B(n388), .Z(n395) );
  XNOR2_X1 U452 ( .A(G99GAT), .B(G106GAT), .ZN(n390) );
  XNOR2_X1 U453 ( .A(n390), .B(KEYINPUT71), .ZN(n434) );
  XOR2_X1 U454 ( .A(n434), .B(G218GAT), .Z(n392) );
  NAND2_X1 U455 ( .A1(G232GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U457 ( .A(G162GAT), .B(n393), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U459 ( .A(n397), .B(n396), .Z(n574) );
  XOR2_X1 U460 ( .A(n574), .B(KEYINPUT36), .Z(n585) );
  XNOR2_X1 U461 ( .A(G183GAT), .B(G127GAT), .ZN(n399) );
  XNOR2_X1 U462 ( .A(G15GAT), .B(G22GAT), .ZN(n423) );
  INV_X1 U463 ( .A(n423), .ZN(n398) );
  XOR2_X1 U464 ( .A(n399), .B(n398), .Z(n412) );
  XOR2_X1 U465 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n401) );
  NAND2_X1 U466 ( .A1(G231GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U468 ( .A(KEYINPUT14), .B(G64GAT), .Z(n403) );
  XNOR2_X1 U469 ( .A(G8GAT), .B(G57GAT), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U471 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U472 ( .A(G71GAT), .B(KEYINPUT13), .Z(n429) );
  XOR2_X1 U473 ( .A(G78GAT), .B(G211GAT), .Z(n407) );
  XNOR2_X1 U474 ( .A(G1GAT), .B(G155GAT), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n429), .B(n408), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U478 ( .A(n412), .B(n411), .Z(n583) );
  INV_X1 U479 ( .A(n583), .ZN(n571) );
  OR2_X1 U480 ( .A1(n585), .A2(n571), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n513) );
  XOR2_X1 U482 ( .A(n416), .B(KEYINPUT30), .Z(n418) );
  NAND2_X1 U483 ( .A1(G229GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U485 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n420) );
  XNOR2_X1 U486 ( .A(G141GAT), .B(G197GAT), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U488 ( .A(n422), .B(n421), .Z(n426) );
  XOR2_X1 U489 ( .A(n424), .B(n423), .Z(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n546) );
  XOR2_X1 U492 ( .A(KEYINPUT69), .B(n546), .Z(n461) );
  INV_X1 U493 ( .A(n461), .ZN(n564) );
  XNOR2_X1 U494 ( .A(n430), .B(n429), .ZN(n444) );
  NAND2_X1 U495 ( .A1(G230GAT), .A2(G233GAT), .ZN(n432) );
  INV_X1 U496 ( .A(KEYINPUT31), .ZN(n431) );
  XOR2_X1 U497 ( .A(KEYINPUT70), .B(KEYINPUT32), .Z(n436) );
  XNOR2_X1 U498 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U501 ( .A(n440), .B(n439), .Z(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n579) );
  NAND2_X1 U504 ( .A1(n564), .A2(n579), .ZN(n482) );
  NOR2_X1 U505 ( .A1(n513), .A2(n482), .ZN(n446) );
  XNOR2_X1 U506 ( .A(KEYINPUT38), .B(KEYINPUT101), .ZN(n445) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n501) );
  NOR2_X1 U508 ( .A1(n517), .A2(n501), .ZN(n449) );
  XNOR2_X1 U509 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n447) );
  NAND2_X1 U510 ( .A1(n579), .A2(KEYINPUT41), .ZN(n453) );
  INV_X1 U511 ( .A(n579), .ZN(n451) );
  INV_X1 U512 ( .A(KEYINPUT41), .ZN(n450) );
  NAND2_X1 U513 ( .A1(n451), .A2(n450), .ZN(n452) );
  NAND2_X1 U514 ( .A1(n453), .A2(n452), .ZN(n454) );
  NOR2_X1 U515 ( .A1(n551), .A2(n546), .ZN(n455) );
  XNOR2_X1 U516 ( .A(n455), .B(KEYINPUT46), .ZN(n457) );
  INV_X1 U517 ( .A(n574), .ZN(n557) );
  NAND2_X1 U518 ( .A1(n583), .A2(n557), .ZN(n456) );
  XNOR2_X1 U519 ( .A(KEYINPUT47), .B(n458), .ZN(n465) );
  NOR2_X1 U520 ( .A1(n585), .A2(n583), .ZN(n460) );
  XNOR2_X1 U521 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n459) );
  XNOR2_X1 U522 ( .A(n460), .B(n459), .ZN(n463) );
  NAND2_X1 U523 ( .A1(n579), .A2(n461), .ZN(n462) );
  NOR2_X1 U524 ( .A1(n463), .A2(n462), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n517), .B(KEYINPUT120), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n527), .A2(n468), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n469), .B(KEYINPUT54), .ZN(n470) );
  NAND2_X1 U529 ( .A1(n470), .A2(n514), .ZN(n559) );
  NOR2_X1 U530 ( .A1(n542), .A2(n559), .ZN(n471) );
  XOR2_X1 U531 ( .A(KEYINPUT124), .B(n471), .Z(n586) );
  NOR2_X1 U532 ( .A1(n586), .A2(n546), .ZN(n473) );
  XNOR2_X1 U533 ( .A(KEYINPUT60), .B(KEYINPUT126), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U535 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n475) );
  INV_X1 U536 ( .A(KEYINPUT96), .ZN(n484) );
  NOR2_X1 U537 ( .A1(n574), .A2(n583), .ZN(n478) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n478), .Z(n479) );
  NOR2_X1 U539 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U540 ( .A(KEYINPUT95), .B(n481), .ZN(n503) );
  NOR2_X1 U541 ( .A1(n503), .A2(n482), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n489) );
  NOR2_X1 U543 ( .A1(n489), .A2(n514), .ZN(n485) );
  XOR2_X1 U544 ( .A(KEYINPUT34), .B(n485), .Z(n486) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  XNOR2_X1 U546 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n488) );
  NOR2_X1 U547 ( .A1(n517), .A2(n489), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(G1325GAT) );
  NOR2_X1 U549 ( .A1(n489), .A2(n563), .ZN(n491) );
  XNOR2_X1 U550 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G15GAT), .B(n492), .ZN(G1326GAT) );
  XNOR2_X1 U553 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n494) );
  NOR2_X1 U554 ( .A1(n528), .A2(n489), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1327GAT) );
  NOR2_X1 U556 ( .A1(n501), .A2(n514), .ZN(n496) );
  XNOR2_X1 U557 ( .A(KEYINPUT39), .B(KEYINPUT102), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U560 ( .A1(n501), .A2(n563), .ZN(n499) );
  XNOR2_X1 U561 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NOR2_X1 U564 ( .A1(n528), .A2(n501), .ZN(n502) );
  XOR2_X1 U565 ( .A(G50GAT), .B(n502), .Z(G1331GAT) );
  XOR2_X1 U566 ( .A(n551), .B(KEYINPUT106), .Z(n567) );
  NAND2_X1 U567 ( .A1(n567), .A2(n546), .ZN(n512) );
  OR2_X1 U568 ( .A1(n503), .A2(n512), .ZN(n509) );
  NOR2_X1 U569 ( .A1(n514), .A2(n509), .ZN(n504) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n504), .Z(n505) );
  XNOR2_X1 U571 ( .A(KEYINPUT42), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U572 ( .A1(n517), .A2(n509), .ZN(n507) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(G1333GAT) );
  NOR2_X1 U575 ( .A1(n563), .A2(n509), .ZN(n508) );
  XOR2_X1 U576 ( .A(G71GAT), .B(n508), .Z(G1334GAT) );
  NOR2_X1 U577 ( .A1(n528), .A2(n509), .ZN(n511) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  OR2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n521) );
  NOR2_X1 U581 ( .A1(n514), .A2(n521), .ZN(n515) );
  XOR2_X1 U582 ( .A(n515), .B(KEYINPUT108), .Z(n516) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n517), .A2(n521), .ZN(n518) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n563), .A2(n521), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  NOR2_X1 U589 ( .A1(n528), .A2(n521), .ZN(n523) );
  XNOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n524), .Z(G1339GAT) );
  INV_X1 U593 ( .A(n525), .ZN(n526) );
  NOR2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n543) );
  NAND2_X1 U595 ( .A1(n528), .A2(n543), .ZN(n529) );
  NOR2_X1 U596 ( .A1(n563), .A2(n529), .ZN(n530) );
  XNOR2_X1 U597 ( .A(KEYINPUT112), .B(n530), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n564), .A2(n539), .ZN(n531) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U601 ( .A1(n567), .A2(n539), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n534), .Z(G1341GAT) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n538) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n536) );
  NAND2_X1 U606 ( .A1(n571), .A2(n539), .ZN(n535) );
  XNOR2_X1 U607 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U608 ( .A(n538), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U610 ( .A1(n539), .A2(n574), .ZN(n540) );
  XNOR2_X1 U611 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n545), .B(KEYINPUT116), .ZN(n556) );
  NOR2_X1 U614 ( .A1(n556), .A2(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(n553) );
  NOR2_X1 U620 ( .A1(n551), .A2(n556), .ZN(n552) );
  XOR2_X1 U621 ( .A(n553), .B(n552), .Z(G1345GAT) );
  NOR2_X1 U622 ( .A1(n556), .A2(n583), .ZN(n555) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  XOR2_X1 U627 ( .A(G169GAT), .B(KEYINPUT121), .Z(n566) );
  NOR2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n561), .B(KEYINPUT55), .ZN(n562) );
  NOR2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n575), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n569) );
  NAND2_X1 U634 ( .A1(n567), .A2(n575), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(n570), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n575), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT122), .ZN(n573) );
  XNOR2_X1 U639 ( .A(G183GAT), .B(n573), .ZN(G1350GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n577) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G190GAT), .B(n578), .ZN(G1351GAT) );
  XNOR2_X1 U644 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n581) );
  NOR2_X1 U645 ( .A1(n579), .A2(n586), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(G204GAT), .B(n582), .Z(G1353GAT) );
  NOR2_X1 U648 ( .A1(n586), .A2(n583), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

