

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599;

  XNOR2_X1 U327 ( .A(n424), .B(n423), .ZN(n425) );
  INV_X1 U328 ( .A(KEYINPUT37), .ZN(n423) );
  XNOR2_X1 U329 ( .A(KEYINPUT38), .B(n467), .ZN(n513) );
  XOR2_X1 U330 ( .A(n341), .B(n340), .Z(n538) );
  XOR2_X1 U331 ( .A(n333), .B(n311), .Z(n532) );
  INV_X1 U332 ( .A(KEYINPUT116), .ZN(n475) );
  XNOR2_X1 U333 ( .A(n475), .B(KEYINPUT47), .ZN(n476) );
  INV_X1 U334 ( .A(G36GAT), .ZN(n305) );
  XNOR2_X1 U335 ( .A(n477), .B(n476), .ZN(n482) );
  XNOR2_X1 U336 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U337 ( .A(n462), .B(n461), .ZN(n463) );
  NOR2_X1 U338 ( .A1(n502), .A2(n374), .ZN(n539) );
  XNOR2_X1 U339 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U340 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U341 ( .A(n426), .B(n425), .ZN(n530) );
  NOR2_X1 U342 ( .A1(n509), .A2(n488), .ZN(n578) );
  XNOR2_X1 U343 ( .A(n489), .B(G190GAT), .ZN(n490) );
  XNOR2_X1 U344 ( .A(n305), .B(KEYINPUT108), .ZN(n468) );
  XNOR2_X1 U345 ( .A(n491), .B(n490), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n469), .B(n468), .ZN(G1329GAT) );
  XNOR2_X1 U347 ( .A(KEYINPUT18), .B(KEYINPUT88), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n295), .B(KEYINPUT89), .ZN(n296) );
  XOR2_X1 U349 ( .A(n296), .B(KEYINPUT17), .Z(n298) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n333) );
  XOR2_X1 U352 ( .A(G190GAT), .B(G92GAT), .Z(n408) );
  XOR2_X1 U353 ( .A(G176GAT), .B(G64GAT), .Z(n447) );
  XOR2_X1 U354 ( .A(KEYINPUT99), .B(n447), .Z(n300) );
  NAND2_X1 U355 ( .A1(G226GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U356 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n408), .B(n301), .ZN(n310) );
  XOR2_X1 U358 ( .A(KEYINPUT91), .B(G211GAT), .Z(n303) );
  XNOR2_X1 U359 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U361 ( .A(G197GAT), .B(n304), .Z(n325) );
  INV_X1 U362 ( .A(n325), .ZN(n308) );
  XOR2_X1 U363 ( .A(G8GAT), .B(G183GAT), .Z(n384) );
  XOR2_X1 U364 ( .A(n384), .B(G218GAT), .Z(n306) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U366 ( .A(KEYINPUT27), .B(n532), .ZN(n373) );
  XOR2_X1 U367 ( .A(G155GAT), .B(KEYINPUT3), .Z(n313) );
  XNOR2_X1 U368 ( .A(KEYINPUT2), .B(KEYINPUT92), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n354) );
  XOR2_X1 U370 ( .A(G218GAT), .B(G162GAT), .Z(n403) );
  XNOR2_X1 U371 ( .A(n354), .B(n403), .ZN(n315) );
  AND2_X1 U372 ( .A1(G228GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U374 ( .A(KEYINPUT24), .B(n316), .Z(n320) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G148GAT), .Z(n318) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n461) );
  XNOR2_X1 U378 ( .A(n461), .B(KEYINPUT23), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n321), .B(KEYINPUT22), .ZN(n323) );
  XOR2_X1 U381 ( .A(G141GAT), .B(G22GAT), .Z(n432) );
  XNOR2_X1 U382 ( .A(G50GAT), .B(n432), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n370) );
  XOR2_X1 U385 ( .A(KEYINPUT90), .B(KEYINPUT87), .Z(n327) );
  XNOR2_X1 U386 ( .A(G43GAT), .B(G183GAT), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n329) );
  XOR2_X1 U388 ( .A(G190GAT), .B(G99GAT), .Z(n328) );
  XNOR2_X1 U389 ( .A(n329), .B(n328), .ZN(n339) );
  XOR2_X1 U390 ( .A(G127GAT), .B(G134GAT), .Z(n331) );
  XNOR2_X1 U391 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U393 ( .A(G113GAT), .B(n332), .Z(n358) );
  XNOR2_X1 U394 ( .A(n358), .B(n333), .ZN(n337) );
  XOR2_X1 U395 ( .A(G176GAT), .B(G71GAT), .Z(n335) );
  XNOR2_X1 U396 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n341) );
  NAND2_X1 U400 ( .A1(G227GAT), .A2(G233GAT), .ZN(n340) );
  INV_X1 U401 ( .A(n538), .ZN(n509) );
  NAND2_X1 U402 ( .A1(n370), .A2(n509), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n342), .B(KEYINPUT101), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n343), .B(KEYINPUT26), .ZN(n583) );
  NAND2_X1 U405 ( .A1(n373), .A2(n583), .ZN(n555) );
  INV_X1 U406 ( .A(n532), .ZN(n484) );
  NOR2_X1 U407 ( .A1(n509), .A2(n484), .ZN(n344) );
  NOR2_X1 U408 ( .A1(n370), .A2(n344), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n345), .B(KEYINPUT25), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n346), .B(KEYINPUT102), .ZN(n347) );
  NAND2_X1 U411 ( .A1(n555), .A2(n347), .ZN(n369) );
  XOR2_X1 U412 ( .A(KEYINPUT96), .B(G57GAT), .Z(n349) );
  XNOR2_X1 U413 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U415 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n351) );
  XNOR2_X1 U416 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U418 ( .A(n353), .B(n352), .Z(n360) );
  XOR2_X1 U419 ( .A(n354), .B(KEYINPUT4), .Z(n356) );
  NAND2_X1 U420 ( .A1(G225GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U421 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n368) );
  XOR2_X1 U424 ( .A(KEYINPUT97), .B(KEYINPUT93), .Z(n362) );
  XNOR2_X1 U425 ( .A(G1GAT), .B(G141GAT), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U427 ( .A(G85GAT), .B(G162GAT), .Z(n364) );
  XNOR2_X1 U428 ( .A(G29GAT), .B(G148GAT), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U430 ( .A(n366), .B(n365), .Z(n367) );
  XOR2_X1 U431 ( .A(n368), .B(n367), .Z(n558) );
  INV_X1 U432 ( .A(n558), .ZN(n505) );
  NAND2_X1 U433 ( .A1(n369), .A2(n505), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n370), .B(KEYINPUT65), .ZN(n372) );
  INV_X1 U435 ( .A(KEYINPUT28), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n502) );
  NAND2_X1 U437 ( .A1(n373), .A2(n558), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n539), .B(KEYINPUT100), .ZN(n375) );
  NAND2_X1 U439 ( .A1(n509), .A2(n375), .ZN(n376) );
  NAND2_X1 U440 ( .A1(n377), .A2(n376), .ZN(n493) );
  INV_X1 U441 ( .A(KEYINPUT13), .ZN(n378) );
  NAND2_X1 U442 ( .A1(KEYINPUT73), .A2(n378), .ZN(n381) );
  INV_X1 U443 ( .A(KEYINPUT73), .ZN(n379) );
  NAND2_X1 U444 ( .A1(n379), .A2(KEYINPUT13), .ZN(n380) );
  NAND2_X1 U445 ( .A1(n381), .A2(n380), .ZN(n383) );
  XNOR2_X1 U446 ( .A(G71GAT), .B(G57GAT), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n383), .B(n382), .ZN(n446) );
  XOR2_X1 U448 ( .A(n446), .B(n384), .Z(n386) );
  NAND2_X1 U449 ( .A1(G231GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U451 ( .A(n387), .B(KEYINPUT12), .Z(n391) );
  XOR2_X1 U452 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n389) );
  XNOR2_X1 U453 ( .A(G15GAT), .B(G1GAT), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n389), .B(n388), .ZN(n436) );
  XNOR2_X1 U455 ( .A(n436), .B(KEYINPUT14), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n399) );
  XOR2_X1 U457 ( .A(G155GAT), .B(G78GAT), .Z(n393) );
  XNOR2_X1 U458 ( .A(G22GAT), .B(G127GAT), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U460 ( .A(KEYINPUT15), .B(KEYINPUT86), .Z(n395) );
  XNOR2_X1 U461 ( .A(G211GAT), .B(G64GAT), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U463 ( .A(n397), .B(n396), .Z(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n592) );
  NAND2_X1 U465 ( .A1(n493), .A2(n592), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n400), .B(KEYINPUT104), .ZN(n422) );
  XOR2_X1 U467 ( .A(KEYINPUT9), .B(KEYINPUT64), .Z(n402) );
  XNOR2_X1 U468 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n404) );
  XOR2_X1 U470 ( .A(n404), .B(n403), .Z(n406) );
  XNOR2_X1 U471 ( .A(G134GAT), .B(G106GAT), .ZN(n405) );
  XNOR2_X1 U472 ( .A(n406), .B(n405), .ZN(n412) );
  XNOR2_X1 U473 ( .A(G99GAT), .B(G85GAT), .ZN(n407) );
  XOR2_X1 U474 ( .A(n407), .B(KEYINPUT76), .Z(n465) );
  XNOR2_X1 U475 ( .A(n465), .B(n408), .ZN(n410) );
  NAND2_X1 U476 ( .A1(G232GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U478 ( .A(n412), .B(n411), .Z(n421) );
  XOR2_X1 U479 ( .A(G29GAT), .B(KEYINPUT8), .Z(n414) );
  XNOR2_X1 U480 ( .A(G43GAT), .B(G36GAT), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U482 ( .A(G50GAT), .B(KEYINPUT7), .Z(n415) );
  XOR2_X1 U483 ( .A(n416), .B(n415), .Z(n441) );
  XOR2_X1 U484 ( .A(KEYINPUT84), .B(KEYINPUT11), .Z(n418) );
  XNOR2_X1 U485 ( .A(KEYINPUT10), .B(KEYINPUT85), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n441), .B(n419), .ZN(n420) );
  XOR2_X1 U488 ( .A(n421), .B(n420), .Z(n567) );
  XNOR2_X1 U489 ( .A(KEYINPUT36), .B(n567), .ZN(n597) );
  NOR2_X1 U490 ( .A1(n422), .A2(n597), .ZN(n426) );
  XNOR2_X1 U491 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n424) );
  XOR2_X1 U492 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n428) );
  XNOR2_X1 U493 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n427) );
  XNOR2_X1 U494 ( .A(n428), .B(n427), .ZN(n440) );
  XOR2_X1 U495 ( .A(G8GAT), .B(G197GAT), .Z(n430) );
  XNOR2_X1 U496 ( .A(G169GAT), .B(G113GAT), .ZN(n429) );
  XNOR2_X1 U497 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U498 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U499 ( .A1(G229GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U500 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U501 ( .A(n435), .B(KEYINPUT69), .Z(n438) );
  XNOR2_X1 U502 ( .A(n436), .B(KEYINPUT66), .ZN(n437) );
  XNOR2_X1 U503 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n442), .B(n441), .ZN(n585) );
  XOR2_X1 U506 ( .A(KEYINPUT72), .B(n585), .Z(n570) );
  XOR2_X1 U507 ( .A(KEYINPUT79), .B(KEYINPUT32), .Z(n444) );
  XNOR2_X1 U508 ( .A(KEYINPUT74), .B(KEYINPUT78), .ZN(n443) );
  XNOR2_X1 U509 ( .A(n444), .B(n443), .ZN(n454) );
  INV_X1 U510 ( .A(n447), .ZN(n445) );
  NAND2_X1 U511 ( .A1(n446), .A2(n445), .ZN(n450) );
  INV_X1 U512 ( .A(n446), .ZN(n448) );
  NAND2_X1 U513 ( .A1(n448), .A2(n447), .ZN(n449) );
  NAND2_X1 U514 ( .A1(n450), .A2(n449), .ZN(n452) );
  NAND2_X1 U515 ( .A1(G230GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U516 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U517 ( .A(n454), .B(n453), .ZN(n464) );
  XOR2_X1 U518 ( .A(KEYINPUT33), .B(G92GAT), .Z(n456) );
  XNOR2_X1 U519 ( .A(G120GAT), .B(G204GAT), .ZN(n455) );
  XNOR2_X1 U520 ( .A(n456), .B(n455), .ZN(n460) );
  XOR2_X1 U521 ( .A(KEYINPUT77), .B(KEYINPUT31), .Z(n458) );
  XNOR2_X1 U522 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n457) );
  XNOR2_X1 U523 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U524 ( .A(n460), .B(n459), .Z(n462) );
  XOR2_X1 U525 ( .A(n466), .B(n465), .Z(n589) );
  NAND2_X1 U526 ( .A1(n570), .A2(n589), .ZN(n495) );
  OR2_X1 U527 ( .A1(n530), .A2(n495), .ZN(n467) );
  NOR2_X1 U528 ( .A1(n513), .A2(n484), .ZN(n469) );
  INV_X1 U529 ( .A(n567), .ZN(n549) );
  INV_X1 U530 ( .A(KEYINPUT41), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n470), .B(n589), .ZN(n561) );
  NOR2_X1 U532 ( .A1(n561), .A2(n585), .ZN(n472) );
  XNOR2_X1 U533 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n471) );
  XNOR2_X1 U534 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U535 ( .A(KEYINPUT114), .B(n592), .ZN(n580) );
  NAND2_X1 U536 ( .A1(n473), .A2(n580), .ZN(n474) );
  NOR2_X1 U537 ( .A1(n549), .A2(n474), .ZN(n477) );
  NOR2_X1 U538 ( .A1(n597), .A2(n592), .ZN(n478) );
  XNOR2_X1 U539 ( .A(KEYINPUT45), .B(n478), .ZN(n479) );
  NAND2_X1 U540 ( .A1(n479), .A2(n589), .ZN(n480) );
  NOR2_X1 U541 ( .A1(n480), .A2(n570), .ZN(n481) );
  NOR2_X1 U542 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U543 ( .A(KEYINPUT48), .B(n483), .ZN(n556) );
  NOR2_X1 U544 ( .A1(n484), .A2(n556), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n485), .B(KEYINPUT54), .ZN(n486) );
  NAND2_X1 U546 ( .A1(n486), .A2(n505), .ZN(n582) );
  NOR2_X1 U547 ( .A1(n582), .A2(n370), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(KEYINPUT55), .ZN(n488) );
  NAND2_X1 U549 ( .A1(n578), .A2(n549), .ZN(n491) );
  XOR2_X1 U550 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n489) );
  XOR2_X1 U551 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n497) );
  NOR2_X1 U552 ( .A1(n549), .A2(n592), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT16), .ZN(n494) );
  NAND2_X1 U554 ( .A1(n494), .A2(n493), .ZN(n520) );
  NOR2_X1 U555 ( .A1(n495), .A2(n520), .ZN(n503) );
  NAND2_X1 U556 ( .A1(n503), .A2(n558), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G1GAT), .B(n498), .ZN(G1324GAT) );
  NAND2_X1 U559 ( .A1(n503), .A2(n532), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U561 ( .A(G15GAT), .B(KEYINPUT35), .Z(n501) );
  NAND2_X1 U562 ( .A1(n503), .A2(n538), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1326GAT) );
  NAND2_X1 U564 ( .A1(n502), .A2(n503), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n504), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U566 ( .A1(n513), .A2(n505), .ZN(n507) );
  XNOR2_X1 U567 ( .A(KEYINPUT107), .B(KEYINPUT39), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U569 ( .A(G29GAT), .B(n508), .Z(G1328GAT) );
  XNOR2_X1 U570 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n511) );
  NOR2_X1 U571 ( .A1(n509), .A2(n513), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U573 ( .A(G43GAT), .B(n512), .ZN(G1330GAT) );
  INV_X1 U574 ( .A(KEYINPUT110), .ZN(n516) );
  INV_X1 U575 ( .A(n502), .ZN(n514) );
  NOR2_X1 U576 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U577 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U578 ( .A(G50GAT), .B(n517), .ZN(G1331GAT) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n518) );
  XNOR2_X1 U580 ( .A(n518), .B(KEYINPUT111), .ZN(n519) );
  XOR2_X1 U581 ( .A(KEYINPUT112), .B(n519), .Z(n522) );
  INV_X1 U582 ( .A(n561), .ZN(n575) );
  NAND2_X1 U583 ( .A1(n585), .A2(n575), .ZN(n529) );
  NOR2_X1 U584 ( .A1(n529), .A2(n520), .ZN(n525) );
  NAND2_X1 U585 ( .A1(n525), .A2(n558), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(G1332GAT) );
  NAND2_X1 U587 ( .A1(n525), .A2(n532), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U589 ( .A1(n538), .A2(n525), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n527) );
  NAND2_X1 U592 ( .A1(n525), .A2(n502), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U594 ( .A(G78GAT), .B(n528), .Z(G1335GAT) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n535) );
  NAND2_X1 U596 ( .A1(n535), .A2(n558), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U598 ( .A1(n532), .A2(n535), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G92GAT), .B(n533), .ZN(G1337GAT) );
  NAND2_X1 U600 ( .A1(n538), .A2(n535), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n534), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U602 ( .A1(n502), .A2(n535), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT44), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  XOR2_X1 U605 ( .A(G113GAT), .B(KEYINPUT117), .Z(n542) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U607 ( .A1(n556), .A2(n540), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n550), .A2(n570), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U611 ( .A1(n550), .A2(n575), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  INV_X1 U613 ( .A(n550), .ZN(n545) );
  NOR2_X1 U614 ( .A1(n580), .A2(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U617 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U619 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n554) );
  XOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT120), .Z(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(G1343GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n566) );
  NOR2_X1 U625 ( .A1(n585), .A2(n566), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G141GAT), .B(KEYINPUT121), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1344GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n566), .ZN(n563) );
  XNOR2_X1 U629 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G148GAT), .B(n564), .ZN(G1345GAT) );
  NOR2_X1 U632 ( .A1(n592), .A2(n566), .ZN(n565) );
  XOR2_X1 U633 ( .A(G155GAT), .B(n565), .Z(G1346GAT) );
  NOR2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U635 ( .A(G162GAT), .B(n568), .Z(n569) );
  XNOR2_X1 U636 ( .A(KEYINPUT122), .B(n569), .ZN(G1347GAT) );
  NAND2_X1 U637 ( .A1(n578), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n573) );
  XNOR2_X1 U640 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n572) );
  XNOR2_X1 U641 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U642 ( .A(KEYINPUT56), .B(n574), .Z(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n575), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(G1349GAT) );
  INV_X1 U645 ( .A(n578), .ZN(n579) );
  NOR2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U647 ( .A(G183GAT), .B(n581), .Z(G1350GAT) );
  INV_X1 U648 ( .A(n582), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n596) );
  NOR2_X1 U650 ( .A1(n585), .A2(n596), .ZN(n587) );
  XNOR2_X1 U651 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G197GAT), .B(n588), .ZN(G1352GAT) );
  NOR2_X1 U654 ( .A1(n589), .A2(n596), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1353GAT) );
  NOR2_X1 U657 ( .A1(n592), .A2(n596), .ZN(n593) );
  XOR2_X1 U658 ( .A(G211GAT), .B(n593), .Z(G1354GAT) );
  XOR2_X1 U659 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n595) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n594) );
  XNOR2_X1 U661 ( .A(n595), .B(n594), .ZN(n599) );
  NOR2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U663 ( .A(n599), .B(n598), .Z(G1355GAT) );
endmodule

