

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776;

  AND2_X1 U375 ( .A1(n735), .A2(n734), .ZN(n443) );
  XNOR2_X1 U376 ( .A(n429), .B(n428), .ZN(n718) );
  NAND2_X1 U377 ( .A1(n430), .A2(n644), .ZN(n429) );
  INV_X1 U378 ( .A(n637), .ZN(n621) );
  NAND2_X1 U379 ( .A1(n373), .A2(n370), .ZN(n582) );
  NOR2_X1 U380 ( .A1(G953), .A2(G237), .ZN(n512) );
  INV_X2 U381 ( .A(G953), .ZN(n768) );
  BUF_X1 U382 ( .A(G143), .Z(n446) );
  XNOR2_X2 U383 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X2 U384 ( .A1(n775), .A2(n415), .ZN(n482) );
  XNOR2_X2 U385 ( .A(n413), .B(KEYINPUT35), .ZN(n775) );
  NOR2_X1 U386 ( .A1(n642), .A2(n584), .ZN(n547) );
  XOR2_X1 U387 ( .A(n728), .B(n727), .Z(n351) );
  XNOR2_X2 U388 ( .A(n590), .B(n589), .ZN(n604) );
  INV_X1 U389 ( .A(n693), .ZN(n642) );
  XNOR2_X2 U390 ( .A(n434), .B(KEYINPUT19), .ZN(n618) );
  XNOR2_X1 U391 ( .A(n401), .B(n596), .ZN(n600) );
  XNOR2_X1 U392 ( .A(n465), .B(n464), .ZN(n577) );
  INV_X1 U393 ( .A(G131), .ZN(n412) );
  XNOR2_X1 U394 ( .A(n736), .B(n737), .ZN(n352) );
  NAND2_X1 U395 ( .A1(n398), .A2(n395), .ZN(n776) );
  NOR2_X1 U396 ( .A1(n438), .A2(n417), .ZN(n416) );
  NOR2_X1 U397 ( .A1(n701), .A2(n700), .ZN(n594) );
  NOR2_X2 U398 ( .A1(n510), .A2(n577), .ZN(n679) );
  XNOR2_X1 U399 ( .A(n524), .B(G472), .ZN(n693) );
  OR2_X1 U400 ( .A1(n655), .A2(G902), .ZN(n524) );
  XNOR2_X1 U401 ( .A(n418), .B(G104), .ZN(n556) );
  XNOR2_X1 U402 ( .A(n412), .B(KEYINPUT71), .ZN(n522) );
  INV_X2 U403 ( .A(G125), .ZN(n393) );
  XOR2_X1 U404 ( .A(KEYINPUT15), .B(G902), .Z(n649) );
  NOR2_X1 U405 ( .A1(n352), .A2(n740), .ZN(G63) );
  XNOR2_X2 U406 ( .A(n550), .B(n743), .ZN(n555) );
  XNOR2_X2 U407 ( .A(G116), .B(G107), .ZN(n502) );
  XNOR2_X1 U408 ( .A(KEYINPUT6), .B(KEYINPUT103), .ZN(n583) );
  AND2_X1 U409 ( .A1(n679), .A2(n388), .ZN(n585) );
  NAND2_X1 U410 ( .A1(n599), .A2(n459), .ZN(n458) );
  INV_X1 U411 ( .A(n364), .ZN(n459) );
  NAND2_X1 U412 ( .A1(n776), .A2(n773), .ZN(n401) );
  INV_X1 U413 ( .A(KEYINPUT77), .ZN(n368) );
  NOR2_X1 U414 ( .A1(n437), .A2(n427), .ZN(n425) );
  INV_X1 U415 ( .A(n460), .ZN(n405) );
  NOR2_X1 U416 ( .A1(n462), .A2(n354), .ZN(n390) );
  AND2_X1 U417 ( .A1(n692), .A2(n642), .ZN(n471) );
  XNOR2_X1 U418 ( .A(n522), .B(G134), .ZN(n756) );
  XNOR2_X1 U419 ( .A(n378), .B(G140), .ZN(n548) );
  INV_X1 U420 ( .A(G137), .ZN(n378) );
  INV_X1 U421 ( .A(G122), .ZN(n418) );
  XNOR2_X1 U422 ( .A(n548), .B(n377), .ZN(n549) );
  INV_X1 U423 ( .A(G104), .ZN(n377) );
  XNOR2_X1 U424 ( .A(G107), .B(G110), .ZN(n468) );
  XNOR2_X1 U425 ( .A(n756), .B(G146), .ZN(n552) );
  AND2_X1 U426 ( .A1(n375), .A2(n374), .ZN(n373) );
  NAND2_X1 U427 ( .A1(n376), .A2(G902), .ZN(n374) );
  OR2_X1 U428 ( .A1(n394), .A2(G902), .ZN(n537) );
  NAND2_X1 U429 ( .A1(n403), .A2(n402), .ZN(n760) );
  NOR2_X1 U430 ( .A1(n460), .A2(n404), .ZN(n402) );
  XNOR2_X1 U431 ( .A(n527), .B(KEYINPUT24), .ZN(n529) );
  XOR2_X1 U432 ( .A(G128), .B(G110), .Z(n527) );
  XOR2_X1 U433 ( .A(G119), .B(KEYINPUT23), .Z(n528) );
  XNOR2_X1 U434 ( .A(n526), .B(n548), .ZN(n757) );
  XOR2_X1 U435 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n499) );
  XNOR2_X1 U436 ( .A(G134), .B(G122), .ZN(n503) );
  INV_X1 U437 ( .A(n679), .ZN(n591) );
  INV_X1 U438 ( .A(KEYINPUT85), .ZN(n564) );
  XNOR2_X1 U439 ( .A(n582), .B(KEYINPUT1), .ZN(n637) );
  INV_X1 U440 ( .A(KEYINPUT33), .ZN(n428) );
  INV_X1 U441 ( .A(n645), .ZN(n430) );
  INV_X1 U442 ( .A(n369), .ZN(n483) );
  AND2_X1 U443 ( .A1(n576), .A2(n574), .ZN(n411) );
  INV_X1 U444 ( .A(n573), .ZN(n574) );
  XNOR2_X1 U445 ( .A(G478), .B(KEYINPUT102), .ZN(n464) );
  OR2_X1 U446 ( .A1(n737), .A2(G902), .ZN(n465) );
  NOR2_X1 U447 ( .A1(n709), .A2(n708), .ZN(n710) );
  INV_X1 U448 ( .A(KEYINPUT73), .ZN(n475) );
  OR2_X1 U449 ( .A1(G237), .A2(G902), .ZN(n563) );
  NAND2_X1 U450 ( .A1(n474), .A2(n372), .ZN(n371) );
  INV_X1 U451 ( .A(G902), .ZN(n372) );
  XNOR2_X1 U452 ( .A(G137), .B(G116), .ZN(n515) );
  XOR2_X1 U453 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n516) );
  XOR2_X1 U454 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n514) );
  NOR2_X1 U455 ( .A1(n601), .A2(n458), .ZN(n457) );
  INV_X1 U456 ( .A(n686), .ZN(n463) );
  NAND2_X1 U457 ( .A1(n601), .A2(n364), .ZN(n461) );
  AND2_X1 U458 ( .A1(n452), .A2(n353), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n440), .B(n558), .ZN(n423) );
  NAND2_X1 U460 ( .A1(n768), .A2(G224), .ZN(n440) );
  XNOR2_X1 U461 ( .A(n470), .B(n469), .ZN(n694) );
  INV_X1 U462 ( .A(KEYINPUT114), .ZN(n469) );
  INV_X1 U463 ( .A(n719), .ZN(n479) );
  XNOR2_X1 U464 ( .A(KEYINPUT38), .B(n588), .ZN(n698) );
  NAND2_X1 U465 ( .A1(G234), .A2(G237), .ZN(n538) );
  XNOR2_X1 U466 ( .A(n497), .B(n450), .ZN(n592) );
  XNOR2_X1 U467 ( .A(n496), .B(G475), .ZN(n450) );
  INV_X1 U468 ( .A(KEYINPUT68), .ZN(n432) );
  XNOR2_X1 U469 ( .A(n419), .B(n556), .ZN(n741) );
  XNOR2_X1 U470 ( .A(n502), .B(n557), .ZN(n419) );
  XNOR2_X1 U471 ( .A(G110), .B(KEYINPUT16), .ZN(n557) );
  XNOR2_X1 U472 ( .A(KEYINPUT12), .B(KEYINPUT96), .ZN(n489) );
  XNOR2_X1 U473 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U474 ( .A(n549), .B(n468), .ZN(n467) );
  XNOR2_X1 U475 ( .A(n477), .B(n476), .ZN(n708) );
  XNOR2_X1 U476 ( .A(KEYINPUT52), .B(KEYINPUT117), .ZN(n476) );
  NAND2_X1 U477 ( .A1(n478), .A2(n356), .ZN(n477) );
  NAND2_X1 U478 ( .A1(n355), .A2(n479), .ZN(n478) );
  AND2_X1 U479 ( .A1(n451), .A2(KEYINPUT2), .ZN(n384) );
  OR2_X1 U480 ( .A1(n554), .A2(n582), .ZN(n595) );
  NAND2_X1 U481 ( .A1(n484), .A2(n638), .ZN(n369) );
  XNOR2_X1 U482 ( .A(n592), .B(KEYINPUT100), .ZN(n510) );
  XNOR2_X1 U483 ( .A(n632), .B(KEYINPUT89), .ZN(n646) );
  XNOR2_X1 U484 ( .A(n433), .B(n531), .ZN(n394) );
  XNOR2_X1 U485 ( .A(n757), .B(n530), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U487 ( .A(n509), .B(n508), .ZN(n737) );
  XNOR2_X1 U488 ( .A(n454), .B(n453), .ZN(n773) );
  XNOR2_X1 U489 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n453) );
  OR2_X1 U490 ( .A1(n595), .A2(n719), .ZN(n454) );
  NAND2_X1 U491 ( .A1(n397), .A2(n396), .ZN(n395) );
  AND2_X1 U492 ( .A1(n400), .A2(n399), .ZN(n398) );
  NOR2_X1 U493 ( .A1(n637), .A2(n587), .ZN(n684) );
  NOR2_X1 U494 ( .A1(n369), .A2(n640), .ZN(n437) );
  AND2_X1 U495 ( .A1(n406), .A2(n411), .ZN(n675) );
  NOR2_X1 U496 ( .A1(n621), .A2(n485), .ZN(n427) );
  NOR2_X2 U497 ( .A1(n625), .A2(n624), .ZN(n668) );
  OR2_X1 U498 ( .A1(n646), .A2(n693), .ZN(n624) );
  INV_X1 U499 ( .A(KEYINPUT56), .ZN(n441) );
  NAND2_X1 U500 ( .A1(n445), .A2(n734), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n729), .B(n351), .ZN(n445) );
  NOR2_X1 U502 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U503 ( .A(n693), .B(n583), .ZN(n644) );
  INV_X1 U504 ( .A(n644), .ZN(n484) );
  OR2_X1 U505 ( .A1(n652), .A2(n651), .ZN(n353) );
  NAND2_X1 U506 ( .A1(n772), .A2(n649), .ZN(n354) );
  XNOR2_X1 U507 ( .A(KEYINPUT51), .B(n696), .ZN(n355) );
  XOR2_X1 U508 ( .A(n707), .B(KEYINPUT116), .Z(n356) );
  XOR2_X1 U509 ( .A(n490), .B(n489), .Z(n357) );
  AND2_X1 U510 ( .A1(n635), .A2(n666), .ZN(n358) );
  INV_X1 U511 ( .A(n474), .ZN(n376) );
  XNOR2_X1 U512 ( .A(n475), .B(G469), .ZN(n474) );
  OR2_X1 U513 ( .A1(n483), .A2(n439), .ZN(n359) );
  XOR2_X1 U514 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n360) );
  AND2_X1 U515 ( .A1(n426), .A2(n427), .ZN(n361) );
  OR2_X1 U516 ( .A1(n651), .A2(n711), .ZN(n362) );
  XOR2_X1 U517 ( .A(n663), .B(n662), .Z(n363) );
  XOR2_X1 U518 ( .A(n602), .B(KEYINPUT48), .Z(n364) );
  NOR2_X1 U519 ( .A1(G952), .A2(n768), .ZN(n740) );
  XNOR2_X1 U520 ( .A(n560), .B(KEYINPUT10), .ZN(n526) );
  BUF_X1 U521 ( .A(n520), .Z(n365) );
  XNOR2_X1 U522 ( .A(n446), .B(G113), .ZN(n491) );
  NAND2_X1 U523 ( .A1(n618), .A2(n617), .ZN(n620) );
  XNOR2_X1 U524 ( .A(n416), .B(n643), .ZN(n415) );
  BUF_X1 U525 ( .A(n775), .Z(n366) );
  BUF_X1 U526 ( .A(n730), .Z(n738) );
  NAND2_X1 U527 ( .A1(n353), .A2(KEYINPUT67), .ZN(n392) );
  NAND2_X1 U528 ( .A1(n381), .A2(n711), .ZN(n383) );
  NAND2_X1 U529 ( .A1(n449), .A2(n367), .ZN(n601) );
  XNOR2_X1 U530 ( .A(n581), .B(n368), .ZN(n367) );
  AND2_X1 U531 ( .A1(n648), .A2(n609), .ZN(n410) );
  NOR2_X1 U532 ( .A1(n713), .A2(n380), .ZN(n715) );
  NAND2_X1 U533 ( .A1(n385), .A2(n714), .ZN(n653) );
  NAND2_X1 U534 ( .A1(n420), .A2(n359), .ZN(n438) );
  OR2_X1 U535 ( .A1(n661), .A2(n371), .ZN(n370) );
  NAND2_X1 U536 ( .A1(n661), .A2(n376), .ZN(n375) );
  INV_X1 U537 ( .A(n379), .ZN(n426) );
  NAND2_X1 U538 ( .A1(n379), .A2(n640), .ZN(n420) );
  XNOR2_X2 U539 ( .A(n633), .B(KEYINPUT22), .ZN(n379) );
  NOR2_X1 U540 ( .A1(n425), .A2(n379), .ZN(n417) );
  INV_X1 U541 ( .A(n383), .ZN(n380) );
  INV_X1 U542 ( .A(n650), .ZN(n381) );
  NAND2_X1 U543 ( .A1(n382), .A2(n392), .ZN(n385) );
  NAND2_X1 U544 ( .A1(n383), .A2(n391), .ZN(n382) );
  NAND2_X1 U545 ( .A1(n384), .A2(n650), .ZN(n714) );
  XNOR2_X2 U546 ( .A(n480), .B(KEYINPUT45), .ZN(n650) );
  NOR2_X1 U547 ( .A1(n732), .A2(G902), .ZN(n497) );
  XNOR2_X1 U548 ( .A(n495), .B(n386), .ZN(n732) );
  XNOR2_X1 U549 ( .A(n387), .B(n493), .ZN(n386) );
  XNOR2_X1 U550 ( .A(n357), .B(n494), .ZN(n387) );
  INV_X1 U551 ( .A(n584), .ZN(n388) );
  NAND2_X1 U552 ( .A1(n389), .A2(n362), .ZN(n452) );
  NAND2_X1 U553 ( .A1(n390), .A2(n405), .ZN(n389) );
  XNOR2_X2 U554 ( .A(n393), .B(G146), .ZN(n560) );
  XNOR2_X1 U555 ( .A(n739), .B(n394), .ZN(n444) );
  NOR2_X1 U556 ( .A1(n591), .A2(n360), .ZN(n396) );
  INV_X1 U557 ( .A(n604), .ZN(n397) );
  NAND2_X1 U558 ( .A1(n591), .A2(n360), .ZN(n399) );
  NAND2_X1 U559 ( .A1(n604), .A2(n360), .ZN(n400) );
  INV_X1 U560 ( .A(n462), .ZN(n403) );
  INV_X1 U561 ( .A(n772), .ZN(n404) );
  AND2_X1 U562 ( .A1(n410), .A2(n575), .ZN(n406) );
  NAND2_X1 U563 ( .A1(n411), .A2(n407), .ZN(n590) );
  AND2_X1 U564 ( .A1(n575), .A2(n698), .ZN(n407) );
  AND2_X1 U565 ( .A1(n426), .A2(n484), .ZN(n639) );
  NOR2_X2 U566 ( .A1(n646), .A2(n718), .ZN(n647) );
  XNOR2_X1 U567 ( .A(n647), .B(KEYINPUT34), .ZN(n414) );
  NAND2_X1 U568 ( .A1(n408), .A2(n456), .ZN(n462) );
  NAND2_X1 U569 ( .A1(n455), .A2(n364), .ZN(n408) );
  XNOR2_X2 U570 ( .A(n409), .B(n432), .ZN(n431) );
  NAND2_X1 U571 ( .A1(n641), .A2(n630), .ZN(n409) );
  NAND2_X1 U572 ( .A1(n414), .A2(n648), .ZN(n413) );
  XNOR2_X1 U573 ( .A(n555), .B(n421), .ZN(n728) );
  XNOR2_X1 U574 ( .A(n741), .B(n422), .ZN(n421) );
  XNOR2_X1 U575 ( .A(n424), .B(n423), .ZN(n422) );
  XNOR2_X1 U576 ( .A(n560), .B(n559), .ZN(n424) );
  XNOR2_X2 U577 ( .A(n759), .B(G101), .ZN(n550) );
  XNOR2_X2 U578 ( .A(n520), .B(n519), .ZN(n759) );
  NAND2_X1 U579 ( .A1(n426), .A2(n437), .ZN(n436) );
  XNOR2_X2 U580 ( .A(n620), .B(n619), .ZN(n632) );
  NAND2_X1 U581 ( .A1(n621), .A2(n431), .ZN(n645) );
  NAND2_X1 U582 ( .A1(n431), .A2(n570), .ZN(n625) );
  NOR2_X1 U583 ( .A1(n621), .A2(n431), .ZN(n687) );
  NOR2_X1 U584 ( .A1(n605), .A2(n434), .ZN(n586) );
  XNOR2_X2 U585 ( .A(n565), .B(n564), .ZN(n434) );
  NAND2_X1 U586 ( .A1(n435), .A2(n436), .ZN(n774) );
  INV_X1 U587 ( .A(n438), .ZN(n435) );
  INV_X1 U588 ( .A(n640), .ZN(n439) );
  XNOR2_X1 U589 ( .A(n442), .B(n441), .ZN(G51) );
  XNOR2_X1 U590 ( .A(n443), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X1 U591 ( .A1(n444), .A2(n740), .ZN(G66) );
  XNOR2_X1 U592 ( .A(n448), .B(n447), .ZN(n655) );
  XNOR2_X1 U593 ( .A(n552), .B(n523), .ZN(n447) );
  INV_X1 U594 ( .A(n555), .ZN(n448) );
  XNOR2_X1 U595 ( .A(n684), .B(KEYINPUT83), .ZN(n449) );
  INV_X1 U596 ( .A(n760), .ZN(n451) );
  NAND2_X1 U597 ( .A1(n600), .A2(n599), .ZN(n455) );
  NAND2_X1 U598 ( .A1(n457), .A2(n600), .ZN(n456) );
  NAND2_X1 U599 ( .A1(n461), .A2(n463), .ZN(n460) );
  XNOR2_X1 U600 ( .A(n553), .B(n466), .ZN(n661) );
  XNOR2_X1 U601 ( .A(n550), .B(n467), .ZN(n466) );
  NAND2_X1 U602 ( .A1(n472), .A2(n471), .ZN(n470) );
  XNOR2_X1 U603 ( .A(n687), .B(n473), .ZN(n472) );
  INV_X1 U604 ( .A(KEYINPUT50), .ZN(n473) );
  XNOR2_X2 U605 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n519) );
  NAND2_X1 U606 ( .A1(n481), .A2(n358), .ZN(n480) );
  XNOR2_X1 U607 ( .A(n482), .B(KEYINPUT44), .ZN(n481) );
  NAND2_X1 U608 ( .A1(n642), .A2(n689), .ZN(n485) );
  XNOR2_X1 U609 ( .A(n664), .B(n363), .ZN(n665) );
  XOR2_X1 U610 ( .A(n732), .B(n731), .Z(n486) );
  INV_X1 U611 ( .A(KEYINPUT84), .ZN(n643) );
  INV_X1 U612 ( .A(KEYINPUT72), .ZN(n602) );
  INV_X1 U613 ( .A(KEYINPUT59), .ZN(n731) );
  INV_X1 U614 ( .A(KEYINPUT0), .ZN(n619) );
  INV_X1 U615 ( .A(n740), .ZN(n734) );
  INV_X1 U616 ( .A(KEYINPUT63), .ZN(n659) );
  NOR2_X1 U617 ( .A1(n665), .A2(n740), .ZN(G54) );
  NAND2_X1 U618 ( .A1(G214), .A2(n512), .ZN(n488) );
  INV_X1 U619 ( .A(n526), .ZN(n487) );
  XNOR2_X1 U620 ( .A(n488), .B(n487), .ZN(n495) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n490) );
  XOR2_X1 U622 ( .A(KEYINPUT98), .B(G140), .Z(n492) );
  XNOR2_X1 U623 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U624 ( .A(n522), .B(n556), .ZN(n494) );
  XNOR2_X1 U625 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n496) );
  NAND2_X1 U626 ( .A1(G234), .A2(n768), .ZN(n498) );
  XNOR2_X1 U627 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U628 ( .A(KEYINPUT70), .B(n500), .Z(n525) );
  NAND2_X1 U629 ( .A1(G217), .A2(n525), .ZN(n509) );
  XNOR2_X1 U630 ( .A(KEYINPUT101), .B(KEYINPUT9), .ZN(n507) );
  XNOR2_X2 U631 ( .A(G128), .B(G143), .ZN(n520) );
  INV_X1 U632 ( .A(n365), .ZN(n501) );
  XNOR2_X1 U633 ( .A(n501), .B(KEYINPUT7), .ZN(n505) );
  XNOR2_X1 U634 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U635 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U636 ( .A(n507), .B(n506), .ZN(n508) );
  NAND2_X1 U637 ( .A1(n510), .A2(n577), .ZN(n603) );
  INV_X1 U638 ( .A(n603), .ZN(n681) );
  NOR2_X1 U639 ( .A1(n679), .A2(n681), .ZN(n702) );
  NAND2_X1 U640 ( .A1(n702), .A2(KEYINPUT47), .ZN(n511) );
  XNOR2_X1 U641 ( .A(n511), .B(KEYINPUT78), .ZN(n568) );
  NAND2_X1 U642 ( .A1(n512), .A2(G210), .ZN(n513) );
  XNOR2_X1 U643 ( .A(n514), .B(n513), .ZN(n518) );
  XNOR2_X1 U644 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U645 ( .A(n518), .B(n517), .Z(n523) );
  XOR2_X1 U646 ( .A(G119), .B(G113), .Z(n521) );
  XNOR2_X1 U647 ( .A(KEYINPUT3), .B(n521), .ZN(n743) );
  NAND2_X1 U648 ( .A1(G221), .A2(n525), .ZN(n531) );
  XOR2_X1 U649 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n535) );
  XOR2_X1 U650 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n533) );
  INV_X1 U651 ( .A(n649), .ZN(n651) );
  NAND2_X1 U652 ( .A1(G234), .A2(n651), .ZN(n532) );
  XNOR2_X1 U653 ( .A(n533), .B(n532), .ZN(n544) );
  NAND2_X1 U654 ( .A1(n544), .A2(G217), .ZN(n534) );
  XNOR2_X1 U655 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X2 U656 ( .A(n537), .B(n536), .ZN(n641) );
  NAND2_X1 U657 ( .A1(G953), .A2(G902), .ZN(n612) );
  XOR2_X1 U658 ( .A(KEYINPUT14), .B(n538), .Z(n616) );
  NOR2_X1 U659 ( .A1(n612), .A2(n616), .ZN(n539) );
  XNOR2_X1 U660 ( .A(n539), .B(KEYINPUT105), .ZN(n540) );
  NOR2_X1 U661 ( .A1(G900), .A2(n540), .ZN(n543) );
  INV_X1 U662 ( .A(n616), .ZN(n541) );
  NAND2_X1 U663 ( .A1(G952), .A2(n541), .ZN(n709) );
  NOR2_X1 U664 ( .A1(G953), .A2(n709), .ZN(n542) );
  NOR2_X1 U665 ( .A1(n543), .A2(n542), .ZN(n573) );
  NOR2_X1 U666 ( .A1(n641), .A2(n573), .ZN(n546) );
  NAND2_X1 U667 ( .A1(G221), .A2(n544), .ZN(n545) );
  XOR2_X1 U668 ( .A(KEYINPUT21), .B(n545), .Z(n630) );
  NAND2_X1 U669 ( .A1(n546), .A2(n630), .ZN(n584) );
  XOR2_X1 U670 ( .A(KEYINPUT28), .B(n547), .Z(n554) );
  AND2_X1 U671 ( .A1(G227), .A2(n768), .ZN(n551) );
  INV_X1 U672 ( .A(n595), .ZN(n566) );
  XOR2_X1 U673 ( .A(KEYINPUT74), .B(KEYINPUT18), .Z(n559) );
  XNOR2_X1 U674 ( .A(KEYINPUT17), .B(KEYINPUT88), .ZN(n558) );
  NOR2_X1 U675 ( .A1(n728), .A2(n649), .ZN(n562) );
  NAND2_X1 U676 ( .A1(G210), .A2(n563), .ZN(n561) );
  XNOR2_X1 U677 ( .A(n562), .B(n561), .ZN(n569) );
  NAND2_X1 U678 ( .A1(G214), .A2(n563), .ZN(n697) );
  NAND2_X1 U679 ( .A1(n569), .A2(n697), .ZN(n565) );
  NAND2_X1 U680 ( .A1(n566), .A2(n618), .ZN(n597) );
  NAND2_X1 U681 ( .A1(n597), .A2(KEYINPUT47), .ZN(n567) );
  NAND2_X1 U682 ( .A1(n568), .A2(n567), .ZN(n580) );
  BUF_X1 U683 ( .A(n569), .Z(n609) );
  INV_X1 U684 ( .A(n609), .ZN(n588) );
  INV_X1 U685 ( .A(n582), .ZN(n570) );
  INV_X1 U686 ( .A(n625), .ZN(n576) );
  XOR2_X1 U687 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n572) );
  NAND2_X1 U688 ( .A1(n693), .A2(n697), .ZN(n571) );
  XNOR2_X1 U689 ( .A(n572), .B(n571), .ZN(n575) );
  INV_X1 U690 ( .A(n577), .ZN(n593) );
  NOR2_X1 U691 ( .A1(n592), .A2(n593), .ZN(n578) );
  XNOR2_X1 U692 ( .A(n578), .B(KEYINPUT104), .ZN(n648) );
  XNOR2_X1 U693 ( .A(n675), .B(KEYINPUT80), .ZN(n579) );
  NOR2_X1 U694 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U695 ( .A1(n644), .A2(n585), .ZN(n605) );
  XOR2_X1 U696 ( .A(KEYINPUT36), .B(n586), .Z(n587) );
  INV_X1 U697 ( .A(KEYINPUT39), .ZN(n589) );
  NAND2_X1 U698 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U699 ( .A1(n593), .A2(n592), .ZN(n700) );
  XNOR2_X1 U700 ( .A(n594), .B(KEYINPUT41), .ZN(n719) );
  XOR2_X1 U701 ( .A(KEYINPUT46), .B(KEYINPUT82), .Z(n596) );
  INV_X1 U702 ( .A(n597), .ZN(n677) );
  XOR2_X1 U703 ( .A(KEYINPUT79), .B(n702), .Z(n627) );
  NOR2_X1 U704 ( .A1(KEYINPUT47), .A2(n627), .ZN(n598) );
  NAND2_X1 U705 ( .A1(n677), .A2(n598), .ZN(n599) );
  NOR2_X1 U706 ( .A1(n604), .A2(n603), .ZN(n686) );
  XOR2_X1 U707 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n608) );
  NOR2_X1 U708 ( .A1(n621), .A2(n605), .ZN(n606) );
  NAND2_X1 U709 ( .A1(n606), .A2(n697), .ZN(n607) );
  XNOR2_X1 U710 ( .A(n608), .B(n607), .ZN(n610) );
  NOR2_X1 U711 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U712 ( .A(n611), .B(KEYINPUT107), .ZN(n772) );
  AND2_X1 U713 ( .A1(n768), .A2(G952), .ZN(n614) );
  NOR2_X1 U714 ( .A1(G898), .A2(n612), .ZN(n613) );
  NOR2_X1 U715 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U716 ( .A1(n616), .A2(n615), .ZN(n617) );
  BUF_X1 U717 ( .A(n632), .Z(n622) );
  NOR2_X1 U718 ( .A1(n642), .A2(n645), .ZN(n695) );
  NAND2_X1 U719 ( .A1(n622), .A2(n695), .ZN(n623) );
  XNOR2_X1 U720 ( .A(n623), .B(KEYINPUT31), .ZN(n682) );
  NOR2_X1 U721 ( .A1(n682), .A2(n668), .ZN(n626) );
  XNOR2_X1 U722 ( .A(n626), .B(KEYINPUT95), .ZN(n629) );
  INV_X1 U723 ( .A(n627), .ZN(n628) );
  NAND2_X1 U724 ( .A1(n629), .A2(n628), .ZN(n635) );
  INV_X1 U725 ( .A(n630), .ZN(n688) );
  NOR2_X1 U726 ( .A1(n688), .A2(n700), .ZN(n631) );
  NAND2_X1 U727 ( .A1(n632), .A2(n631), .ZN(n633) );
  INV_X1 U728 ( .A(n641), .ZN(n689) );
  NOR2_X1 U729 ( .A1(n621), .A2(n689), .ZN(n634) );
  NAND2_X1 U730 ( .A1(n639), .A2(n634), .ZN(n666) );
  XNOR2_X1 U731 ( .A(KEYINPUT66), .B(KEYINPUT75), .ZN(n636) );
  XNOR2_X1 U732 ( .A(n636), .B(KEYINPUT32), .ZN(n640) );
  NOR2_X1 U733 ( .A1(n637), .A2(n641), .ZN(n638) );
  INV_X1 U734 ( .A(KEYINPUT2), .ZN(n711) );
  NAND2_X1 U735 ( .A1(KEYINPUT2), .A2(KEYINPUT67), .ZN(n652) );
  XNOR2_X2 U736 ( .A(n653), .B(KEYINPUT65), .ZN(n730) );
  NAND2_X1 U737 ( .A1(n730), .A2(G472), .ZN(n657) );
  XOR2_X1 U738 ( .A(KEYINPUT62), .B(KEYINPUT87), .Z(n654) );
  XNOR2_X1 U739 ( .A(n657), .B(n656), .ZN(n658) );
  NOR2_X2 U740 ( .A1(n658), .A2(n740), .ZN(n660) );
  XNOR2_X1 U741 ( .A(n660), .B(n659), .ZN(G57) );
  NAND2_X1 U742 ( .A1(n738), .A2(G469), .ZN(n664) );
  XNOR2_X1 U743 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n663) );
  XNOR2_X1 U744 ( .A(n661), .B(KEYINPUT57), .ZN(n662) );
  XNOR2_X1 U745 ( .A(G101), .B(n666), .ZN(G3) );
  NAND2_X1 U746 ( .A1(n668), .A2(n679), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n667), .B(G104), .ZN(G6) );
  XOR2_X1 U748 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n670) );
  NAND2_X1 U749 ( .A1(n668), .A2(n681), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n670), .B(n669), .ZN(n672) );
  XOR2_X1 U751 ( .A(G107), .B(KEYINPUT111), .Z(n671) );
  XNOR2_X1 U752 ( .A(n672), .B(n671), .ZN(G9) );
  XOR2_X1 U753 ( .A(G110), .B(n361), .Z(G12) );
  XOR2_X1 U754 ( .A(G128), .B(KEYINPUT29), .Z(n674) );
  NAND2_X1 U755 ( .A1(n681), .A2(n677), .ZN(n673) );
  XNOR2_X1 U756 ( .A(n674), .B(n673), .ZN(G30) );
  XOR2_X1 U757 ( .A(n675), .B(n446), .Z(n676) );
  XNOR2_X1 U758 ( .A(KEYINPUT112), .B(n676), .ZN(G45) );
  NAND2_X1 U759 ( .A1(n677), .A2(n679), .ZN(n678) );
  XNOR2_X1 U760 ( .A(n678), .B(G146), .ZN(G48) );
  NAND2_X1 U761 ( .A1(n682), .A2(n679), .ZN(n680) );
  XNOR2_X1 U762 ( .A(n680), .B(G113), .ZN(G15) );
  NAND2_X1 U763 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U764 ( .A(n683), .B(G116), .ZN(G18) );
  XNOR2_X1 U765 ( .A(G125), .B(n684), .ZN(n685) );
  XNOR2_X1 U766 ( .A(n685), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U767 ( .A(G134), .B(n686), .Z(G36) );
  NAND2_X1 U768 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U769 ( .A(n690), .B(KEYINPUT113), .ZN(n691) );
  XNOR2_X1 U770 ( .A(KEYINPUT49), .B(n691), .ZN(n692) );
  NOR2_X1 U771 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U772 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U773 ( .A1(n700), .A2(n699), .ZN(n705) );
  NOR2_X1 U774 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U775 ( .A(KEYINPUT115), .B(n703), .Z(n704) );
  NOR2_X1 U776 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U777 ( .A1(n706), .A2(n718), .ZN(n707) );
  XOR2_X1 U778 ( .A(KEYINPUT118), .B(n710), .Z(n717) );
  NAND2_X1 U779 ( .A1(n711), .A2(n760), .ZN(n712) );
  XNOR2_X1 U780 ( .A(KEYINPUT81), .B(n712), .ZN(n713) );
  NAND2_X1 U781 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U782 ( .A1(n717), .A2(n716), .ZN(n721) );
  NOR2_X1 U783 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U784 ( .A(n722), .B(KEYINPUT119), .ZN(n723) );
  NOR2_X1 U785 ( .A1(G953), .A2(n723), .ZN(n724) );
  XNOR2_X1 U786 ( .A(KEYINPUT53), .B(n724), .ZN(G75) );
  XOR2_X1 U787 ( .A(KEYINPUT86), .B(KEYINPUT76), .Z(n726) );
  XNOR2_X1 U788 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n725) );
  XNOR2_X1 U789 ( .A(n726), .B(n725), .ZN(n727) );
  NAND2_X1 U790 ( .A1(G210), .A2(n730), .ZN(n729) );
  NAND2_X1 U791 ( .A1(n730), .A2(G475), .ZN(n733) );
  XNOR2_X1 U792 ( .A(n733), .B(n486), .ZN(n735) );
  NAND2_X1 U793 ( .A1(n738), .A2(G478), .ZN(n736) );
  NAND2_X1 U794 ( .A1(G217), .A2(n738), .ZN(n739) );
  XOR2_X1 U795 ( .A(n741), .B(KEYINPUT123), .Z(n742) );
  XNOR2_X1 U796 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U797 ( .A(n744), .B(G101), .ZN(n746) );
  NOR2_X1 U798 ( .A1(n768), .A2(G898), .ZN(n745) );
  NOR2_X1 U799 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U800 ( .A(KEYINPUT124), .B(n747), .ZN(n755) );
  NAND2_X1 U801 ( .A1(n650), .A2(n768), .ZN(n748) );
  XNOR2_X1 U802 ( .A(n748), .B(KEYINPUT122), .ZN(n753) );
  XOR2_X1 U803 ( .A(KEYINPUT61), .B(KEYINPUT121), .Z(n750) );
  NAND2_X1 U804 ( .A1(G224), .A2(G953), .ZN(n749) );
  XNOR2_X1 U805 ( .A(n750), .B(n749), .ZN(n751) );
  NAND2_X1 U806 ( .A1(n751), .A2(G898), .ZN(n752) );
  NAND2_X1 U807 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U808 ( .A(n755), .B(n754), .ZN(G69) );
  XOR2_X1 U809 ( .A(n756), .B(n757), .Z(n758) );
  XNOR2_X1 U810 ( .A(n759), .B(n758), .ZN(n764) );
  INV_X1 U811 ( .A(n764), .ZN(n761) );
  XNOR2_X1 U812 ( .A(n761), .B(n760), .ZN(n762) );
  NOR2_X1 U813 ( .A1(G953), .A2(n762), .ZN(n763) );
  XNOR2_X1 U814 ( .A(KEYINPUT125), .B(n763), .ZN(n771) );
  XNOR2_X1 U815 ( .A(G227), .B(n764), .ZN(n765) );
  NAND2_X1 U816 ( .A1(n765), .A2(G900), .ZN(n766) );
  XOR2_X1 U817 ( .A(KEYINPUT126), .B(n766), .Z(n767) );
  NOR2_X1 U818 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U819 ( .A(KEYINPUT127), .B(n769), .ZN(n770) );
  NAND2_X1 U820 ( .A1(n771), .A2(n770), .ZN(G72) );
  XNOR2_X1 U821 ( .A(G140), .B(n772), .ZN(G42) );
  XNOR2_X1 U822 ( .A(n773), .B(G137), .ZN(G39) );
  XOR2_X1 U823 ( .A(n774), .B(G119), .Z(G21) );
  XOR2_X1 U824 ( .A(n366), .B(G122), .Z(G24) );
  XNOR2_X1 U825 ( .A(G131), .B(n776), .ZN(G33) );
endmodule

