

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(G1384), .A2(G164), .ZN(n772) );
  XNOR2_X2 U553 ( .A(n547), .B(KEYINPUT88), .ZN(G164) );
  NOR2_X1 U554 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  NOR2_X1 U555 ( .A1(n692), .A2(n1012), .ZN(n694) );
  AND2_X1 U556 ( .A1(n807), .A2(n806), .ZN(n809) );
  XNOR2_X2 U557 ( .A(n538), .B(KEYINPUT66), .ZN(n609) );
  XOR2_X1 U558 ( .A(n774), .B(KEYINPUT90), .Z(n519) );
  INV_X1 U559 ( .A(KEYINPUT64), .ZN(n693) );
  XNOR2_X1 U560 ( .A(n694), .B(n693), .ZN(n702) );
  XNOR2_X1 U561 ( .A(KEYINPUT29), .B(KEYINPUT101), .ZN(n716) );
  XNOR2_X1 U562 ( .A(n717), .B(n716), .ZN(n721) );
  INV_X1 U563 ( .A(G2104), .ZN(n541) );
  NOR2_X1 U564 ( .A1(n519), .A2(n805), .ZN(n806) );
  XOR2_X1 U565 ( .A(KEYINPUT0), .B(G543), .Z(n629) );
  INV_X1 U566 ( .A(KEYINPUT106), .ZN(n808) );
  XNOR2_X1 U567 ( .A(KEYINPUT68), .B(n525), .ZN(n649) );
  NOR2_X1 U568 ( .A1(G651), .A2(n629), .ZN(n643) );
  INV_X1 U569 ( .A(KEYINPUT74), .ZN(n535) );
  XNOR2_X1 U570 ( .A(n535), .B(KEYINPUT8), .ZN(n536) );
  XNOR2_X1 U571 ( .A(G168), .B(n536), .ZN(G286) );
  NAND2_X1 U572 ( .A1(n643), .A2(G51), .ZN(n522) );
  XNOR2_X1 U573 ( .A(KEYINPUT67), .B(G651), .ZN(n524) );
  NOR2_X1 U574 ( .A1(G543), .A2(n524), .ZN(n520) );
  XOR2_X1 U575 ( .A(KEYINPUT1), .B(n520), .Z(n645) );
  NAND2_X1 U576 ( .A1(G63), .A2(n645), .ZN(n521) );
  NAND2_X1 U577 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U578 ( .A(KEYINPUT6), .B(n523), .ZN(n532) );
  NOR2_X1 U579 ( .A1(n629), .A2(n524), .ZN(n525) );
  NAND2_X1 U580 ( .A1(n649), .A2(G76), .ZN(n526) );
  XNOR2_X1 U581 ( .A(KEYINPUT72), .B(n526), .ZN(n529) );
  NOR2_X1 U582 ( .A1(G651), .A2(G543), .ZN(n644) );
  NAND2_X1 U583 ( .A1(n644), .A2(G89), .ZN(n527) );
  XNOR2_X1 U584 ( .A(KEYINPUT4), .B(n527), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U586 ( .A(n530), .B(KEYINPUT5), .Z(n531) );
  NOR2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U588 ( .A(KEYINPUT73), .B(n533), .Z(n534) );
  XOR2_X1 U589 ( .A(KEYINPUT7), .B(n534), .Z(G168) );
  XOR2_X2 U590 ( .A(KEYINPUT17), .B(n537), .Z(n887) );
  NAND2_X1 U591 ( .A1(G138), .A2(n887), .ZN(n540) );
  NOR2_X1 U592 ( .A1(n541), .A2(G2105), .ZN(n538) );
  NAND2_X1 U593 ( .A1(G102), .A2(n609), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n546) );
  NAND2_X1 U595 ( .A1(n541), .A2(G2105), .ZN(n542) );
  XNOR2_X2 U596 ( .A(n542), .B(KEYINPUT65), .ZN(n883) );
  NAND2_X1 U597 ( .A1(G126), .A2(n883), .ZN(n544) );
  AND2_X1 U598 ( .A1(G2105), .A2(G2104), .ZN(n884) );
  NAND2_X1 U599 ( .A1(G114), .A2(n884), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n884), .A2(G113), .ZN(n550) );
  NAND2_X1 U603 ( .A1(n609), .A2(G101), .ZN(n548) );
  XOR2_X1 U604 ( .A(KEYINPUT23), .B(n548), .Z(n549) );
  AND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U606 ( .A1(G125), .A2(n883), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G137), .A2(n887), .ZN(n551) );
  AND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n553) );
  AND2_X1 U609 ( .A1(n554), .A2(n553), .ZN(G160) );
  NAND2_X1 U610 ( .A1(n645), .A2(G64), .ZN(n555) );
  XOR2_X1 U611 ( .A(KEYINPUT70), .B(n555), .Z(n562) );
  NAND2_X1 U612 ( .A1(G90), .A2(n644), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G77), .A2(n649), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U615 ( .A(n558), .B(KEYINPUT9), .ZN(n560) );
  NAND2_X1 U616 ( .A1(G52), .A2(n643), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U618 ( .A1(n562), .A2(n561), .ZN(G171) );
  AND2_X1 U619 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U620 ( .A(G57), .ZN(G237) );
  NAND2_X1 U621 ( .A1(G88), .A2(n644), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G75), .A2(n649), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n643), .A2(G50), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G62), .A2(n645), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U628 ( .A(KEYINPUT84), .B(n569), .Z(G303) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U630 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U631 ( .A(G223), .ZN(n825) );
  NAND2_X1 U632 ( .A1(n825), .A2(G567), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  XNOR2_X1 U634 ( .A(KEYINPUT71), .B(KEYINPUT13), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n644), .A2(G81), .ZN(n572) );
  XNOR2_X1 U636 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G68), .A2(n649), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(n576), .B(n575), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G56), .A2(n645), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n577), .Z(n578) );
  NOR2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n643), .A2(G43), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n1012) );
  INV_X1 U645 ( .A(G860), .ZN(n600) );
  OR2_X1 U646 ( .A1(n1012), .A2(n600), .ZN(G153) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  NAND2_X1 U648 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U649 ( .A1(G92), .A2(n644), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G79), .A2(n649), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n643), .A2(G54), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G66), .A2(n645), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U656 ( .A(KEYINPUT15), .B(n588), .Z(n1000) );
  INV_X1 U657 ( .A(n1000), .ZN(n701) );
  INV_X1 U658 ( .A(G868), .ZN(n656) );
  NAND2_X1 U659 ( .A1(n701), .A2(n656), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U661 ( .A1(G78), .A2(n649), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G53), .A2(n643), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n644), .A2(G91), .ZN(n594) );
  NAND2_X1 U665 ( .A1(G65), .A2(n645), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n997) );
  INV_X1 U668 ( .A(n997), .ZN(G299) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n597) );
  XOR2_X1 U670 ( .A(KEYINPUT75), .B(n597), .Z(n599) );
  NOR2_X1 U671 ( .A1(G286), .A2(n656), .ZN(n598) );
  NOR2_X1 U672 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U673 ( .A1(n600), .A2(G559), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n601), .A2(n1000), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U676 ( .A1(G868), .A2(n1012), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n1000), .A2(G868), .ZN(n603) );
  NOR2_X1 U678 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U679 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G123), .A2(n883), .ZN(n606) );
  XNOR2_X1 U681 ( .A(n606), .B(KEYINPUT18), .ZN(n614) );
  NAND2_X1 U682 ( .A1(G111), .A2(n884), .ZN(n608) );
  NAND2_X1 U683 ( .A1(G135), .A2(n887), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n609), .A2(G99), .ZN(n610) );
  XOR2_X1 U686 ( .A(KEYINPUT76), .B(n610), .Z(n611) );
  NOR2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n971) );
  XNOR2_X1 U689 ( .A(n971), .B(G2096), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n615), .B(KEYINPUT77), .ZN(n617) );
  INV_X1 U691 ( .A(G2100), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U693 ( .A1(G559), .A2(n1000), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n618), .B(n1012), .ZN(n664) );
  NOR2_X1 U695 ( .A1(G860), .A2(n664), .ZN(n628) );
  NAND2_X1 U696 ( .A1(n643), .A2(G55), .ZN(n620) );
  NAND2_X1 U697 ( .A1(G67), .A2(n645), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U699 ( .A(KEYINPUT80), .B(n621), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G93), .A2(n644), .ZN(n622) );
  XNOR2_X1 U701 ( .A(KEYINPUT79), .B(n622), .ZN(n623) );
  NOR2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n649), .A2(G80), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n661) );
  XOR2_X1 U705 ( .A(n661), .B(KEYINPUT78), .Z(n627) );
  XNOR2_X1 U706 ( .A(n628), .B(n627), .ZN(G145) );
  NAND2_X1 U707 ( .A1(G49), .A2(n643), .ZN(n631) );
  NAND2_X1 U708 ( .A1(G87), .A2(n629), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U710 ( .A1(n645), .A2(n632), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n633) );
  XOR2_X1 U712 ( .A(KEYINPUT81), .B(n633), .Z(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(G288) );
  NAND2_X1 U714 ( .A1(n643), .A2(G47), .ZN(n637) );
  NAND2_X1 U715 ( .A1(G60), .A2(n645), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U717 ( .A(KEYINPUT69), .B(n638), .ZN(n642) );
  NAND2_X1 U718 ( .A1(G85), .A2(n644), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G72), .A2(n649), .ZN(n639) );
  AND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(G290) );
  NAND2_X1 U722 ( .A1(n643), .A2(G48), .ZN(n654) );
  NAND2_X1 U723 ( .A1(n644), .A2(G86), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G61), .A2(n645), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U726 ( .A(KEYINPUT82), .B(n648), .ZN(n652) );
  NAND2_X1 U727 ( .A1(n649), .A2(G73), .ZN(n650) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(n650), .Z(n651) );
  NOR2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U731 ( .A(KEYINPUT83), .B(n655), .Z(G305) );
  AND2_X1 U732 ( .A1(n656), .A2(n661), .ZN(n657) );
  XNOR2_X1 U733 ( .A(n657), .B(KEYINPUT85), .ZN(n667) );
  XNOR2_X1 U734 ( .A(G288), .B(KEYINPUT19), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n997), .B(G303), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n660), .B(G290), .ZN(n662) );
  XNOR2_X1 U738 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(G305), .ZN(n899) );
  XNOR2_X1 U740 ( .A(n899), .B(n664), .ZN(n665) );
  NAND2_X1 U741 ( .A1(G868), .A2(n665), .ZN(n666) );
  NAND2_X1 U742 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U744 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U747 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U748 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U749 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n673) );
  NAND2_X1 U750 ( .A1(G132), .A2(G82), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n674), .A2(G96), .ZN(n675) );
  NOR2_X1 U753 ( .A1(n675), .A2(G218), .ZN(n676) );
  XNOR2_X1 U754 ( .A(n676), .B(KEYINPUT87), .ZN(n830) );
  NAND2_X1 U755 ( .A1(n830), .A2(G2106), .ZN(n680) );
  NAND2_X1 U756 ( .A1(G120), .A2(G108), .ZN(n677) );
  NOR2_X1 U757 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U758 ( .A1(G69), .A2(n678), .ZN(n831) );
  NAND2_X1 U759 ( .A1(n831), .A2(G567), .ZN(n679) );
  NAND2_X1 U760 ( .A1(n680), .A2(n679), .ZN(n832) );
  NAND2_X1 U761 ( .A1(G483), .A2(G661), .ZN(n681) );
  NOR2_X1 U762 ( .A1(n832), .A2(n681), .ZN(n829) );
  NAND2_X1 U763 ( .A1(n829), .A2(G36), .ZN(G176) );
  AND2_X1 U764 ( .A1(G160), .A2(G40), .ZN(n770) );
  NAND2_X2 U765 ( .A1(n772), .A2(n770), .ZN(n736) );
  NAND2_X1 U766 ( .A1(G8), .A2(n736), .ZN(n766) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n682) );
  XOR2_X1 U768 ( .A(n682), .B(KEYINPUT24), .Z(n683) );
  NOR2_X1 U769 ( .A1(n766), .A2(n683), .ZN(n761) );
  XOR2_X1 U770 ( .A(G1981), .B(G305), .Z(n994) );
  NOR2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n684) );
  XOR2_X1 U772 ( .A(KEYINPUT104), .B(n684), .Z(n1009) );
  NOR2_X1 U773 ( .A1(n766), .A2(n1009), .ZN(n685) );
  NAND2_X1 U774 ( .A1(KEYINPUT33), .A2(n685), .ZN(n686) );
  NAND2_X1 U775 ( .A1(n994), .A2(n686), .ZN(n759) );
  NOR2_X1 U776 ( .A1(G303), .A2(G1971), .ZN(n1018) );
  INV_X1 U777 ( .A(n1009), .ZN(n687) );
  NOR2_X1 U778 ( .A1(n1018), .A2(n687), .ZN(n753) );
  INV_X1 U779 ( .A(n736), .ZN(n688) );
  XNOR2_X1 U780 ( .A(G1996), .B(KEYINPUT98), .ZN(n948) );
  NAND2_X1 U781 ( .A1(n688), .A2(n948), .ZN(n689) );
  XNOR2_X1 U782 ( .A(n689), .B(KEYINPUT26), .ZN(n691) );
  NAND2_X1 U783 ( .A1(n736), .A2(G1341), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n692) );
  OR2_X2 U785 ( .A1(n702), .A2(n701), .ZN(n699) );
  INV_X1 U786 ( .A(G2067), .ZN(n944) );
  NOR2_X1 U787 ( .A1(n736), .A2(n944), .ZN(n695) );
  XNOR2_X1 U788 ( .A(n695), .B(KEYINPUT99), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n736), .A2(G1348), .ZN(n696) );
  NAND2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U792 ( .A(n700), .B(KEYINPUT100), .ZN(n704) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n711) );
  NAND2_X1 U795 ( .A1(G1956), .A2(n736), .ZN(n705) );
  XNOR2_X1 U796 ( .A(KEYINPUT97), .B(n705), .ZN(n709) );
  XOR2_X1 U797 ( .A(KEYINPUT27), .B(KEYINPUT96), .Z(n707) );
  NAND2_X1 U798 ( .A1(n688), .A2(G2072), .ZN(n706) );
  XOR2_X1 U799 ( .A(n707), .B(n706), .Z(n708) );
  NOR2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U801 ( .A1(n997), .A2(n712), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n715) );
  NOR2_X1 U803 ( .A1(n997), .A2(n712), .ZN(n713) );
  XOR2_X1 U804 ( .A(n713), .B(KEYINPUT28), .Z(n714) );
  NAND2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n717) );
  XOR2_X1 U806 ( .A(KEYINPUT25), .B(G2078), .Z(n949) );
  NOR2_X1 U807 ( .A1(n949), .A2(n736), .ZN(n719) );
  NOR2_X1 U808 ( .A1(n688), .A2(G1961), .ZN(n718) );
  NOR2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n727) );
  OR2_X1 U810 ( .A1(G301), .A2(n727), .ZN(n720) );
  NAND2_X1 U811 ( .A1(n721), .A2(n720), .ZN(n745) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n766), .ZN(n732) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n736), .ZN(n731) );
  NOR2_X1 U814 ( .A1(n732), .A2(n731), .ZN(n722) );
  NAND2_X1 U815 ( .A1(G8), .A2(n722), .ZN(n723) );
  XNOR2_X1 U816 ( .A(KEYINPUT30), .B(n723), .ZN(n724) );
  XOR2_X1 U817 ( .A(KEYINPUT102), .B(n724), .Z(n726) );
  INV_X1 U818 ( .A(G168), .ZN(n725) );
  NAND2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n727), .A2(G301), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U822 ( .A(n730), .B(KEYINPUT31), .ZN(n743) );
  AND2_X1 U823 ( .A1(n745), .A2(n743), .ZN(n735) );
  AND2_X1 U824 ( .A1(G8), .A2(n731), .ZN(n733) );
  OR2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n734) );
  OR2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n752) );
  INV_X1 U827 ( .A(G8), .ZN(n742) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n766), .ZN(n738) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U830 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U831 ( .A1(G303), .A2(n739), .ZN(n740) );
  XOR2_X1 U832 ( .A(KEYINPUT103), .B(n740), .Z(n741) );
  OR2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n746) );
  AND2_X1 U834 ( .A1(n743), .A2(n746), .ZN(n744) );
  NAND2_X1 U835 ( .A1(n745), .A2(n744), .ZN(n749) );
  INV_X1 U836 ( .A(n746), .ZN(n747) );
  OR2_X1 U837 ( .A1(n747), .A2(G286), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U839 ( .A(n750), .B(KEYINPUT32), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n764) );
  AND2_X1 U841 ( .A1(n753), .A2(n764), .ZN(n756) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n1010) );
  INV_X1 U843 ( .A(n766), .ZN(n754) );
  NAND2_X1 U844 ( .A1(n1010), .A2(n754), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U846 ( .A1(n757), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n769) );
  NOR2_X1 U849 ( .A1(G303), .A2(G2090), .ZN(n762) );
  XOR2_X1 U850 ( .A(KEYINPUT105), .B(n762), .Z(n763) );
  NAND2_X1 U851 ( .A1(G8), .A2(n763), .ZN(n765) );
  NAND2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n769), .A2(n768), .ZN(n807) );
  INV_X1 U855 ( .A(n770), .ZN(n771) );
  NOR2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n820) );
  XOR2_X1 U857 ( .A(G1986), .B(KEYINPUT89), .Z(n773) );
  XNOR2_X1 U858 ( .A(G290), .B(n773), .ZN(n1008) );
  NAND2_X1 U859 ( .A1(n820), .A2(n1008), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n609), .A2(G105), .ZN(n775) );
  XNOR2_X1 U861 ( .A(n775), .B(KEYINPUT38), .ZN(n782) );
  NAND2_X1 U862 ( .A1(G129), .A2(n883), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G141), .A2(n887), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U865 ( .A1(G117), .A2(n884), .ZN(n778) );
  XNOR2_X1 U866 ( .A(KEYINPUT93), .B(n778), .ZN(n779) );
  NOR2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n782), .A2(n781), .ZN(n867) );
  NAND2_X1 U869 ( .A1(G1996), .A2(n867), .ZN(n783) );
  XNOR2_X1 U870 ( .A(n783), .B(KEYINPUT94), .ZN(n792) );
  NAND2_X1 U871 ( .A1(G119), .A2(n883), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G107), .A2(n884), .ZN(n784) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G131), .A2(n887), .ZN(n787) );
  NAND2_X1 U875 ( .A1(G95), .A2(n609), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U878 ( .A(KEYINPUT92), .B(n790), .Z(n866) );
  NAND2_X1 U879 ( .A1(n866), .A2(G1991), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n812) );
  INV_X1 U881 ( .A(n812), .ZN(n803) );
  XNOR2_X1 U882 ( .A(G2067), .B(KEYINPUT37), .ZN(n793) );
  XOR2_X1 U883 ( .A(n793), .B(KEYINPUT91), .Z(n818) );
  NAND2_X1 U884 ( .A1(G128), .A2(n883), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G116), .A2(n884), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U887 ( .A(n796), .B(KEYINPUT35), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G140), .A2(n887), .ZN(n798) );
  NAND2_X1 U889 ( .A1(G104), .A2(n609), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U891 ( .A(KEYINPUT34), .B(n799), .Z(n800) );
  NAND2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U893 ( .A(n802), .B(KEYINPUT36), .Z(n861) );
  OR2_X1 U894 ( .A1(n818), .A2(n861), .ZN(n816) );
  NAND2_X1 U895 ( .A1(n803), .A2(n816), .ZN(n987) );
  NAND2_X1 U896 ( .A1(n820), .A2(n987), .ZN(n804) );
  XNOR2_X1 U897 ( .A(KEYINPUT95), .B(n804), .ZN(n805) );
  XNOR2_X1 U898 ( .A(n809), .B(n808), .ZN(n823) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n867), .ZN(n969) );
  NOR2_X1 U900 ( .A1(G1991), .A2(n866), .ZN(n974) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n810) );
  XOR2_X1 U902 ( .A(n810), .B(KEYINPUT107), .Z(n811) );
  NOR2_X1 U903 ( .A1(n974), .A2(n811), .ZN(n813) );
  NOR2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U905 ( .A1(n969), .A2(n814), .ZN(n815) );
  XNOR2_X1 U906 ( .A(n815), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U908 ( .A1(n818), .A2(n861), .ZN(n975) );
  NAND2_X1 U909 ( .A1(n819), .A2(n975), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U912 ( .A(n824), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U913 ( .A1(n825), .A2(G2106), .ZN(n826) );
  XOR2_X1 U914 ( .A(KEYINPUT109), .B(n826), .Z(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U916 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n829), .A2(n828), .ZN(G188) );
  NOR2_X1 U919 ( .A1(n831), .A2(n830), .ZN(G325) );
  XOR2_X1 U920 ( .A(KEYINPUT110), .B(G325), .Z(G261) );
  XNOR2_X1 U921 ( .A(G108), .B(KEYINPUT121), .ZN(G238) );
  INV_X1 U923 ( .A(G132), .ZN(G219) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G82), .ZN(G220) );
  INV_X1 U927 ( .A(n832), .ZN(G319) );
  XOR2_X1 U928 ( .A(G2678), .B(KEYINPUT43), .Z(n834) );
  XNOR2_X1 U929 ( .A(KEYINPUT42), .B(KEYINPUT111), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U931 ( .A(KEYINPUT112), .B(G2090), .Z(n836) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2072), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U934 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U935 ( .A(G2096), .B(G2100), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n842) );
  XOR2_X1 U937 ( .A(G2078), .B(G2084), .Z(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1976), .B(G1961), .Z(n844) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1986), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U942 ( .A(G1981), .B(G1971), .Z(n846) );
  XNOR2_X1 U943 ( .A(G1966), .B(G1956), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U946 ( .A(KEYINPUT113), .B(G2474), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U948 ( .A(G1991), .B(KEYINPUT41), .Z(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G112), .A2(n884), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G100), .A2(n609), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n860) );
  NAND2_X1 U953 ( .A1(G136), .A2(n887), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n855), .B(KEYINPUT114), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G124), .A2(n883), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n856), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U958 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U959 ( .A(n861), .B(G164), .Z(n862) );
  XNOR2_X1 U960 ( .A(n862), .B(n971), .ZN(n871) );
  XOR2_X1 U961 ( .A(KEYINPUT46), .B(KEYINPUT118), .Z(n864) );
  XNOR2_X1 U962 ( .A(KEYINPUT119), .B(KEYINPUT48), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U964 ( .A(G160), .B(n865), .ZN(n869) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U967 ( .A(n871), .B(n870), .Z(n882) );
  XNOR2_X1 U968 ( .A(KEYINPUT47), .B(KEYINPUT117), .ZN(n875) );
  NAND2_X1 U969 ( .A1(G127), .A2(n883), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G115), .A2(n884), .ZN(n872) );
  NAND2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n875), .B(n874), .ZN(n880) );
  NAND2_X1 U973 ( .A1(G103), .A2(n609), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n876), .B(KEYINPUT116), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G139), .A2(n887), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n978) );
  XNOR2_X1 U978 ( .A(n978), .B(G162), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n895) );
  NAND2_X1 U980 ( .A1(G130), .A2(n883), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G118), .A2(n884), .ZN(n885) );
  NAND2_X1 U982 ( .A1(n886), .A2(n885), .ZN(n893) );
  NAND2_X1 U983 ( .A1(n887), .A2(G142), .ZN(n888) );
  XOR2_X1 U984 ( .A(KEYINPUT115), .B(n888), .Z(n890) );
  NAND2_X1 U985 ( .A1(G106), .A2(n609), .ZN(n889) );
  NAND2_X1 U986 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U987 ( .A(n891), .B(KEYINPUT45), .Z(n892) );
  NOR2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U989 ( .A(n895), .B(n894), .Z(n896) );
  NOR2_X1 U990 ( .A1(G37), .A2(n896), .ZN(G395) );
  XNOR2_X1 U991 ( .A(G171), .B(n1012), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n897), .B(G286), .ZN(n898) );
  XOR2_X1 U993 ( .A(n898), .B(KEYINPUT120), .Z(n901) );
  XNOR2_X1 U994 ( .A(n1000), .B(n899), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U997 ( .A(G2438), .B(G2435), .Z(n904) );
  XNOR2_X1 U998 ( .A(G2443), .B(G2430), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1000 ( .A(n905), .B(G2454), .Z(n907) );
  XNOR2_X1 U1001 ( .A(G1341), .B(G1348), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1003 ( .A(G2451), .B(G2427), .Z(n909) );
  XNOR2_X1 U1004 ( .A(KEYINPUT108), .B(G2446), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(n911), .B(n910), .Z(n912) );
  NAND2_X1 U1007 ( .A1(G14), .A2(n912), .ZN(n918) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G69), .ZN(G235) );
  INV_X1 U1016 ( .A(n918), .ZN(G401) );
  XOR2_X1 U1017 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n929) );
  XNOR2_X1 U1018 ( .A(KEYINPUT59), .B(G1348), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n919), .B(G4), .ZN(n927) );
  XNOR2_X1 U1020 ( .A(G1956), .B(G20), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(G1341), .B(G19), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(n920), .B(KEYINPUT124), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(G6), .B(G1981), .ZN(n921) );
  NOR2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1025 ( .A(KEYINPUT125), .B(n923), .ZN(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(n929), .B(n928), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(G1966), .B(G21), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(G1961), .B(G5), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n941) );
  XNOR2_X1 U1033 ( .A(G1986), .B(G24), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(G23), .B(G1976), .ZN(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(G1971), .B(KEYINPUT127), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(n936), .B(G22), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(KEYINPUT58), .B(n939), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1041 ( .A(KEYINPUT61), .B(n942), .Z(n943) );
  NOR2_X1 U1042 ( .A1(G16), .A2(n943), .ZN(n967) );
  INV_X1 U1043 ( .A(KEYINPUT55), .ZN(n989) );
  XNOR2_X1 U1044 ( .A(G2090), .B(G35), .ZN(n958) );
  XNOR2_X1 U1045 ( .A(G26), .B(n944), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(n945), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(G1991), .B(G25), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(G33), .B(G2072), .ZN(n946) );
  NOR2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(n948), .B(G32), .ZN(n951) );
  XNOR2_X1 U1051 ( .A(G27), .B(n949), .ZN(n950) );
  NOR2_X1 U1052 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(KEYINPUT53), .B(n956), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1057 ( .A(G2084), .B(G34), .Z(n959) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(n959), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(n989), .B(n962), .ZN(n964) );
  INV_X1 U1061 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n965), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n993) );
  XOR2_X1 U1065 ( .A(G2090), .B(G162), .Z(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1067 ( .A(KEYINPUT51), .B(n970), .Z(n985) );
  XNOR2_X1 U1068 ( .A(G160), .B(G2084), .ZN(n972) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n983) );
  XOR2_X1 U1072 ( .A(G2078), .B(KEYINPUT122), .Z(n977) );
  XNOR2_X1 U1073 ( .A(G164), .B(n977), .ZN(n980) );
  XOR2_X1 U1074 ( .A(G2072), .B(n978), .Z(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1076 ( .A(KEYINPUT50), .B(n981), .Z(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT52), .B(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n991), .A2(G29), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n1022) );
  XOR2_X1 U1084 ( .A(KEYINPUT56), .B(G16), .Z(n1020) );
  XNOR2_X1 U1085 ( .A(G1966), .B(G168), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n996), .B(KEYINPUT57), .ZN(n1006) );
  XNOR2_X1 U1088 ( .A(G171), .B(G1961), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(n997), .B(G1956), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(n1000), .B(G1348), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(G1971), .A2(G303), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1016) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(KEYINPUT123), .B(n1011), .Z(n1014) );
  XNOR2_X1 U1099 ( .A(G1341), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1104 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1105 ( .A(n1023), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
  INV_X1 U1107 ( .A(G303), .ZN(G166) );
endmodule

