//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G217));
  OR4_X1    g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(G567), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(new_n466), .B2(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n465), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n465), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT69), .Z(G160));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT70), .Z(new_n481));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n482));
  INV_X1    g057(.A(G2104), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(KEYINPUT68), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n465), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n481), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  OAI211_X1 g069(.A(G138), .B(new_n465), .C1(new_n467), .C2(new_n468), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n496), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n495), .A2(KEYINPUT4), .B1(new_n473), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n467), .B2(new_n468), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n465), .B2(G114), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n504));
  OR2_X1    g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n502), .A2(new_n504), .A3(new_n505), .A4(G2104), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT72), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n500), .A2(KEYINPUT72), .A3(new_n506), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n498), .B1(new_n508), .B2(new_n509), .ZN(G164));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n516), .A2(KEYINPUT74), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT73), .A3(G50), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n513), .A2(new_n518), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n520), .A2(new_n524), .B1(G88), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n516), .A2(KEYINPUT74), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n517), .A2(new_n527), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n519), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n519), .A2(new_n531), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  INV_X1    g114(.A(G89), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n537), .B(new_n539), .C1(new_n525), .C2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n536), .A2(new_n541), .ZN(G168));
  INV_X1    g117(.A(new_n513), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  INV_X1    g119(.A(G77), .ZN(new_n545));
  INV_X1    g120(.A(G543), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n543), .A2(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT76), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n549));
  OAI221_X1 g124(.A(new_n549), .B1(new_n545), .B2(new_n546), .C1(new_n543), .C2(new_n544), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n548), .A2(G651), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n526), .A2(G90), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n533), .A2(new_n534), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n551), .B(new_n552), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT77), .ZN(G171));
  NAND2_X1  g131(.A1(new_n535), .A2(G43), .ZN(new_n557));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n543), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n515), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n562), .B1(new_n561), .B2(new_n560), .ZN(new_n563));
  XOR2_X1   g138(.A(KEYINPUT79), .B(G81), .Z(new_n564));
  NAND2_X1  g139(.A1(new_n526), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n557), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT80), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  INV_X1    g148(.A(KEYINPUT81), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n522), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n518), .A2(KEYINPUT81), .A3(G53), .A4(G543), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n576), .A2(KEYINPUT9), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n574), .B(new_n579), .C1(new_n522), .C2(new_n575), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n526), .A2(G91), .ZN(new_n581));
  INV_X1    g156(.A(G65), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n511), .B2(new_n512), .ZN(new_n583));
  AND2_X1   g158(.A1(G78), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n578), .A2(new_n580), .A3(new_n581), .A4(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  INV_X1    g162(.A(G168), .ZN(G286));
  NAND2_X1  g163(.A1(new_n526), .A2(G87), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n519), .A2(G49), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n513), .A2(new_n593), .A3(G61), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT83), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n593), .B1(new_n513), .B2(G61), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n526), .A2(G86), .B1(new_n519), .B2(G48), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G305));
  AND2_X1   g176(.A1(new_n535), .A2(G47), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n603), .A2(new_n515), .B1(new_n604), .B2(new_n525), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(new_n526), .A2(G92), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT10), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(new_n515), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n535), .A2(G54), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g191(.A(new_n615), .B1(G171), .B2(G868), .ZN(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G299), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G168), .B2(new_n618), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(G168), .B2(new_n618), .ZN(G280));
  INV_X1    g196(.A(new_n614), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n566), .A2(new_n618), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n614), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g203(.A(new_n471), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n473), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n635));
  INV_X1    g210(.A(G135), .ZN(new_n636));
  INV_X1    g211(.A(G123), .ZN(new_n637));
  OAI221_X1 g212(.A(new_n635), .B1(new_n487), .B2(new_n636), .C1(new_n637), .C2(new_n490), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n633), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT84), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2430), .Z(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n647), .B(new_n651), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(G14), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n653), .ZN(G401));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2084), .B(G2090), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n658), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT87), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT86), .ZN(new_n669));
  INV_X1    g244(.A(new_n662), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n669), .B1(new_n670), .B2(new_n658), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2096), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n667), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n675), .A2(new_n680), .A3(new_n678), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n680), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n683));
  AOI211_X1 g258(.A(new_n679), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT89), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G229));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G22), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G166), .B2(new_n693), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1971), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(KEYINPUT93), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(KEYINPUT93), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n693), .A2(G23), .ZN(new_n699));
  INV_X1    g274(.A(G288), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n693), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT33), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1976), .ZN(new_n703));
  MUX2_X1   g278(.A(G6), .B(G305), .S(G16), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT92), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n697), .A2(new_n698), .A3(new_n703), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G25), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n488), .A2(G131), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n491), .A2(G119), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n465), .A2(G107), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n714), .B(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT90), .Z(new_n719));
  OAI21_X1  g294(.A(new_n713), .B1(new_n719), .B2(new_n712), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  AND2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n693), .A2(G24), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n606), .B2(new_n693), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(G1986), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n726), .A2(G1986), .ZN(new_n728));
  NOR4_X1   g303(.A1(new_n723), .A2(new_n724), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n710), .A2(new_n711), .A3(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT36), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n712), .A2(G35), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G162), .B2(new_n712), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G2090), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT103), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT103), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n693), .A2(G20), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT23), .Z(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G299), .B2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1956), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n736), .A2(new_n737), .A3(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT104), .Z(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n622), .A2(G16), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G4), .B2(G16), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  INV_X1    g322(.A(G2078), .ZN(new_n748));
  NOR2_X1   g323(.A1(G164), .A2(new_n712), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G27), .B2(new_n712), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n567), .A2(G16), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G16), .B2(G19), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT94), .B(G1341), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n751), .B1(new_n748), .B2(new_n750), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n746), .A2(new_n747), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n693), .A2(G21), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G168), .B2(new_n693), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n638), .A2(new_n712), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT100), .Z(new_n762));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(G28), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n712), .B1(new_n763), .B2(G28), .ZN(new_n765));
  AND2_X1   g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NOR2_X1   g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  OAI22_X1  g342(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n753), .A2(new_n754), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n756), .A2(new_n760), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n712), .A2(G32), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n488), .A2(G141), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n491), .A2(G129), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT26), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n777), .A2(new_n778), .B1(G105), .B2(new_n629), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n773), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n772), .B1(new_n781), .B2(new_n712), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT99), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT27), .B(G1996), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(G160), .A2(G29), .ZN(new_n786));
  INV_X1    g361(.A(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n787), .B2(KEYINPUT24), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(KEYINPUT24), .B2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G2084), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR4_X1   g367(.A1(new_n755), .A2(new_n771), .A3(new_n785), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n734), .A2(G2090), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT102), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n712), .A2(G26), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT28), .Z(new_n797));
  OR2_X1    g372(.A1(G104), .A2(G2105), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n798), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT95), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n488), .A2(G140), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n491), .A2(G128), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(KEYINPUT96), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(KEYINPUT96), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n797), .B1(new_n807), .B2(G29), .ZN(new_n808));
  INV_X1    g383(.A(G2067), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n795), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n712), .A2(G33), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(KEYINPUT97), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(KEYINPUT97), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n814), .A2(G2105), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT25), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n488), .B2(G139), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT98), .Z(new_n821));
  OAI21_X1  g396(.A(new_n812), .B1(new_n821), .B2(new_n712), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(G2072), .Z(new_n823));
  INV_X1    g398(.A(KEYINPUT101), .ZN(new_n824));
  OR3_X1    g399(.A1(new_n824), .A2(G5), .A3(G16), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(G5), .B2(G16), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n825), .B(new_n826), .C1(G301), .C2(new_n693), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1961), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n793), .A2(new_n811), .A3(new_n823), .A4(new_n828), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n731), .A2(new_n744), .A3(new_n829), .ZN(G311));
  INV_X1    g405(.A(G311), .ZN(G150));
  NOR2_X1   g406(.A1(new_n614), .A2(new_n623), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n543), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n837), .A2(G651), .B1(new_n526), .B2(G93), .ZN(new_n838));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n553), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT106), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n567), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n566), .A2(new_n840), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n834), .B(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n841), .A2(new_n847), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  AND2_X1   g427(.A1(new_n805), .A2(new_n806), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n500), .A2(new_n506), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n498), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n807), .A2(new_n855), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n857), .A2(new_n781), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n781), .B1(new_n857), .B2(new_n858), .ZN(new_n860));
  OR3_X1    g435(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT108), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT108), .B1(new_n859), .B2(new_n860), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n862), .A3(new_n821), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT109), .ZN(new_n864));
  OR3_X1    g439(.A1(new_n859), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n859), .B2(new_n860), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n820), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n491), .A2(G130), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n465), .A2(G118), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(G142), .B2(new_n488), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(new_n631), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n718), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT110), .ZN(new_n877));
  INV_X1    g452(.A(new_n875), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n863), .A2(new_n867), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G160), .B(new_n638), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT107), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n493), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n868), .A2(KEYINPUT110), .A3(new_n875), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n883), .B1(new_n868), .B2(new_n875), .ZN(new_n886));
  AOI21_X1  g461(.A(G37), .B1(new_n886), .B2(new_n879), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(KEYINPUT111), .B(KEYINPUT40), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(G395));
  INV_X1    g465(.A(new_n844), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n626), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n844), .B1(G559), .B2(new_n614), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n622), .A2(G299), .ZN(new_n894));
  INV_X1    g469(.A(G299), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n614), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(KEYINPUT112), .A3(new_n896), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n614), .A2(KEYINPUT112), .A3(new_n895), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n892), .A2(new_n893), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n894), .A2(new_n896), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n892), .A2(new_n893), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT42), .B1(new_n901), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n892), .A2(new_n893), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n905), .A2(new_n902), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n908), .B(new_n900), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n606), .B(G303), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n700), .B(G305), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n907), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n907), .B2(new_n911), .ZN(new_n917));
  OAI21_X1  g492(.A(G868), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n841), .A2(G868), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(G295));
  INV_X1    g495(.A(KEYINPUT113), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n918), .A2(new_n921), .A3(new_n919), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n918), .B2(new_n919), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(G331));
  NAND2_X1  g499(.A1(G301), .A2(G168), .ZN(new_n925));
  NAND2_X1  g500(.A1(G171), .A2(G286), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n891), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n844), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n910), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n899), .B1(new_n928), .B2(new_n891), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(KEYINPUT114), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT114), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n927), .A2(new_n935), .A3(new_n844), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(new_n914), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n914), .B1(new_n932), .B2(new_n937), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT43), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n934), .A2(new_n929), .A3(new_n936), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n903), .A2(new_n904), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(new_n899), .B2(new_n904), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n943), .A2(new_n945), .B1(new_n930), .B2(new_n933), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n938), .B(new_n939), .C1(new_n946), .C2(new_n914), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n942), .B1(KEYINPUT43), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n940), .ZN(new_n951));
  INV_X1    g526(.A(new_n941), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT43), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n947), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n950), .A2(new_n956), .ZN(G397));
  XNOR2_X1  g532(.A(new_n807), .B(new_n809), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n781), .ZN(new_n959));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n498), .B2(new_n854), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G40), .ZN(new_n964));
  OR3_X1    g539(.A1(new_n472), .A2(new_n476), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n959), .A2(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n963), .A2(G1996), .A3(new_n965), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT46), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n968), .A2(KEYINPUT46), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  INV_X1    g547(.A(G1996), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n780), .B(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n958), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n719), .A3(new_n722), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(G2067), .B2(new_n807), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n966), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n718), .B(new_n722), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n966), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n982));
  INV_X1    g557(.A(G1986), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n606), .A2(new_n983), .A3(new_n966), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT48), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n972), .B(new_n978), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT127), .Z(new_n989));
  XNOR2_X1  g564(.A(new_n606), .B(new_n983), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n966), .B1(new_n980), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  NOR2_X1   g567(.A1(G168), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT51), .B1(new_n993), .B2(KEYINPUT121), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n472), .A2(new_n476), .A3(new_n964), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n963), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT116), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n963), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  NOR2_X1   g574(.A1(G164), .A2(G1384), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT45), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n995), .B1(new_n961), .B2(KEYINPUT50), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1002), .A2(new_n759), .B1(new_n1006), .B2(new_n791), .ZN(new_n1007));
  AOI211_X1 g582(.A(new_n992), .B(new_n994), .C1(G168), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n993), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1009), .B(new_n994), .C1(new_n1007), .C2(new_n992), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  OAI22_X1  g586(.A1(new_n1008), .A2(new_n1011), .B1(new_n1009), .B2(new_n1007), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G305), .A2(G1981), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n599), .A2(new_n1014), .A3(new_n600), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1013), .B(new_n1015), .C1(KEYINPUT115), .C2(KEYINPUT49), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n965), .A2(new_n961), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(new_n992), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n700), .A2(G1976), .ZN(new_n1023));
  INV_X1    g598(.A(G1976), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT52), .B1(G288), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n473), .A2(new_n497), .ZN(new_n1027));
  AOI211_X1 g602(.A(new_n496), .B(G2105), .C1(new_n484), .C2(new_n485), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT4), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n854), .ZN(new_n1031));
  AOI21_X1  g606(.A(G1384), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n995), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1023), .A2(new_n1033), .A3(G8), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1022), .A2(new_n1026), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1971), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n995), .B1(new_n961), .B2(new_n962), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n500), .A2(KEYINPUT72), .A3(new_n506), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1030), .B1(new_n1040), .B2(new_n507), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT45), .B1(new_n1041), .B2(new_n960), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1041), .A2(new_n1003), .A3(new_n960), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n961), .A2(KEYINPUT50), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n995), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(G2090), .ZN(new_n1048));
  OAI21_X1  g623(.A(G8), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G303), .A2(G8), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT55), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1005), .ZN(new_n1053));
  INV_X1    g628(.A(G2090), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1053), .B(new_n1054), .C1(new_n1003), .C2(new_n1000), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n992), .B1(new_n1055), .B2(new_n1043), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1050), .B(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1037), .A2(new_n1052), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1036), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(KEYINPUT123), .A3(new_n1052), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n1002), .B2(G2078), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1001), .A2(new_n999), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(KEYINPUT122), .A3(new_n748), .A4(new_n997), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1069), .A3(KEYINPUT53), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n748), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1053), .B1(new_n1003), .B2(new_n1000), .ZN(new_n1074));
  INV_X1    g649(.A(G1961), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1072), .A2(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1070), .A2(G301), .A3(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT53), .B(new_n748), .C1(new_n961), .C2(new_n962), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n996), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT124), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1080), .A2(KEYINPUT124), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT54), .B(new_n1077), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n1085));
  AOI21_X1  g660(.A(G301), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1080), .A2(G171), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1012), .A2(new_n1065), .A3(new_n1084), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n965), .B1(KEYINPUT45), .B2(new_n1032), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n962), .B1(G164), .B2(G1384), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n973), .A3(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT58), .B(G1341), .Z(new_n1094));
  NAND2_X1  g669(.A1(new_n1033), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1090), .B1(new_n1096), .B2(new_n567), .ZN(new_n1097));
  AOI211_X1 g672(.A(KEYINPUT59), .B(new_n566), .C1(new_n1093), .C2(new_n1095), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1071), .A2(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n895), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1102), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G299), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n1107));
  INV_X1    g682(.A(G1956), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1047), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1107), .B1(new_n1047), .B2(new_n1108), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1101), .B(new_n1106), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1091), .A2(new_n1100), .A3(new_n1092), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1047), .A2(new_n1108), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT117), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1047), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1111), .B1(new_n1116), .B2(new_n1106), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1099), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1112), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1118), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1101), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1121), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1124), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1119), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1119), .B(KEYINPUT120), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1074), .A2(new_n747), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1020), .A2(new_n809), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(KEYINPUT60), .A3(new_n614), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n622), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1137), .A2(new_n1139), .B1(new_n1138), .B2(new_n1135), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1131), .A2(new_n1132), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1126), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1136), .A2(new_n614), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1111), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1089), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n1147));
  AOI21_X1  g722(.A(G1966), .B1(new_n1068), .B2(new_n997), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1074), .A2(G2084), .ZN(new_n1149));
  OAI211_X1 g724(.A(G8), .B(G168), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1147), .B1(new_n1060), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1056), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1147), .B1(new_n1152), .B2(new_n1051), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n1063), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1151), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1059), .A2(new_n1036), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1022), .A2(new_n1024), .A3(new_n700), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1015), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1021), .B2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n993), .A2(KEYINPUT121), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1007), .A2(new_n992), .ZN(new_n1163));
  OAI211_X1 g738(.A(KEYINPUT51), .B(new_n1162), .C1(new_n1163), .C2(new_n993), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1161), .B1(new_n1164), .B2(new_n1010), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1065), .B(new_n1086), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1160), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g744(.A(KEYINPUT125), .B(new_n991), .C1(new_n1146), .C2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1062), .A2(new_n1064), .A3(new_n1086), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1012), .B2(KEYINPUT62), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1172), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1145), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1140), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1178), .B2(new_n1132), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1176), .B1(new_n1179), .B2(new_n1089), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT125), .B1(new_n1180), .B2(new_n991), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n989), .B1(new_n1171), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g757(.A1(G401), .A2(G227), .A3(new_n463), .ZN(new_n1184));
  NOR2_X1   g758(.A1(G229), .A2(new_n1184), .ZN(new_n1185));
  AND3_X1   g759(.A1(new_n1185), .A2(new_n948), .A3(new_n888), .ZN(G308));
  NAND3_X1  g760(.A1(new_n1185), .A2(new_n948), .A3(new_n888), .ZN(G225));
endmodule


