

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(G651), .A2(n633), .ZN(n655) );
  NAND2_X1 U552 ( .A1(G8), .A2(n746), .ZN(n779) );
  XOR2_X1 U553 ( .A(n585), .B(KEYINPUT14), .Z(n515) );
  NAND2_X2 U554 ( .A1(n782), .A2(n698), .ZN(n730) );
  NOR2_X1 U555 ( .A1(n742), .A2(n741), .ZN(n743) );
  AND2_X2 U556 ( .A1(n541), .A2(G2104), .ZN(n866) );
  NOR2_X2 U557 ( .A1(n696), .A2(G1384), .ZN(n782) );
  NOR2_X1 U558 ( .A1(n730), .A2(n918), .ZN(n700) );
  NAND2_X1 U559 ( .A1(n752), .A2(G8), .ZN(n754) );
  INV_X1 U560 ( .A(KEYINPUT32), .ZN(n753) );
  NOR2_X1 U561 ( .A1(G1966), .A2(n779), .ZN(n760) );
  XOR2_X1 U562 ( .A(KEYINPUT13), .B(n582), .Z(n583) );
  INV_X1 U563 ( .A(G2105), .ZN(n541) );
  INV_X1 U564 ( .A(n723), .ZN(n724) );
  INV_X1 U565 ( .A(KEYINPUT28), .ZN(n718) );
  NOR2_X1 U566 ( .A1(n762), .A2(n761), .ZN(n771) );
  XNOR2_X1 U567 ( .A(n754), .B(n753), .ZN(n762) );
  XNOR2_X1 U568 ( .A(n536), .B(n535), .ZN(n546) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n535) );
  XNOR2_X1 U570 ( .A(n534), .B(KEYINPUT64), .ZN(n536) );
  INV_X1 U571 ( .A(KEYINPUT17), .ZN(n534) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n654) );
  NOR2_X2 U573 ( .A1(n633), .A2(n526), .ZN(n658) );
  XNOR2_X1 U574 ( .A(n538), .B(n537), .ZN(n539) );
  INV_X1 U575 ( .A(KEYINPUT23), .ZN(n537) );
  NOR2_X2 U576 ( .A1(G2104), .A2(n541), .ZN(n871) );
  NAND2_X1 U577 ( .A1(n586), .A2(n515), .ZN(n989) );
  NOR2_X1 U578 ( .A1(n583), .A2(n516), .ZN(n586) );
  XOR2_X1 U579 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  BUF_X1 U580 ( .A(n697), .Z(G160) );
  XNOR2_X2 U581 ( .A(n730), .B(KEYINPUT93), .ZN(n723) );
  AND2_X1 U582 ( .A1(n655), .A2(G43), .ZN(n516) );
  AND2_X1 U583 ( .A1(n817), .A2(n812), .ZN(n517) );
  AND2_X1 U584 ( .A1(n781), .A2(n780), .ZN(n518) );
  NAND2_X1 U585 ( .A1(n774), .A2(n779), .ZN(n519) );
  INV_X1 U586 ( .A(KEYINPUT26), .ZN(n699) );
  NOR2_X1 U587 ( .A1(n733), .A2(n760), .ZN(n734) );
  INV_X1 U588 ( .A(G168), .ZN(n735) );
  INV_X1 U589 ( .A(KEYINPUT92), .ZN(n731) );
  BUF_X1 U590 ( .A(n730), .Z(n746) );
  AND2_X1 U591 ( .A1(n825), .A2(n517), .ZN(n813) );
  INV_X1 U592 ( .A(KEYINPUT103), .ZN(n815) );
  BUF_X1 U593 ( .A(n546), .Z(n867) );
  NAND2_X1 U594 ( .A1(G89), .A2(n654), .ZN(n520) );
  XNOR2_X1 U595 ( .A(n520), .B(KEYINPUT76), .ZN(n521) );
  XNOR2_X1 U596 ( .A(n521), .B(KEYINPUT4), .ZN(n524) );
  XNOR2_X1 U597 ( .A(G543), .B(KEYINPUT0), .ZN(n522) );
  XNOR2_X1 U598 ( .A(n522), .B(KEYINPUT65), .ZN(n633) );
  INV_X1 U599 ( .A(G651), .ZN(n526) );
  NAND2_X1 U600 ( .A1(G76), .A2(n658), .ZN(n523) );
  NAND2_X1 U601 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U602 ( .A(n525), .B(KEYINPUT5), .ZN(n532) );
  NOR2_X1 U603 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X2 U604 ( .A(KEYINPUT1), .B(n527), .Z(n662) );
  NAND2_X1 U605 ( .A1(G63), .A2(n662), .ZN(n529) );
  NAND2_X1 U606 ( .A1(G51), .A2(n655), .ZN(n528) );
  NAND2_X1 U607 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U608 ( .A(KEYINPUT6), .B(n530), .Z(n531) );
  NAND2_X1 U609 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U610 ( .A(n533), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U611 ( .A1(G137), .A2(n546), .ZN(n540) );
  NAND2_X1 U612 ( .A1(G101), .A2(n866), .ZN(n538) );
  NAND2_X1 U613 ( .A1(n540), .A2(n539), .ZN(n545) );
  NAND2_X1 U614 ( .A1(G125), .A2(n871), .ZN(n543) );
  AND2_X1 U615 ( .A1(G2104), .A2(G2105), .ZN(n872) );
  NAND2_X1 U616 ( .A1(G113), .A2(n872), .ZN(n542) );
  NAND2_X1 U617 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U618 ( .A1(n545), .A2(n544), .ZN(n697) );
  NAND2_X1 U619 ( .A1(n546), .A2(G138), .ZN(n548) );
  NAND2_X1 U620 ( .A1(n866), .A2(G102), .ZN(n547) );
  NAND2_X1 U621 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U622 ( .A(n549), .B(KEYINPUT86), .ZN(n553) );
  NAND2_X1 U623 ( .A1(G126), .A2(n871), .ZN(n551) );
  NAND2_X1 U624 ( .A1(G114), .A2(n872), .ZN(n550) );
  NAND2_X1 U625 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U626 ( .A1(n553), .A2(n552), .ZN(n696) );
  BUF_X1 U627 ( .A(n696), .Z(G164) );
  XOR2_X1 U628 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n556) );
  XNOR2_X1 U629 ( .A(G1341), .B(G1348), .ZN(n555) );
  XNOR2_X1 U630 ( .A(n556), .B(n555), .ZN(n566) );
  XOR2_X1 U631 ( .A(G2446), .B(G2435), .Z(n558) );
  XNOR2_X1 U632 ( .A(G2430), .B(KEYINPUT108), .ZN(n557) );
  XNOR2_X1 U633 ( .A(n558), .B(n557), .ZN(n562) );
  XOR2_X1 U634 ( .A(G2438), .B(KEYINPUT107), .Z(n560) );
  XNOR2_X1 U635 ( .A(G2427), .B(G2454), .ZN(n559) );
  XNOR2_X1 U636 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U637 ( .A(n562), .B(n561), .Z(n564) );
  XNOR2_X1 U638 ( .A(G2443), .B(G2451), .ZN(n563) );
  XNOR2_X1 U639 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U640 ( .A(n566), .B(n565), .ZN(n567) );
  AND2_X1 U641 ( .A1(n567), .A2(G14), .ZN(G401) );
  AND2_X1 U642 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U643 ( .A(G57), .ZN(G237) );
  INV_X1 U644 ( .A(G132), .ZN(G219) );
  NAND2_X1 U645 ( .A1(n658), .A2(G77), .ZN(n568) );
  XNOR2_X1 U646 ( .A(n568), .B(KEYINPUT68), .ZN(n570) );
  NAND2_X1 U647 ( .A1(G90), .A2(n654), .ZN(n569) );
  NAND2_X1 U648 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U649 ( .A(n571), .B(KEYINPUT9), .ZN(n573) );
  NAND2_X1 U650 ( .A1(G52), .A2(n655), .ZN(n572) );
  NAND2_X1 U651 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U652 ( .A1(G64), .A2(n662), .ZN(n574) );
  XNOR2_X1 U653 ( .A(KEYINPUT67), .B(n574), .ZN(n575) );
  NOR2_X1 U654 ( .A1(n576), .A2(n575), .ZN(G171) );
  NAND2_X1 U655 ( .A1(G7), .A2(G661), .ZN(n577) );
  XNOR2_X1 U656 ( .A(n577), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U657 ( .A(G223), .ZN(n834) );
  NAND2_X1 U658 ( .A1(n834), .A2(G567), .ZN(n578) );
  XOR2_X1 U659 ( .A(KEYINPUT11), .B(n578), .Z(G234) );
  XOR2_X1 U660 ( .A(G860), .B(KEYINPUT72), .Z(n608) );
  NAND2_X1 U661 ( .A1(n654), .A2(G81), .ZN(n579) );
  XNOR2_X1 U662 ( .A(n579), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U663 ( .A1(G68), .A2(n658), .ZN(n580) );
  NAND2_X1 U664 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U665 ( .A1(G56), .A2(n662), .ZN(n584) );
  XNOR2_X1 U666 ( .A(n584), .B(KEYINPUT71), .ZN(n585) );
  OR2_X1 U667 ( .A1(n608), .A2(n989), .ZN(G153) );
  INV_X1 U668 ( .A(G868), .ZN(n673) );
  NOR2_X1 U669 ( .A1(n673), .A2(G171), .ZN(n587) );
  XNOR2_X1 U670 ( .A(n587), .B(KEYINPUT73), .ZN(n598) );
  NAND2_X1 U671 ( .A1(G92), .A2(n654), .ZN(n588) );
  XNOR2_X1 U672 ( .A(n588), .B(KEYINPUT74), .ZN(n595) );
  NAND2_X1 U673 ( .A1(G66), .A2(n662), .ZN(n590) );
  NAND2_X1 U674 ( .A1(G54), .A2(n655), .ZN(n589) );
  NAND2_X1 U675 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U676 ( .A1(G79), .A2(n658), .ZN(n591) );
  XNOR2_X1 U677 ( .A(KEYINPUT75), .B(n591), .ZN(n592) );
  NOR2_X1 U678 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U679 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X2 U680 ( .A(KEYINPUT15), .B(n596), .ZN(n1001) );
  OR2_X1 U681 ( .A1(G868), .A2(n1001), .ZN(n597) );
  NAND2_X1 U682 ( .A1(n598), .A2(n597), .ZN(G284) );
  NAND2_X1 U683 ( .A1(G65), .A2(n662), .ZN(n600) );
  NAND2_X1 U684 ( .A1(G53), .A2(n655), .ZN(n599) );
  NAND2_X1 U685 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U686 ( .A1(G78), .A2(n658), .ZN(n602) );
  NAND2_X1 U687 ( .A1(G91), .A2(n654), .ZN(n601) );
  NAND2_X1 U688 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U689 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U690 ( .A(n605), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U691 ( .A1(G286), .A2(G868), .ZN(n607) );
  NAND2_X1 U692 ( .A1(G299), .A2(n673), .ZN(n606) );
  NAND2_X1 U693 ( .A1(n607), .A2(n606), .ZN(G297) );
  NAND2_X1 U694 ( .A1(n608), .A2(G559), .ZN(n609) );
  NAND2_X1 U695 ( .A1(n609), .A2(n1001), .ZN(n610) );
  XNOR2_X1 U696 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U697 ( .A1(G559), .A2(n673), .ZN(n611) );
  NAND2_X1 U698 ( .A1(n1001), .A2(n611), .ZN(n612) );
  XNOR2_X1 U699 ( .A(n612), .B(KEYINPUT77), .ZN(n614) );
  NOR2_X1 U700 ( .A1(n989), .A2(G868), .ZN(n613) );
  NOR2_X1 U701 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U702 ( .A1(G99), .A2(n866), .ZN(n616) );
  NAND2_X1 U703 ( .A1(G111), .A2(n872), .ZN(n615) );
  NAND2_X1 U704 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U705 ( .A1(n871), .A2(G123), .ZN(n617) );
  XOR2_X1 U706 ( .A(KEYINPUT18), .B(n617), .Z(n618) );
  NOR2_X1 U707 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U708 ( .A1(G135), .A2(n867), .ZN(n620) );
  NAND2_X1 U709 ( .A1(n621), .A2(n620), .ZN(n971) );
  XNOR2_X1 U710 ( .A(G2096), .B(n971), .ZN(n622) );
  NOR2_X1 U711 ( .A1(G2100), .A2(n622), .ZN(n623) );
  XOR2_X1 U712 ( .A(KEYINPUT78), .B(n623), .Z(G156) );
  NAND2_X1 U713 ( .A1(n1001), .A2(G559), .ZN(n671) );
  XNOR2_X1 U714 ( .A(n989), .B(n671), .ZN(n624) );
  NOR2_X1 U715 ( .A1(n624), .A2(G860), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n654), .A2(G93), .ZN(n627) );
  NAND2_X1 U717 ( .A1(G80), .A2(n658), .ZN(n625) );
  XOR2_X1 U718 ( .A(KEYINPUT79), .B(n625), .Z(n626) );
  NAND2_X1 U719 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U720 ( .A1(G67), .A2(n662), .ZN(n629) );
  NAND2_X1 U721 ( .A1(G55), .A2(n655), .ZN(n628) );
  NAND2_X1 U722 ( .A1(n629), .A2(n628), .ZN(n630) );
  OR2_X1 U723 ( .A1(n631), .A2(n630), .ZN(n674) );
  XOR2_X1 U724 ( .A(n632), .B(n674), .Z(G145) );
  NAND2_X1 U725 ( .A1(G49), .A2(n655), .ZN(n635) );
  NAND2_X1 U726 ( .A1(G87), .A2(n633), .ZN(n634) );
  NAND2_X1 U727 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U728 ( .A1(n662), .A2(n636), .ZN(n638) );
  NAND2_X1 U729 ( .A1(G651), .A2(G74), .ZN(n637) );
  NAND2_X1 U730 ( .A1(n638), .A2(n637), .ZN(G288) );
  NAND2_X1 U731 ( .A1(G75), .A2(n658), .ZN(n640) );
  NAND2_X1 U732 ( .A1(G88), .A2(n654), .ZN(n639) );
  NAND2_X1 U733 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U734 ( .A1(G62), .A2(n662), .ZN(n641) );
  XNOR2_X1 U735 ( .A(KEYINPUT81), .B(n641), .ZN(n642) );
  NOR2_X1 U736 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U737 ( .A1(n655), .A2(G50), .ZN(n644) );
  NAND2_X1 U738 ( .A1(n645), .A2(n644), .ZN(G303) );
  INV_X1 U739 ( .A(G303), .ZN(G166) );
  XOR2_X1 U740 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n647) );
  NAND2_X1 U741 ( .A1(G73), .A2(n658), .ZN(n646) );
  XNOR2_X1 U742 ( .A(n647), .B(n646), .ZN(n651) );
  NAND2_X1 U743 ( .A1(G86), .A2(n654), .ZN(n649) );
  NAND2_X1 U744 ( .A1(G61), .A2(n662), .ZN(n648) );
  NAND2_X1 U745 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U746 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U747 ( .A1(n655), .A2(G48), .ZN(n652) );
  NAND2_X1 U748 ( .A1(n653), .A2(n652), .ZN(G305) );
  NAND2_X1 U749 ( .A1(G85), .A2(n654), .ZN(n657) );
  NAND2_X1 U750 ( .A1(G47), .A2(n655), .ZN(n656) );
  NAND2_X1 U751 ( .A1(n657), .A2(n656), .ZN(n661) );
  NAND2_X1 U752 ( .A1(G72), .A2(n658), .ZN(n659) );
  XOR2_X1 U753 ( .A(KEYINPUT66), .B(n659), .Z(n660) );
  NOR2_X1 U754 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U755 ( .A1(n662), .A2(G60), .ZN(n663) );
  NAND2_X1 U756 ( .A1(n664), .A2(n663), .ZN(G290) );
  XNOR2_X1 U757 ( .A(KEYINPUT19), .B(G299), .ZN(n665) );
  XNOR2_X1 U758 ( .A(n665), .B(G288), .ZN(n668) );
  XNOR2_X1 U759 ( .A(G166), .B(n989), .ZN(n666) );
  XNOR2_X1 U760 ( .A(n666), .B(G305), .ZN(n667) );
  XNOR2_X1 U761 ( .A(n668), .B(n667), .ZN(n670) );
  XOR2_X1 U762 ( .A(G290), .B(n674), .Z(n669) );
  XNOR2_X1 U763 ( .A(n670), .B(n669), .ZN(n886) );
  XOR2_X1 U764 ( .A(n886), .B(n671), .Z(n672) );
  NAND2_X1 U765 ( .A1(G868), .A2(n672), .ZN(n676) );
  NAND2_X1 U766 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U767 ( .A1(n676), .A2(n675), .ZN(G295) );
  XNOR2_X1 U768 ( .A(KEYINPUT20), .B(KEYINPUT83), .ZN(n679) );
  NAND2_X1 U769 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XNOR2_X1 U770 ( .A(n677), .B(KEYINPUT82), .ZN(n678) );
  XNOR2_X1 U771 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U772 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U773 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U774 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U775 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U776 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U777 ( .A1(G220), .A2(G219), .ZN(n683) );
  XOR2_X1 U778 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U779 ( .A1(G218), .A2(n684), .ZN(n685) );
  XNOR2_X1 U780 ( .A(KEYINPUT84), .B(n685), .ZN(n686) );
  NAND2_X1 U781 ( .A1(n686), .A2(G96), .ZN(n841) );
  NAND2_X1 U782 ( .A1(G2106), .A2(n841), .ZN(n687) );
  XOR2_X1 U783 ( .A(KEYINPUT85), .B(n687), .Z(n691) );
  NAND2_X1 U784 ( .A1(G69), .A2(G120), .ZN(n688) );
  NOR2_X1 U785 ( .A1(G237), .A2(n688), .ZN(n689) );
  NAND2_X1 U786 ( .A1(G108), .A2(n689), .ZN(n840) );
  NAND2_X1 U787 ( .A1(G567), .A2(n840), .ZN(n690) );
  NAND2_X1 U788 ( .A1(n691), .A2(n690), .ZN(n890) );
  NAND2_X1 U789 ( .A1(G661), .A2(G483), .ZN(n692) );
  NOR2_X1 U790 ( .A1(n890), .A2(n692), .ZN(n839) );
  NAND2_X1 U791 ( .A1(n839), .A2(G36), .ZN(G176) );
  INV_X1 U792 ( .A(G171), .ZN(G301) );
  NOR2_X1 U793 ( .A1(G2090), .A2(G303), .ZN(n693) );
  XOR2_X1 U794 ( .A(KEYINPUT101), .B(n693), .Z(n694) );
  NAND2_X1 U795 ( .A1(G8), .A2(n694), .ZN(n695) );
  XNOR2_X1 U796 ( .A(KEYINPUT102), .B(n695), .ZN(n773) );
  NAND2_X1 U797 ( .A1(n697), .A2(G40), .ZN(n783) );
  INV_X1 U798 ( .A(n783), .ZN(n698) );
  INV_X1 U799 ( .A(G1996), .ZN(n918) );
  XNOR2_X1 U800 ( .A(n700), .B(n699), .ZN(n702) );
  NAND2_X1 U801 ( .A1(n746), .A2(G1341), .ZN(n701) );
  NAND2_X1 U802 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U803 ( .A1(n703), .A2(n989), .ZN(n709) );
  NAND2_X1 U804 ( .A1(n1001), .A2(n709), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n723), .A2(G2067), .ZN(n705) );
  NAND2_X1 U806 ( .A1(G1348), .A2(n746), .ZN(n704) );
  NAND2_X1 U807 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U808 ( .A(n706), .B(KEYINPUT94), .ZN(n707) );
  NAND2_X1 U809 ( .A1(n708), .A2(n707), .ZN(n711) );
  OR2_X1 U810 ( .A1(n709), .A2(n1001), .ZN(n710) );
  NAND2_X1 U811 ( .A1(n711), .A2(n710), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n723), .A2(G2072), .ZN(n712) );
  XNOR2_X1 U813 ( .A(n712), .B(KEYINPUT27), .ZN(n714) );
  INV_X1 U814 ( .A(G1956), .ZN(n938) );
  NOR2_X1 U815 ( .A1(n938), .A2(n723), .ZN(n713) );
  NOR2_X1 U816 ( .A1(n714), .A2(n713), .ZN(n717) );
  INV_X1 U817 ( .A(G299), .ZN(n1000) );
  NAND2_X1 U818 ( .A1(n717), .A2(n1000), .ZN(n715) );
  NAND2_X1 U819 ( .A1(n716), .A2(n715), .ZN(n721) );
  NOR2_X1 U820 ( .A1(n717), .A2(n1000), .ZN(n719) );
  XNOR2_X1 U821 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U822 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U823 ( .A(n722), .B(KEYINPUT29), .ZN(n729) );
  XOR2_X1 U824 ( .A(G2078), .B(KEYINPUT25), .Z(n925) );
  NOR2_X1 U825 ( .A1(n925), .A2(n724), .ZN(n727) );
  INV_X1 U826 ( .A(n746), .ZN(n725) );
  NOR2_X1 U827 ( .A1(n725), .A2(G1961), .ZN(n726) );
  NOR2_X1 U828 ( .A1(n727), .A2(n726), .ZN(n737) );
  NOR2_X1 U829 ( .A1(G301), .A2(n737), .ZN(n728) );
  NOR2_X1 U830 ( .A1(n729), .A2(n728), .ZN(n742) );
  NOR2_X1 U831 ( .A1(n730), .A2(G2084), .ZN(n732) );
  XNOR2_X1 U832 ( .A(n732), .B(n731), .ZN(n756) );
  NAND2_X1 U833 ( .A1(G8), .A2(n756), .ZN(n733) );
  XNOR2_X1 U834 ( .A(n734), .B(KEYINPUT30), .ZN(n736) );
  AND2_X1 U835 ( .A1(n736), .A2(n735), .ZN(n739) );
  AND2_X1 U836 ( .A1(G301), .A2(n737), .ZN(n738) );
  NOR2_X1 U837 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U838 ( .A(n740), .B(KEYINPUT31), .ZN(n741) );
  XNOR2_X1 U839 ( .A(n743), .B(KEYINPUT95), .ZN(n755) );
  NAND2_X1 U840 ( .A1(n755), .A2(G286), .ZN(n744) );
  XNOR2_X1 U841 ( .A(n744), .B(KEYINPUT96), .ZN(n751) );
  NOR2_X1 U842 ( .A1(G1971), .A2(n779), .ZN(n745) );
  XNOR2_X1 U843 ( .A(KEYINPUT97), .B(n745), .ZN(n749) );
  NOR2_X1 U844 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U845 ( .A1(G166), .A2(n747), .ZN(n748) );
  NAND2_X1 U846 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U847 ( .A1(n751), .A2(n750), .ZN(n752) );
  INV_X1 U848 ( .A(n756), .ZN(n757) );
  NAND2_X1 U849 ( .A1(G8), .A2(n757), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n755), .A2(n758), .ZN(n759) );
  NOR2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n994) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n992) );
  XNOR2_X1 U854 ( .A(KEYINPUT98), .B(n992), .ZN(n763) );
  NOR2_X1 U855 ( .A1(n994), .A2(n763), .ZN(n764) );
  NOR2_X1 U856 ( .A1(n779), .A2(n764), .ZN(n765) );
  NOR2_X1 U857 ( .A1(n771), .A2(n765), .ZN(n767) );
  NAND2_X1 U858 ( .A1(G288), .A2(G1976), .ZN(n766) );
  XNOR2_X1 U859 ( .A(n766), .B(KEYINPUT99), .ZN(n1005) );
  NOR2_X1 U860 ( .A1(n767), .A2(n1005), .ZN(n768) );
  NOR2_X1 U861 ( .A1(n768), .A2(KEYINPUT33), .ZN(n770) );
  XNOR2_X1 U862 ( .A(KEYINPUT100), .B(G1981), .ZN(n769) );
  XNOR2_X1 U863 ( .A(n769), .B(G305), .ZN(n1009) );
  NOR2_X1 U864 ( .A1(n770), .A2(n1009), .ZN(n775) );
  NOR2_X1 U865 ( .A1(n775), .A2(n771), .ZN(n772) );
  NAND2_X1 U866 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U867 ( .A1(n994), .A2(KEYINPUT33), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n775), .A2(n776), .ZN(n781) );
  NOR2_X1 U869 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XOR2_X1 U870 ( .A(n777), .B(KEYINPUT24), .Z(n778) );
  OR2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n519), .A2(n518), .ZN(n814) );
  NOR2_X1 U873 ( .A1(n782), .A2(n783), .ZN(n829) );
  NAND2_X1 U874 ( .A1(n866), .A2(G104), .ZN(n784) );
  XNOR2_X1 U875 ( .A(n784), .B(KEYINPUT88), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G140), .A2(n867), .ZN(n785) );
  NAND2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(n787), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n872), .A2(G116), .ZN(n788) );
  XOR2_X1 U880 ( .A(KEYINPUT89), .B(n788), .Z(n790) );
  NAND2_X1 U881 ( .A1(n871), .A2(G128), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U883 ( .A(n791), .B(KEYINPUT35), .Z(n792) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U885 ( .A(KEYINPUT36), .B(n794), .Z(n795) );
  XOR2_X1 U886 ( .A(KEYINPUT90), .B(n795), .Z(n883) );
  XOR2_X1 U887 ( .A(G2067), .B(KEYINPUT37), .Z(n796) );
  XNOR2_X1 U888 ( .A(KEYINPUT87), .B(n796), .ZN(n827) );
  NOR2_X1 U889 ( .A1(n883), .A2(n827), .ZN(n981) );
  NAND2_X1 U890 ( .A1(n829), .A2(n981), .ZN(n825) );
  NAND2_X1 U891 ( .A1(n871), .A2(G129), .ZN(n798) );
  NAND2_X1 U892 ( .A1(G141), .A2(n867), .ZN(n797) );
  NAND2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n866), .A2(G105), .ZN(n799) );
  XOR2_X1 U895 ( .A(KEYINPUT38), .B(n799), .Z(n800) );
  NOR2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n872), .A2(G117), .ZN(n802) );
  NAND2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n862) );
  AND2_X1 U899 ( .A1(n862), .A2(G1996), .ZN(n970) );
  NAND2_X1 U900 ( .A1(n871), .A2(G119), .ZN(n806) );
  NAND2_X1 U901 ( .A1(G95), .A2(n866), .ZN(n804) );
  XOR2_X1 U902 ( .A(KEYINPUT91), .B(n804), .Z(n805) );
  NAND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n872), .A2(G107), .ZN(n808) );
  NAND2_X1 U905 ( .A1(G131), .A2(n867), .ZN(n807) );
  NAND2_X1 U906 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n810), .A2(n809), .ZN(n878) );
  INV_X1 U908 ( .A(G1991), .ZN(n818) );
  NOR2_X1 U909 ( .A1(n878), .A2(n818), .ZN(n968) );
  OR2_X1 U910 ( .A1(n970), .A2(n968), .ZN(n811) );
  NAND2_X1 U911 ( .A1(n811), .A2(n829), .ZN(n817) );
  XNOR2_X1 U912 ( .A(G1986), .B(G290), .ZN(n993) );
  NAND2_X1 U913 ( .A1(n829), .A2(n993), .ZN(n812) );
  NAND2_X1 U914 ( .A1(n814), .A2(n813), .ZN(n816) );
  XNOR2_X1 U915 ( .A(n816), .B(n815), .ZN(n832) );
  NOR2_X1 U916 ( .A1(G1996), .A2(n862), .ZN(n974) );
  INV_X1 U917 ( .A(n817), .ZN(n822) );
  AND2_X1 U918 ( .A1(n818), .A2(n878), .ZN(n967) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n819) );
  XNOR2_X1 U920 ( .A(KEYINPUT104), .B(n819), .ZN(n820) );
  NOR2_X1 U921 ( .A1(n967), .A2(n820), .ZN(n821) );
  NOR2_X1 U922 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U923 ( .A1(n974), .A2(n823), .ZN(n824) );
  XNOR2_X1 U924 ( .A(KEYINPUT39), .B(n824), .ZN(n826) );
  NAND2_X1 U925 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n883), .A2(n827), .ZN(n985) );
  NAND2_X1 U927 ( .A1(n828), .A2(n985), .ZN(n830) );
  NAND2_X1 U928 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n834), .ZN(G217) );
  NAND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n836) );
  INV_X1 U933 ( .A(G661), .ZN(n835) );
  NOR2_X1 U934 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n837), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U937 ( .A1(n839), .A2(n838), .ZN(G188) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G69), .ZN(G235) );
  NOR2_X1 U942 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n842), .B(KEYINPUT110), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  NAND2_X1 U945 ( .A1(G124), .A2(n871), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n843), .B(KEYINPUT44), .ZN(n845) );
  NAND2_X1 U947 ( .A1(n866), .A2(G100), .ZN(n844) );
  NAND2_X1 U948 ( .A1(n845), .A2(n844), .ZN(n849) );
  NAND2_X1 U949 ( .A1(n872), .A2(G112), .ZN(n847) );
  NAND2_X1 U950 ( .A1(G136), .A2(n867), .ZN(n846) );
  NAND2_X1 U951 ( .A1(n847), .A2(n846), .ZN(n848) );
  NOR2_X1 U952 ( .A1(n849), .A2(n848), .ZN(G162) );
  NAND2_X1 U953 ( .A1(n866), .A2(G106), .ZN(n851) );
  NAND2_X1 U954 ( .A1(G142), .A2(n867), .ZN(n850) );
  NAND2_X1 U955 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n852), .B(KEYINPUT45), .ZN(n854) );
  NAND2_X1 U957 ( .A1(G118), .A2(n872), .ZN(n853) );
  NAND2_X1 U958 ( .A1(n854), .A2(n853), .ZN(n857) );
  NAND2_X1 U959 ( .A1(G130), .A2(n871), .ZN(n855) );
  XNOR2_X1 U960 ( .A(KEYINPUT113), .B(n855), .ZN(n856) );
  NOR2_X1 U961 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U962 ( .A(G164), .B(n858), .ZN(n882) );
  XOR2_X1 U963 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n860) );
  XNOR2_X1 U964 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n859) );
  XNOR2_X1 U965 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U966 ( .A(n971), .B(n861), .ZN(n864) );
  XOR2_X1 U967 ( .A(G160), .B(n862), .Z(n863) );
  XNOR2_X1 U968 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U969 ( .A(n865), .B(G162), .Z(n880) );
  NAND2_X1 U970 ( .A1(n866), .A2(G103), .ZN(n869) );
  NAND2_X1 U971 ( .A1(G139), .A2(n867), .ZN(n868) );
  NAND2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U973 ( .A(KEYINPUT114), .B(n870), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G127), .A2(n871), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G115), .A2(n872), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n963) );
  XNOR2_X1 U979 ( .A(n878), .B(n963), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n885) );
  NOR2_X1 U983 ( .A1(G37), .A2(n885), .ZN(G395) );
  XNOR2_X1 U984 ( .A(n1001), .B(G286), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n888), .B(G171), .ZN(n889) );
  NOR2_X1 U987 ( .A1(G37), .A2(n889), .ZN(G397) );
  XNOR2_X1 U988 ( .A(KEYINPUT111), .B(n890), .ZN(G319) );
  XOR2_X1 U989 ( .A(G2100), .B(G2096), .Z(n892) );
  XNOR2_X1 U990 ( .A(KEYINPUT42), .B(G2678), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U992 ( .A(KEYINPUT43), .B(G2090), .Z(n894) );
  XNOR2_X1 U993 ( .A(G2067), .B(G2072), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U995 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U996 ( .A(G2078), .B(G2084), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(G227) );
  XNOR2_X1 U998 ( .A(G1986), .B(KEYINPUT112), .ZN(n908) );
  XOR2_X1 U999 ( .A(G1981), .B(G1971), .Z(n900) );
  XNOR2_X1 U1000 ( .A(G1966), .B(G1961), .ZN(n899) );
  XNOR2_X1 U1001 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U1002 ( .A(G1976), .B(G1956), .Z(n902) );
  XNOR2_X1 U1003 ( .A(G1996), .B(G1991), .ZN(n901) );
  XNOR2_X1 U1004 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1005 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1006 ( .A(G2474), .B(KEYINPUT41), .ZN(n905) );
  XNOR2_X1 U1007 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(n908), .B(n907), .ZN(G229) );
  OR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n909) );
  XOR2_X1 U1011 ( .A(KEYINPUT117), .B(n909), .Z(n910) );
  XNOR2_X1 U1012 ( .A(n910), .B(KEYINPUT49), .ZN(n911) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n911), .ZN(n912) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n912), .ZN(n913) );
  NOR2_X1 U1015 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n915), .B(KEYINPUT118), .ZN(G308) );
  INV_X1 U1017 ( .A(G308), .ZN(G225) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1019 ( .A(G1991), .B(G25), .ZN(n917) );
  XNOR2_X1 U1020 ( .A(G33), .B(G2072), .ZN(n916) );
  NOR2_X1 U1021 ( .A1(n917), .A2(n916), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(G32), .B(n918), .ZN(n919) );
  NAND2_X1 U1023 ( .A1(n919), .A2(G28), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(KEYINPUT120), .B(G2067), .ZN(n920) );
  XNOR2_X1 U1025 ( .A(G26), .B(n920), .ZN(n921) );
  NOR2_X1 U1026 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(G27), .B(n925), .ZN(n926) );
  NOR2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1030 ( .A(KEYINPUT53), .B(n928), .Z(n931) );
  XOR2_X1 U1031 ( .A(KEYINPUT54), .B(G34), .Z(n929) );
  XNOR2_X1 U1032 ( .A(G2084), .B(n929), .ZN(n930) );
  NAND2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(G35), .B(G2090), .ZN(n932) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1036 ( .A(KEYINPUT121), .B(n934), .Z(n935) );
  NOR2_X1 U1037 ( .A1(G29), .A2(n935), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(KEYINPUT55), .B(n936), .ZN(n1023) );
  XNOR2_X1 U1039 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n937) );
  XNOR2_X1 U1040 ( .A(n937), .B(KEYINPUT61), .ZN(n959) );
  XNOR2_X1 U1041 ( .A(G20), .B(n938), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(G1341), .B(G19), .ZN(n940) );
  XNOR2_X1 U1043 ( .A(G1981), .B(G6), .ZN(n939) );
  NOR2_X1 U1044 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1045 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1046 ( .A(KEYINPUT59), .B(G1348), .Z(n943) );
  XNOR2_X1 U1047 ( .A(G4), .B(n943), .ZN(n944) );
  NOR2_X1 U1048 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1049 ( .A(KEYINPUT60), .B(n946), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G21), .ZN(n948) );
  XNOR2_X1 U1051 ( .A(G5), .B(G1961), .ZN(n947) );
  NOR2_X1 U1052 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1053 ( .A1(n950), .A2(n949), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(G1986), .B(G24), .ZN(n952) );
  XNOR2_X1 U1055 ( .A(G1971), .B(G22), .ZN(n951) );
  NOR2_X1 U1056 ( .A1(n952), .A2(n951), .ZN(n954) );
  XOR2_X1 U1057 ( .A(G1976), .B(G23), .Z(n953) );
  NAND2_X1 U1058 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1059 ( .A(KEYINPUT58), .B(n955), .ZN(n956) );
  NOR2_X1 U1060 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1061 ( .A(n959), .B(n958), .ZN(n960) );
  NOR2_X1 U1062 ( .A1(G16), .A2(n960), .ZN(n961) );
  XNOR2_X1 U1063 ( .A(KEYINPUT127), .B(n961), .ZN(n962) );
  NAND2_X1 U1064 ( .A1(n962), .A2(G11), .ZN(n1021) );
  XOR2_X1 U1065 ( .A(G2072), .B(n963), .Z(n965) );
  XOR2_X1 U1066 ( .A(G164), .B(G2078), .Z(n964) );
  NOR2_X1 U1067 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1068 ( .A(KEYINPUT50), .B(n966), .Z(n984) );
  NOR2_X1 U1069 ( .A1(n968), .A2(n967), .ZN(n979) );
  XOR2_X1 U1070 ( .A(G160), .B(G2084), .Z(n969) );
  NOR2_X1 U1071 ( .A1(n970), .A2(n969), .ZN(n972) );
  NAND2_X1 U1072 ( .A1(n972), .A2(n971), .ZN(n977) );
  XOR2_X1 U1073 ( .A(G2090), .B(G162), .Z(n973) );
  NOR2_X1 U1074 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1075 ( .A(n975), .B(KEYINPUT51), .ZN(n976) );
  NOR2_X1 U1076 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1077 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1079 ( .A(KEYINPUT119), .B(n982), .ZN(n983) );
  NOR2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(n987), .B(KEYINPUT52), .ZN(n988) );
  NAND2_X1 U1083 ( .A1(n988), .A2(G29), .ZN(n1019) );
  XNOR2_X1 U1084 ( .A(KEYINPUT56), .B(G16), .ZN(n1017) );
  XNOR2_X1 U1085 ( .A(G1341), .B(KEYINPUT124), .ZN(n990) );
  XNOR2_X1 U1086 ( .A(n990), .B(n989), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1090 ( .A(G1961), .B(G301), .Z(n997) );
  XNOR2_X1 U1091 ( .A(KEYINPUT123), .B(n997), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1015) );
  XNOR2_X1 U1093 ( .A(n1000), .B(G1956), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(n1001), .B(G1348), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(G1971), .A2(G303), .ZN(n1002) );
  NAND2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(G168), .B(G1966), .Z(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1101 ( .A(KEYINPUT57), .B(n1010), .Z(n1011) );
  XOR2_X1 U1102 ( .A(KEYINPUT122), .B(n1011), .Z(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

