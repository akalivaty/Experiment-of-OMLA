//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960;
  NAND2_X1  g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT7), .ZN(new_n203));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204));
  INV_X1    g003(.A(G85gat), .ZN(new_n205));
  INV_X1    g004(.A(G92gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(KEYINPUT8), .A2(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G99gat), .B(G106gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT15), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  OAI22_X1  g013(.A1(KEYINPUT91), .A2(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT91), .A2(KEYINPUT14), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT92), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n217), .A2(KEYINPUT92), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n214), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT94), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n212), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  INV_X1    g025(.A(G50gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(KEYINPUT94), .A3(G43gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n229), .A2(KEYINPUT95), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n217), .B1(KEYINPUT93), .B2(new_n214), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT93), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n213), .A2(new_n232), .B1(G29gat), .B2(G36gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(KEYINPUT95), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n230), .A2(new_n231), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n211), .B1(new_n223), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(G232gat), .A2(G233gat), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n237), .A2(KEYINPUT41), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT100), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT100), .B1(new_n236), .B2(new_n238), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n223), .A2(new_n235), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT17), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT17), .B1(new_n223), .B2(new_n235), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(new_n210), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n241), .A2(new_n242), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G190gat), .B(G218gat), .Z(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n245), .A2(new_n247), .ZN(new_n251));
  INV_X1    g050(.A(new_n242), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n236), .A2(KEYINPUT100), .A3(new_n238), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n249), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT101), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n254), .B2(new_n255), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n237), .A2(KEYINPUT41), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(G134gat), .ZN(new_n261));
  INV_X1    g060(.A(G162gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n259), .A2(KEYINPUT102), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT102), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT101), .B1(new_n248), .B2(new_n249), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n267), .B2(new_n263), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n257), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT102), .B1(new_n259), .B2(new_n264), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n266), .A3(new_n263), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n270), .A2(new_n256), .A3(new_n271), .A4(new_n250), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G57gat), .B(G64gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT97), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G71gat), .A2(G78gat), .ZN(new_n278));
  OR2_X1    g077(.A1(G71gat), .A2(G78gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT9), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n278), .B(new_n279), .C1(new_n275), .C2(new_n280), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT98), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT98), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n282), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT21), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G127gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G231gat), .ZN(new_n293));
  INV_X1    g092(.A(G233gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n290), .B(G127gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(G231gat), .A3(G233gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G15gat), .B(G22gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT16), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(G1gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(G1gat), .B2(new_n299), .ZN(new_n302));
  INV_X1    g101(.A(G8gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(new_n288), .B2(new_n289), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT99), .B(G155gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n298), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n298), .A2(new_n307), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n311));
  XNOR2_X1  g110(.A(G183gat), .B(G211gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n308), .A2(new_n313), .A3(new_n309), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n274), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G113gat), .B(G141gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(G197gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT11), .ZN(new_n321));
  INV_X1    g120(.A(G169gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT12), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n304), .B1(new_n246), .B2(KEYINPUT96), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n304), .A2(KEYINPUT96), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n223), .B(new_n235), .C1(new_n326), .C2(KEYINPUT17), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G229gat), .A2(G233gat), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT18), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT18), .ZN(new_n331));
  INV_X1    g130(.A(new_n329), .ZN(new_n332));
  AOI211_X1 g131(.A(new_n331), .B(new_n332), .C1(new_n325), .C2(new_n327), .ZN(new_n333));
  INV_X1    g132(.A(new_n304), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n243), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n329), .B(KEYINPUT13), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n330), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT90), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n324), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n324), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n328), .A2(new_n329), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n331), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n328), .A2(KEYINPUT18), .A3(new_n329), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g145(.A(KEYINPUT90), .B(new_n342), .C1(new_n346), .C2(new_n338), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G230gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(new_n294), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n210), .B1(new_n285), .B2(new_n287), .ZN(new_n353));
  XOR2_X1   g152(.A(KEYINPUT103), .B(KEYINPUT10), .Z(new_n354));
  NOR2_X1   g153(.A1(new_n211), .A2(new_n284), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n210), .A2(KEYINPUT10), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n288), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n352), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n288), .A2(new_n211), .ZN(new_n361));
  INV_X1    g160(.A(new_n355), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n352), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G120gat), .B(G148gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(G176gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(G204gat), .ZN(new_n366));
  OR3_X1    g165(.A1(new_n360), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(new_n360), .B2(new_n363), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n349), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT34), .ZN(new_n372));
  NAND2_X1  g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT23), .ZN(new_n375));
  NOR3_X1   g174(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT66), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT25), .B1(new_n380), .B2(KEYINPUT23), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT67), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT67), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(KEYINPUT66), .B(new_n373), .C1(new_n375), .C2(new_n376), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n379), .A2(new_n382), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT68), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT23), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n380), .B(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n386), .B(KEYINPUT64), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n388), .B1(G183gat), .B2(G190gat), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n373), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n386), .B1(new_n399), .B2(KEYINPUT67), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n381), .B1(new_n403), .B2(new_n390), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n404), .A2(KEYINPUT68), .A3(new_n379), .A4(new_n392), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n395), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT27), .B(G183gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(G190gat), .ZN(new_n409));
  OR2_X1    g208(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n380), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT70), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT26), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(KEYINPUT65), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT26), .B1(new_n374), .B2(new_n413), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n373), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G183gat), .A2(G190gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n411), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n406), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G134gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(G127gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT71), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT71), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(new_n421), .A3(G127gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT72), .B(G127gat), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n423), .B(new_n425), .C1(new_n426), .C2(new_n421), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT73), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(G113gat), .B(G120gat), .Z(new_n430));
  INV_X1    g229(.A(KEYINPUT1), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n291), .A2(KEYINPUT72), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n291), .A2(KEYINPUT72), .ZN(new_n434));
  OAI21_X1  g233(.A(G134gat), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n435), .A2(KEYINPUT73), .A3(new_n423), .A4(new_n425), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n291), .A2(G134gat), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n430), .A2(new_n431), .A3(new_n438), .A4(new_n422), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT74), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n439), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT74), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n420), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n406), .A2(new_n443), .A3(new_n419), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n372), .B1(new_n449), .B2(KEYINPUT77), .ZN(new_n450));
  INV_X1    g249(.A(new_n448), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n445), .B2(new_n446), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT77), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT34), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n445), .A2(new_n451), .A3(new_n446), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n456), .B1(KEYINPUT32), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G15gat), .B(G43gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT75), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(G71gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(G99gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(KEYINPUT33), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n456), .A2(KEYINPUT32), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT76), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT76), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n456), .A2(new_n467), .A3(KEYINPUT32), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n455), .A2(new_n463), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT34), .B1(new_n452), .B2(new_n453), .ZN(new_n471));
  INV_X1    g270(.A(new_n454), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n469), .A2(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT36), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n470), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n469), .A2(new_n463), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n472), .A2(new_n471), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n455), .A2(new_n469), .A3(new_n463), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT36), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n482));
  XNOR2_X1  g281(.A(G1gat), .B(G29gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G57gat), .B(G85gat), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G225gat), .A2(G233gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G141gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(G148gat), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT81), .B(G141gat), .ZN(new_n493));
  INV_X1    g292(.A(G148gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G155gat), .A2(G162gat), .ZN(new_n496));
  INV_X1    g295(.A(G155gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n262), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n496), .B1(new_n498), .B2(KEYINPUT2), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT2), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n494), .A2(G141gat), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(new_n491), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n498), .A2(new_n496), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n495), .A2(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n437), .A2(new_n439), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n437), .B2(new_n439), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n489), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g307(.A(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT3), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT3), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n442), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT4), .ZN(new_n514));
  INV_X1    g313(.A(new_n505), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n489), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n504), .B(KEYINPUT82), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n440), .A3(KEYINPUT4), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n508), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n513), .A2(KEYINPUT4), .B1(new_n517), .B2(new_n440), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT4), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n442), .A2(new_n521), .A3(new_n509), .ZN(new_n522));
  NOR4_X1   g321(.A1(new_n520), .A2(KEYINPUT5), .A3(new_n489), .A4(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n487), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n520), .A2(new_n522), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n489), .A2(KEYINPUT5), .ZN(new_n528));
  INV_X1    g327(.A(new_n508), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n437), .A2(new_n439), .B1(new_n511), .B2(new_n504), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n521), .B1(new_n530), .B2(new_n510), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n488), .B(new_n518), .C1(new_n531), .C2(new_n505), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  AOI211_X1 g332(.A(KEYINPUT84), .B(KEYINPUT6), .C1(new_n533), .C2(new_n486), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n526), .B1(new_n534), .B2(new_n524), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT29), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n420), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G226gat), .A2(G233gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G197gat), .B(G204gat), .ZN(new_n540));
  INV_X1    g339(.A(G211gat), .ZN(new_n541));
  INV_X1    g340(.A(G218gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n540), .B1(KEYINPUT22), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G211gat), .B(G218gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n538), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT79), .B1(new_n420), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT79), .ZN(new_n549));
  AOI211_X1 g348(.A(new_n549), .B(new_n538), .C1(new_n406), .C2(new_n419), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n539), .B(new_n546), .C1(new_n548), .C2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT80), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n420), .A2(new_n547), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n549), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n420), .A2(KEYINPUT79), .A3(new_n547), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n557), .A2(KEYINPUT80), .A3(new_n546), .A4(new_n539), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n547), .B1(new_n420), .B2(new_n536), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT78), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n546), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n554), .A2(KEYINPUT78), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n561), .B(new_n562), .C1(new_n559), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n553), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G8gat), .B(G36gat), .Z(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(G64gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n206), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n568), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n553), .A2(new_n558), .A3(new_n564), .A4(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(KEYINPUT30), .A3(new_n571), .ZN(new_n572));
  OR3_X1    g371(.A1(new_n565), .A2(KEYINPUT30), .A3(new_n568), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n535), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n512), .A2(new_n536), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n562), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT3), .B1(new_n546), .B2(new_n536), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n504), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(G228gat), .A3(G233gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(G228gat), .A2(G233gat), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n576), .B(new_n580), .C1(new_n517), .C2(new_n577), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT31), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT31), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n579), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G78gat), .B(G106gat), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n583), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n583), .B2(new_n585), .ZN(new_n590));
  XNOR2_X1  g389(.A(G22gat), .B(G50gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n583), .A2(new_n585), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n586), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n591), .B1(new_n595), .B2(new_n588), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n481), .B(KEYINPUT85), .C1(new_n574), .C2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT85), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n572), .A2(new_n573), .ZN(new_n600));
  INV_X1    g399(.A(new_n535), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n474), .B1(new_n470), .B2(new_n473), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n478), .A2(KEYINPUT36), .A3(new_n479), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n599), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT40), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n608));
  INV_X1    g407(.A(new_n522), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n517), .A2(new_n440), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n611), .B2(new_n531), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT86), .B1(new_n612), .B2(new_n489), .ZN(new_n613));
  OAI211_X1 g412(.A(KEYINPUT86), .B(new_n489), .C1(new_n520), .C2(new_n522), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n608), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT86), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n527), .B2(new_n488), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n505), .A2(new_n506), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n608), .B1(new_n619), .B2(new_n488), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n616), .A2(new_n621), .A3(new_n486), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT87), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n519), .A2(new_n523), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n527), .A2(new_n528), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n529), .A2(new_n532), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT87), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n607), .A2(new_n622), .B1(new_n628), .B2(new_n487), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n622), .A2(new_n607), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n572), .A2(new_n629), .A3(new_n573), .A4(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT88), .B(KEYINPUT37), .Z(new_n633));
  NAND4_X1  g432(.A1(new_n553), .A2(new_n558), .A3(new_n564), .A4(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n634), .A2(new_n568), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n565), .A2(KEYINPUT37), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n557), .A2(new_n562), .A3(new_n539), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n561), .B(new_n546), .C1(new_n559), .C2(new_n563), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n639), .A3(KEYINPUT37), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n634), .A2(new_n632), .A3(new_n568), .A4(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n623), .B1(new_n519), .B2(new_n523), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT87), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n487), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT6), .B1(new_n533), .B2(new_n486), .ZN(new_n645));
  INV_X1    g444(.A(new_n524), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n644), .A2(new_n645), .B1(new_n646), .B2(KEYINPUT6), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n641), .A2(new_n647), .A3(new_n571), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n631), .B(new_n597), .C1(new_n637), .C2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n598), .A2(new_n606), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n593), .A2(new_n596), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n651), .B1(new_n479), .B2(new_n478), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n574), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT35), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n651), .A2(KEYINPUT35), .A3(new_n647), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n478), .A2(KEYINPUT89), .A3(new_n479), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT89), .B1(new_n478), .B2(new_n479), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n600), .B(new_n655), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  AOI211_X1 g459(.A(new_n318), .B(new_n371), .C1(new_n650), .C2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n535), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g462(.A1(new_n572), .A2(new_n573), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n300), .A2(new_n303), .ZN(new_n665));
  NAND2_X1  g464(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n666));
  AND4_X1   g465(.A1(new_n664), .A2(new_n661), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n303), .B1(new_n661), .B2(new_n664), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT42), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(KEYINPUT42), .B2(new_n667), .ZN(G1325gat));
  NOR2_X1   g469(.A1(new_n657), .A2(new_n658), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(G15gat), .B1(new_n661), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n605), .A2(G15gat), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(new_n661), .B2(new_n674), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n661), .A2(new_n651), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  AOI21_X1  g477(.A(new_n274), .B1(new_n650), .B2(new_n660), .ZN(new_n679));
  INV_X1    g478(.A(new_n317), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n679), .A2(new_n680), .A3(new_n370), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n219), .A3(new_n535), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT104), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT104), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT45), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n683), .A2(KEYINPUT45), .A3(new_n684), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n317), .B(KEYINPUT105), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n689), .A2(new_n370), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n650), .A2(new_n660), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n273), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n597), .B1(new_n637), .B2(new_n648), .ZN(new_n693));
  AND4_X1   g492(.A1(new_n573), .A2(new_n572), .A3(new_n629), .A4(new_n630), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n604), .B(new_n603), .C1(new_n574), .C2(new_n597), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT106), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n602), .A2(new_n605), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n699), .A3(new_n649), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n274), .B1(new_n701), .B2(new_n660), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n690), .B(new_n692), .C1(new_n702), .C2(KEYINPUT44), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT107), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n697), .A2(new_n700), .B1(new_n654), .B2(new_n659), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(new_n274), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n707), .A2(new_n708), .A3(new_n690), .A4(new_n692), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n601), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n687), .B(new_n688), .C1(new_n710), .C2(new_n219), .ZN(G1328gat));
  NAND3_X1  g510(.A1(new_n681), .A2(new_n220), .A3(new_n664), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(KEYINPUT46), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n713), .A2(KEYINPUT46), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n600), .B1(new_n704), .B2(new_n709), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n220), .B2(new_n717), .ZN(G1329gat));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719));
  INV_X1    g518(.A(G43gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n709), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n721), .B2(new_n605), .ZN(new_n722));
  INV_X1    g521(.A(new_n681), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n723), .A2(G43gat), .A3(new_n671), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n719), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n724), .ZN(new_n726));
  OAI21_X1  g525(.A(G43gat), .B1(new_n703), .B2(new_n481), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(KEYINPUT47), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(G1330gat));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n227), .B1(new_n721), .B2(new_n651), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n651), .B1(new_n723), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n227), .B1(new_n681), .B2(KEYINPUT109), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n730), .B1(new_n731), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G50gat), .B1(new_n703), .B2(new_n597), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n737), .B(KEYINPUT48), .C1(new_n733), .C2(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1331gat));
  NOR3_X1   g538(.A1(new_n706), .A2(new_n318), .A3(new_n348), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n369), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n535), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g543(.A1(new_n741), .A2(new_n600), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(G1333gat));
  INV_X1    g548(.A(G71gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n671), .B(KEYINPUT110), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n742), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G71gat), .B1(new_n741), .B2(new_n481), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n742), .A2(new_n651), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g557(.A1(new_n707), .A2(new_n692), .ZN(new_n759));
  INV_X1    g558(.A(new_n369), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n317), .A2(new_n760), .A3(new_n348), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(new_n535), .A3(new_n761), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n762), .A2(KEYINPUT111), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(KEYINPUT111), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(G85gat), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n317), .A2(new_n348), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n702), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n767), .A2(KEYINPUT112), .A3(KEYINPUT51), .ZN(new_n768));
  NAND2_X1  g567(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n769));
  OR2_X1    g568(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n702), .A2(new_n766), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n772), .A2(new_n205), .A3(new_n535), .A4(new_n369), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n765), .A2(new_n773), .ZN(G1336gat));
  NAND4_X1  g573(.A1(new_n707), .A2(new_n664), .A3(new_n692), .A4(new_n761), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G92gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT113), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n600), .A2(G92gat), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n768), .A2(new_n369), .A3(new_n771), .A4(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n775), .A2(new_n780), .A3(G92gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT52), .ZN(new_n783));
  XOR2_X1   g582(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n784));
  NAND3_X1  g583(.A1(new_n779), .A2(new_n776), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1337gat));
  NAND3_X1  g585(.A1(new_n772), .A2(new_n369), .A3(new_n672), .ZN(new_n787));
  INV_X1    g586(.A(G99gat), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n759), .A2(new_n761), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n481), .A2(new_n788), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n790), .ZN(G1338gat));
  NAND4_X1  g590(.A1(new_n707), .A2(new_n651), .A3(new_n692), .A4(new_n761), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G106gat), .ZN(new_n793));
  INV_X1    g592(.A(G106gat), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n768), .A2(new_n794), .A3(new_n369), .A4(new_n771), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n795), .B2(new_n597), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT53), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n798), .B(new_n793), .C1(new_n795), .C2(new_n597), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1339gat));
  NOR2_X1   g599(.A1(new_n664), .A2(new_n601), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802));
  INV_X1    g601(.A(new_n354), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n361), .A2(new_n803), .A3(new_n362), .ZN(new_n804));
  INV_X1    g603(.A(new_n358), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n351), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n359), .A2(new_n806), .A3(KEYINPUT54), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT115), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n359), .A2(new_n806), .A3(new_n809), .A4(KEYINPUT54), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g610(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n812));
  NAND2_X1  g611(.A1(new_n360), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n366), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n367), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT117), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n811), .A2(new_n366), .A3(new_n813), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n817), .A2(new_n818), .B1(new_n341), .B2(new_n347), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n814), .A2(new_n820), .A3(new_n367), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n816), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n339), .A2(new_n324), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n328), .A2(new_n329), .B1(new_n335), .B2(new_n337), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n323), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n369), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n826), .B(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n273), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n823), .A2(new_n825), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n269), .B2(new_n272), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n818), .A2(new_n817), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n816), .A4(new_n821), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n689), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n318), .A2(new_n369), .A3(new_n348), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n802), .B1(new_n838), .B2(new_n597), .ZN(new_n839));
  AOI211_X1 g638(.A(KEYINPUT119), .B(new_n651), .C1(new_n835), .C2(new_n837), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n672), .B(new_n801), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n349), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n601), .B1(new_n835), .B2(new_n837), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n652), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT120), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(KEYINPUT120), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n600), .A3(new_n846), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n349), .A2(G113gat), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n842), .B1(new_n847), .B2(new_n848), .ZN(G1340gat));
  NOR2_X1   g648(.A1(new_n760), .A2(G120gat), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n845), .A2(new_n600), .A3(new_n846), .A4(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G120gat), .B1(new_n841), .B2(new_n760), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT121), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n855), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1341gat));
  INV_X1    g656(.A(new_n426), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n847), .B2(new_n680), .ZN(new_n859));
  OR3_X1    g658(.A1(new_n841), .A2(new_n858), .A3(new_n689), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OR4_X1    g661(.A1(new_n861), .A2(new_n841), .A3(new_n858), .A4(new_n689), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n859), .A2(new_n862), .A3(new_n863), .ZN(G1342gat));
  AND3_X1   g663(.A1(new_n845), .A2(new_n600), .A3(new_n846), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT56), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n865), .A2(new_n866), .A3(new_n421), .A4(new_n273), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n841), .B2(new_n274), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n845), .A2(new_n421), .A3(new_n600), .A4(new_n846), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT56), .B1(new_n869), .B2(new_n274), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(G1343gat));
  AOI21_X1  g670(.A(new_n597), .B1(new_n835), .B2(new_n837), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n826), .ZN(new_n875));
  INV_X1    g674(.A(new_n815), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n819), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n833), .B1(new_n877), .B2(new_n273), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n836), .B1(new_n878), .B2(new_n680), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT57), .B1(new_n879), .B2(new_n597), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n605), .A2(new_n601), .A3(new_n664), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n874), .A2(new_n880), .A3(new_n348), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n493), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT123), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n651), .B1(new_n843), .B2(new_n885), .ZN(new_n886));
  AOI211_X1 g685(.A(KEYINPUT124), .B(new_n601), .C1(new_n835), .C2(new_n837), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n605), .A2(new_n664), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n888), .A2(new_n490), .A3(new_n348), .A4(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n882), .A2(new_n891), .A3(new_n493), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n884), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT58), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT58), .B1(new_n882), .B2(new_n493), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n890), .A2(KEYINPUT125), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT125), .B1(new_n890), .B2(new_n895), .ZN(new_n897));
  OAI22_X1  g696(.A1(new_n893), .A2(new_n894), .B1(new_n896), .B2(new_n897), .ZN(G1344gat));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n874), .A2(new_n880), .A3(new_n881), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n760), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n494), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n872), .A2(new_n873), .ZN(new_n903));
  OR3_X1    g702(.A1(new_n879), .A2(KEYINPUT57), .A3(new_n597), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n903), .A2(new_n369), .A3(new_n904), .A4(new_n881), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n899), .B1(new_n905), .B2(G148gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n889), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n369), .A2(new_n494), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n902), .A2(new_n906), .B1(new_n907), .B2(new_n908), .ZN(G1345gat));
  NOR3_X1   g708(.A1(new_n900), .A2(new_n497), .A3(new_n689), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n888), .A2(new_n317), .A3(new_n889), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n497), .ZN(G1346gat));
  NOR3_X1   g711(.A1(new_n900), .A2(new_n262), .A3(new_n274), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n888), .A2(new_n273), .A3(new_n889), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n262), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n600), .A2(new_n535), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n751), .B(new_n916), .C1(new_n839), .C2(new_n840), .ZN(new_n917));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n349), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n838), .A2(new_n652), .A3(new_n916), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n322), .A3(new_n348), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n918), .A2(new_n921), .ZN(G1348gat));
  INV_X1    g721(.A(G176gat), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n917), .A2(new_n923), .A3(new_n760), .ZN(new_n924));
  AOI21_X1  g723(.A(G176gat), .B1(new_n920), .B2(new_n369), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  OAI21_X1  g725(.A(G183gat), .B1(new_n917), .B2(new_n689), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n920), .A2(new_n317), .A3(new_n407), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g729(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n931));
  OAI211_X1 g730(.A(G190gat), .B(new_n931), .C1(new_n917), .C2(new_n274), .ZN(new_n932));
  NOR2_X1   g731(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR3_X1    g733(.A1(new_n919), .A2(G190gat), .A3(new_n274), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n933), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G1351gat));
  NAND2_X1  g736(.A1(new_n481), .A2(new_n916), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n903), .A2(new_n904), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n349), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n872), .A2(new_n939), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n349), .A2(G197gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G1352gat));
  NAND3_X1  g743(.A1(new_n903), .A2(new_n369), .A3(new_n904), .ZN(new_n945));
  OAI21_X1  g744(.A(G204gat), .B1(new_n945), .B2(new_n938), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n942), .A2(G204gat), .A3(new_n760), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT127), .A3(new_n947), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT127), .B1(new_n948), .B2(new_n947), .ZN(new_n950));
  OAI221_X1 g749(.A(new_n946), .B1(new_n947), .B2(new_n948), .C1(new_n949), .C2(new_n950), .ZN(G1353gat));
  OR2_X1    g750(.A1(new_n940), .A2(new_n680), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n953));
  OAI211_X1 g752(.A(KEYINPUT63), .B(G211gat), .C1(new_n940), .C2(new_n680), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n317), .A2(new_n541), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n953), .A2(new_n955), .B1(new_n942), .B2(new_n956), .ZN(G1354gat));
  OAI21_X1  g756(.A(new_n542), .B1(new_n942), .B2(new_n274), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n273), .A2(G218gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n940), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(G1355gat));
endmodule


