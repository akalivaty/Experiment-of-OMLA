//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND3_X1  g0014(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n203), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(new_n225), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n235), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G45), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(KEYINPUT66), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT66), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G1), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n258), .B1(G33), .B2(G41), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n252), .B2(new_n248), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n257), .B1(G226), .B2(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G223), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(KEYINPUT67), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT67), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G1698), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n269), .A2(new_n271), .A3(G222), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n259), .B1(G77), .B2(new_n265), .C1(new_n268), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G179), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(new_n274), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n258), .ZN(new_n279));
  XOR2_X1   g0079(.A(KEYINPUT8), .B(G58), .Z(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  INV_X1    g0081(.A(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(G20), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n209), .A2(KEYINPUT68), .A3(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n280), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G150), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT69), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n283), .A2(new_n284), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  OAI211_X1 g0090(.A(KEYINPUT69), .B(new_n287), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n279), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G50), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n278), .A2(new_n258), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(new_n298), .A3(new_n295), .ZN(new_n299));
  INV_X1    g0099(.A(new_n295), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT70), .B1(new_n300), .B2(new_n279), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n299), .A2(new_n301), .B1(new_n208), .B2(G20), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n296), .B1(new_n302), .B2(G50), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n277), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT73), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n294), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(new_n294), .B2(new_n303), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT9), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n304), .A2(KEYINPUT73), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT9), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(new_n308), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n274), .A2(G200), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n274), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n306), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  AOI211_X1 g0120(.A(KEYINPUT10), .B(new_n318), .C1(new_n311), .C2(new_n314), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n305), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n257), .B1(G244), .B2(new_n261), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n267), .B1(new_n263), .B2(new_n264), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G238), .ZN(new_n325));
  AND2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G107), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n269), .B(new_n271), .C1(new_n326), .C2(new_n327), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n325), .B(new_n329), .C1(new_n225), .C2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(G1), .B(G13), .C1(new_n282), .C2(new_n252), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n334), .A2(G179), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n280), .A2(new_n286), .B1(G20), .B2(G77), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT15), .B(G87), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT71), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n336), .B1(new_n338), .B2(new_n289), .ZN(new_n339));
  INV_X1    g0139(.A(G77), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n339), .A2(new_n279), .B1(new_n340), .B2(new_n300), .ZN(new_n341));
  OR3_X1    g0141(.A1(new_n300), .A2(new_n279), .A3(KEYINPUT72), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n208), .A2(G20), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT72), .B1(new_n300), .B2(new_n279), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n342), .A2(G77), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n334), .A2(new_n276), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n335), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n334), .A2(G200), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n334), .A2(new_n317), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n346), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n349), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n302), .A2(new_n280), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n280), .A2(new_n295), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT7), .B1(new_n328), .B2(new_n209), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT7), .ZN(new_n359));
  NOR4_X1   g0159(.A1(new_n326), .A2(new_n327), .A3(new_n359), .A4(G20), .ZN(new_n360));
  OAI21_X1  g0160(.A(G68), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n224), .A2(new_n218), .ZN(new_n362));
  OAI21_X1  g0162(.A(G20), .B1(new_n362), .B2(new_n202), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n286), .A2(G159), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n297), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n361), .A2(KEYINPUT16), .A3(new_n366), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n357), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(G226), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n372), .B(new_n373), .C1(new_n330), .C2(new_n266), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n259), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n261), .A2(G232), .B1(new_n253), .B2(new_n255), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n375), .A2(G190), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n375), .B2(new_n376), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT79), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n375), .A2(new_n376), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G200), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n375), .A2(G190), .A3(new_n376), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT79), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n371), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n380), .B1(new_n377), .B2(new_n379), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n383), .A2(KEYINPUT79), .A3(new_n384), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(KEYINPUT17), .A3(new_n371), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n382), .A2(new_n276), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(G179), .B2(new_n382), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n393), .B1(new_n371), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n263), .A2(new_n209), .A3(new_n264), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n359), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n264), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n218), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n368), .B1(new_n400), .B2(new_n365), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(new_n370), .A3(new_n279), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n355), .B1(new_n302), .B2(new_n280), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G179), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n375), .A2(new_n405), .A3(new_n376), .ZN(new_n406));
  AOI21_X1  g0206(.A(G169), .B1(new_n375), .B2(new_n376), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(KEYINPUT18), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n396), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n353), .A2(new_n388), .A3(new_n392), .A4(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n269), .A2(new_n271), .A3(G226), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G232), .A2(G1698), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n328), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G97), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n259), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n261), .A2(G238), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT74), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n253), .A2(new_n420), .A3(new_n255), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n420), .B1(new_n253), .B2(new_n255), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n419), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT13), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT75), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n256), .A2(KEYINPUT74), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n421), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n417), .A3(new_n429), .A4(new_n419), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n430), .A2(G190), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n427), .A2(new_n421), .B1(G238), .B2(new_n261), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n429), .B1(new_n432), .B2(new_n417), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT75), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n426), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT76), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n426), .A2(new_n431), .A3(new_n435), .A4(KEYINPUT76), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT77), .B1(new_n209), .B2(G68), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n209), .A2(new_n282), .ZN(new_n442));
  INV_X1    g0242(.A(G50), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n286), .A2(KEYINPUT77), .A3(G50), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n444), .B(new_n445), .C1(new_n340), .C2(new_n289), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n446), .A2(KEYINPUT78), .A3(new_n279), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT78), .B1(new_n446), .B2(new_n279), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT11), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n279), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT78), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT11), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n446), .A2(KEYINPUT78), .A3(new_n279), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n342), .A2(G68), .A3(new_n343), .A4(new_n344), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n300), .A2(new_n218), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n457), .B(KEYINPUT12), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n449), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n378), .B1(new_n425), .B2(new_n430), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n440), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n430), .ZN(new_n465));
  OAI21_X1  g0265(.A(G169), .B1(new_n465), .B2(new_n433), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT14), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n426), .A2(new_n435), .A3(G179), .A4(new_n430), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT14), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n469), .B(G169), .C1(new_n465), .C2(new_n433), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n460), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n464), .A2(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n322), .A2(new_n411), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(G20), .B1(G33), .B2(G283), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(G33), .B2(new_n226), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n476), .B(new_n279), .C1(new_n209), .C2(G116), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT20), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G116), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n208), .B2(G33), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n342), .A2(new_n344), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT87), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT87), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n342), .A2(new_n484), .A3(new_n344), .A4(new_n481), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n300), .A2(new_n480), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n479), .A2(new_n483), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n227), .B1(new_n263), .B2(new_n264), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n269), .A2(new_n271), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n489), .A2(new_n490), .B1(new_n328), .B2(G303), .ZN(new_n491));
  OAI211_X1 g0291(.A(G264), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n333), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT81), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT5), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(G41), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n252), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n248), .A2(G1), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(G41), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(G270), .A3(new_n333), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n208), .A2(G45), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n502), .B1(new_n495), .B2(G41), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n503), .A2(G274), .A3(new_n497), .A4(new_n496), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n493), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G190), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n488), .B(new_n507), .C1(new_n378), .C2(new_n506), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT21), .ZN(new_n509));
  OAI21_X1  g0309(.A(G257), .B1(new_n326), .B2(new_n327), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n269), .A2(new_n271), .ZN(new_n511));
  INV_X1    g0311(.A(G303), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n510), .A2(new_n511), .B1(new_n265), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n492), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n259), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n504), .A3(new_n501), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G169), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n509), .B1(new_n488), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(KEYINPUT21), .B(G169), .C1(new_n493), .C2(new_n505), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n515), .A2(G179), .A3(new_n504), .A4(new_n501), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n521), .A2(KEYINPUT88), .A3(new_n487), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT88), .B1(new_n521), .B2(new_n487), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n508), .B(new_n518), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n500), .A2(G257), .A3(new_n333), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n504), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n324), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  INV_X1    g0329(.A(G244), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n330), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n490), .A2(new_n265), .A3(KEYINPUT4), .A4(G244), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n527), .B1(new_n533), .B2(new_n259), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT6), .ZN(new_n535));
  INV_X1    g0335(.A(G107), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n226), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n535), .B1(new_n537), .B2(new_n205), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(KEYINPUT6), .A3(G97), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(G20), .B1(G77), .B2(new_n286), .ZN(new_n541));
  OAI21_X1  g0341(.A(G107), .B1(new_n358), .B2(new_n360), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n297), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n300), .A2(new_n226), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n297), .B(new_n295), .C1(G1), .C2(new_n282), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(new_n226), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n534), .A2(G169), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n533), .A2(new_n259), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT80), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n533), .A2(KEYINPUT80), .A3(new_n259), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n527), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n547), .B1(new_n552), .B2(new_n405), .ZN(new_n553));
  INV_X1    g0353(.A(new_n527), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n533), .A2(KEYINPUT80), .A3(new_n259), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT80), .B1(new_n533), .B2(new_n259), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT82), .B1(new_n557), .B2(G200), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n543), .A2(new_n546), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT83), .ZN(new_n560));
  AND4_X1   g0360(.A1(new_n560), .A2(new_n548), .A3(G190), .A4(new_n554), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n534), .B2(G190), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n557), .A2(KEYINPUT82), .A3(G200), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n553), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n545), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G87), .ZN(new_n568));
  OAI211_X1 g0368(.A(G244), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G116), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n569), .B(new_n570), .C1(new_n330), .C2(new_n219), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n259), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n502), .A2(KEYINPUT84), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT84), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(new_n208), .A3(G45), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n259), .A2(new_n221), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n576), .A2(new_n577), .B1(G274), .B2(new_n498), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n378), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G190), .B2(new_n579), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n283), .A2(G97), .A3(new_n284), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n265), .A2(new_n209), .A3(G68), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n209), .B1(new_n415), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(G87), .B2(new_n206), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT85), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n584), .A2(KEYINPUT85), .A3(new_n585), .A4(new_n587), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n279), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT86), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n338), .A2(new_n300), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n593), .B1(new_n592), .B2(new_n594), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n568), .B(new_n581), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n338), .A2(new_n545), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n592), .A2(new_n594), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT86), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n572), .A2(G179), .A3(new_n578), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n333), .A2(G250), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n573), .A2(new_n575), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n604), .A2(new_n605), .B1(new_n254), .B2(new_n502), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n259), .B2(new_n571), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n603), .B1(new_n607), .B2(new_n276), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n597), .B1(new_n602), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n500), .A2(G264), .A3(new_n333), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT92), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT92), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n500), .A2(new_n613), .A3(G264), .A4(new_n333), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(G257), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n616));
  NAND2_X1  g0416(.A1(G33), .A2(G294), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n616), .B(new_n617), .C1(new_n330), .C2(new_n221), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n259), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n615), .A2(new_n504), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n504), .A3(new_n611), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n620), .A2(G200), .B1(G190), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n265), .A2(new_n209), .A3(G87), .ZN(new_n623));
  XOR2_X1   g0423(.A(KEYINPUT89), .B(KEYINPUT22), .Z(new_n624));
  XNOR2_X1  g0424(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT24), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT23), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(new_n536), .A3(G20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT90), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n627), .B2(new_n536), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n628), .A2(KEYINPUT90), .B1(new_n631), .B2(G20), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n625), .A2(new_n626), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n626), .B1(new_n625), .B2(new_n633), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n279), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n300), .A2(new_n536), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT91), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n639), .A3(KEYINPUT25), .ZN(new_n640));
  XOR2_X1   g0440(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n641));
  OAI221_X1 g0441(.A(new_n640), .B1(new_n638), .B2(new_n641), .C1(new_n545), .C2(new_n536), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n622), .A2(new_n637), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n621), .A2(G169), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n612), .A2(new_n614), .B1(new_n259), .B2(new_n618), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n504), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n645), .B1(new_n647), .B2(new_n405), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n623), .A2(new_n624), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n623), .A2(new_n624), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n633), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT24), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n297), .B1(new_n653), .B2(new_n634), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n648), .B1(new_n654), .B2(new_n642), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n644), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n610), .A2(new_n656), .ZN(new_n657));
  AND4_X1   g0457(.A1(new_n474), .A2(new_n525), .A3(new_n566), .A4(new_n657), .ZN(G372));
  NAND2_X1  g0458(.A1(new_n388), .A2(new_n392), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n464), .A2(new_n349), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n472), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT95), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n404), .A2(new_n662), .A3(new_n408), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n404), .B2(new_n408), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n663), .A2(new_n664), .A3(new_n393), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT95), .B1(new_n371), .B2(new_n395), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n404), .A2(new_n662), .A3(new_n408), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT18), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n320), .A2(new_n321), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n670), .A2(new_n671), .B1(new_n304), .B2(new_n277), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n521), .A2(new_n487), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n655), .A2(new_n518), .A3(new_n673), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n600), .A2(new_n601), .B1(G87), .B2(new_n567), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n595), .A2(new_n596), .B1(new_n338), .B2(new_n545), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT93), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n608), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n603), .B(KEYINPUT93), .C1(new_n607), .C2(new_n276), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n675), .A2(new_n581), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n566), .A2(new_n674), .A3(new_n644), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n680), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n597), .B(new_n553), .C1(new_n602), .C2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n676), .A2(new_n608), .ZN(new_n688));
  XOR2_X1   g0488(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n688), .A2(new_n553), .A3(new_n597), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n682), .A2(new_n683), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n474), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n672), .A2(new_n694), .ZN(G369));
  NAND2_X1  g0495(.A1(new_n518), .A2(new_n673), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT96), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G213), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n698), .A2(new_n699), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  XOR2_X1   g0504(.A(KEYINPUT97), .B(G343), .Z(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n488), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n696), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n524), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n707), .B1(new_n637), .B2(new_n643), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n656), .A2(new_n713), .B1(new_n655), .B2(new_n707), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n717), .A2(new_n707), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(new_n655), .A3(new_n644), .ZN(new_n719));
  INV_X1    g0519(.A(new_n707), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n655), .B2(new_n720), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n716), .A2(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n212), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n216), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n693), .A2(new_n707), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n597), .B(new_n553), .C1(new_n602), .C2(new_n609), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(KEYINPUT100), .A3(new_n689), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n683), .A2(KEYINPUT26), .A3(new_n553), .A4(new_n597), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT100), .B1(new_n733), .B2(new_n689), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n553), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT82), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n552), .B2(new_n378), .ZN(new_n741));
  INV_X1    g0541(.A(new_n562), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n534), .A2(new_n560), .A3(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n741), .A2(new_n744), .A3(new_n559), .A4(new_n565), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n681), .A2(new_n739), .A3(new_n745), .A4(new_n644), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n655), .B(new_n518), .C1(new_n522), .C2(new_n523), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n683), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(KEYINPUT29), .B(new_n707), .C1(new_n738), .C2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n657), .A2(new_n566), .A3(new_n525), .A4(new_n707), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n516), .A2(new_n405), .A3(new_n579), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n620), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n557), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT30), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n548), .A2(new_n607), .A3(new_n554), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n615), .A2(new_n619), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n520), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n755), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n506), .A2(new_n646), .A3(G179), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n761), .A2(new_n756), .A3(KEYINPUT30), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n754), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT98), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT31), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n707), .A2(new_n765), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n764), .B1(new_n763), .B2(new_n766), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n757), .A2(new_n759), .A3(new_n755), .ZN(new_n770));
  OAI21_X1  g0570(.A(KEYINPUT30), .B1(new_n761), .B2(new_n756), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n770), .A2(new_n771), .B1(new_n753), .B2(new_n557), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT99), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n720), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n754), .B(new_n773), .C1(new_n760), .C2(new_n762), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n765), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n751), .A2(new_n769), .A3(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n732), .A2(new_n750), .B1(G330), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n729), .B1(new_n779), .B2(G1), .ZN(G364));
  XOR2_X1   g0580(.A(new_n711), .B(KEYINPUT101), .Z(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G13), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n208), .B1(new_n784), .B2(G45), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n724), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n782), .B(new_n788), .C1(G330), .C2(new_n710), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT102), .Z(new_n790));
  NAND2_X1  g0590(.A1(new_n212), .A2(new_n265), .ZN(new_n791));
  INV_X1    g0591(.A(G355), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n792), .B1(G116), .B2(new_n212), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n243), .A2(G45), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n212), .A2(new_n328), .ZN(new_n795));
  INV_X1    g0595(.A(new_n216), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n249), .A2(new_n251), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n793), .B1(new_n794), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n258), .B1(G20), .B2(new_n276), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n787), .B1(new_n799), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n317), .A2(new_n378), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n209), .A2(G179), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n209), .A2(new_n405), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G190), .A2(G200), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n512), .A2(new_n809), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(KEYINPUT33), .B(G317), .Z(new_n815));
  NOR2_X1   g0615(.A1(new_n378), .A2(G190), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n808), .A2(new_n816), .ZN(new_n818));
  INV_X1    g0618(.A(G283), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n815), .A2(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n317), .A2(G179), .A3(G200), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n209), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G294), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n810), .A2(new_n807), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n265), .B1(new_n827), .B2(G326), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n810), .A2(G190), .A3(new_n378), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n808), .A2(new_n811), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n830), .A2(G322), .B1(new_n832), .B2(G329), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n821), .A2(new_n825), .A3(new_n828), .A4(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n826), .A2(new_n443), .B1(new_n812), .B2(new_n340), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n829), .A2(new_n224), .B1(new_n809), .B2(new_n220), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G159), .ZN(new_n838));
  OR3_X1    g0638(.A1(new_n831), .A2(KEYINPUT32), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT32), .B1(new_n831), .B2(new_n838), .ZN(new_n840));
  INV_X1    g0640(.A(new_n818), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n328), .B1(new_n841), .B2(G107), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n837), .A2(new_n839), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n823), .A2(new_n226), .B1(new_n817), .B2(new_n218), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT103), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n834), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n806), .B1(new_n846), .B2(new_n803), .ZN(new_n847));
  INV_X1    g0647(.A(new_n802), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n710), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n790), .A2(new_n849), .ZN(G396));
  NOR2_X1   g0650(.A1(new_n348), .A2(new_n720), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n346), .A2(new_n720), .B1(new_n352), .B2(new_n350), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n853), .B2(new_n349), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n730), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n854), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n693), .A2(new_n707), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n778), .A2(G330), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n787), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n265), .B1(new_n809), .B2(new_n443), .ZN(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n818), .A2(new_n218), .B1(new_n831), .B2(new_n863), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n862), .B(new_n864), .C1(G58), .C2(new_n824), .ZN(new_n865));
  INV_X1    g0665(.A(G137), .ZN(new_n866));
  INV_X1    g0666(.A(G150), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n826), .A2(new_n866), .B1(new_n817), .B2(new_n867), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT105), .Z(new_n869));
  INV_X1    g0669(.A(G143), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n869), .B1(new_n870), .B2(new_n829), .C1(new_n838), .C2(new_n812), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT34), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n865), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n872), .B2(new_n871), .ZN(new_n874));
  INV_X1    g0674(.A(new_n817), .ZN(new_n875));
  AOI22_X1  g0675(.A1(G283), .A2(new_n875), .B1(new_n841), .B2(G87), .ZN(new_n876));
  INV_X1    g0676(.A(new_n812), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n265), .B1(new_n877), .B2(G116), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n876), .B(new_n878), .C1(new_n226), .C2(new_n823), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n809), .A2(new_n536), .B1(new_n831), .B2(new_n813), .ZN(new_n880));
  INV_X1    g0680(.A(G294), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n829), .A2(new_n881), .B1(new_n826), .B2(new_n512), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT104), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n803), .B1(new_n874), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n803), .A2(new_n800), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n788), .B1(new_n340), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n885), .B(new_n887), .C1(new_n856), .C2(new_n801), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n861), .A2(new_n888), .ZN(G384));
  NOR3_X1   g0689(.A1(new_n216), .A2(new_n340), .A3(new_n362), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n201), .A2(new_n218), .ZN(new_n891));
  OAI211_X1 g0691(.A(G1), .B(new_n783), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT106), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT36), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n480), .B(new_n215), .C1(new_n540), .C2(KEYINPUT35), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(KEYINPUT35), .B2(new_n540), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n893), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n894), .B2(new_n896), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n388), .A2(new_n410), .A3(new_n392), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n703), .B1(new_n402), .B2(new_n403), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n404), .A2(new_n408), .ZN(new_n903));
  INV_X1    g0703(.A(new_n901), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n386), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n901), .B1(new_n391), .B2(new_n371), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n908), .A3(new_n903), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n902), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n902), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n899), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n707), .B1(new_n763), .B2(KEYINPUT99), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(KEYINPUT31), .A3(new_n775), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n751), .A2(new_n777), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n462), .B1(new_n438), .B2(new_n439), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n460), .B(new_n720), .C1(new_n917), .C2(new_n471), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n720), .A2(new_n460), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n464), .A2(new_n472), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n854), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n913), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n666), .A2(new_n667), .ZN(new_n924));
  AOI211_X1 g0724(.A(KEYINPUT108), .B(new_n908), .C1(new_n924), .C2(new_n907), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n388), .B(new_n392), .C1(new_n665), .C2(new_n668), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n925), .B1(new_n926), .B2(new_n901), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n386), .B(new_n904), .C1(new_n663), .C2(new_n664), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT37), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(KEYINPUT108), .A3(new_n909), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n916), .B(new_n921), .C1(new_n931), .C2(new_n911), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n923), .B1(new_n932), .B2(KEYINPUT40), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT109), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n474), .A2(new_n916), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(G330), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n918), .A2(new_n920), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n851), .B(KEYINPUT107), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n940), .B1(new_n857), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n912), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n902), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n944), .A2(KEYINPUT39), .A3(new_n945), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n472), .A2(new_n720), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT108), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n928), .A2(new_n950), .A3(KEYINPUT37), .ZN(new_n951));
  INV_X1    g0751(.A(new_n668), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n666), .A2(KEYINPUT18), .A3(new_n667), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n659), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n930), .B(new_n951), .C1(new_n954), .C2(new_n904), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT38), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n911), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n948), .B(new_n949), .C1(new_n957), .C2(KEYINPUT39), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n669), .A2(new_n703), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n947), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n732), .A2(new_n750), .A3(new_n474), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n672), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n960), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n938), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(KEYINPUT110), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n965), .B1(new_n208), .B2(new_n784), .C1(new_n963), .C2(new_n938), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n964), .A2(KEYINPUT110), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n898), .B1(new_n966), .B2(new_n967), .ZN(G367));
  NAND2_X1  g0768(.A1(new_n745), .A2(new_n739), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n707), .A2(new_n559), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n969), .A2(new_n970), .B1(new_n739), .B2(new_n707), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n971), .A2(KEYINPUT111), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(KEYINPUT111), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n719), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT42), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n739), .B1(new_n974), .B2(new_n655), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n707), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n683), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n675), .A2(new_n707), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n681), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n983), .B2(new_n981), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT43), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n979), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n976), .A2(new_n986), .A3(new_n985), .A4(new_n978), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OR3_X1    g0791(.A1(new_n991), .A2(new_n715), .A3(new_n974), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n991), .B1(new_n715), .B2(new_n974), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n724), .B(KEYINPUT41), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n974), .A2(new_n721), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT44), .Z(new_n996));
  NOR2_X1   g0796(.A1(new_n974), .A2(new_n721), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n716), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n719), .B1(new_n714), .B2(new_n718), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1001), .A2(new_n711), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n782), .B2(new_n1001), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n996), .A2(new_n715), .A3(new_n998), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1000), .A2(new_n779), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n994), .B1(new_n1005), .B2(new_n779), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n992), .B(new_n993), .C1(new_n1006), .C2(new_n786), .ZN(new_n1007));
  AND3_X1   g0807(.A1(new_n239), .A2(new_n212), .A3(new_n328), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n804), .B1(new_n338), .B2(new_n212), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n787), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n826), .A2(new_n813), .B1(new_n817), .B2(new_n881), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n265), .B(new_n1011), .C1(G97), .C2(new_n841), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n824), .A2(G107), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n809), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(G116), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT46), .ZN(new_n1016));
  INV_X1    g0816(.A(G317), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n829), .A2(new_n512), .B1(new_n831), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G283), .B2(new_n877), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1012), .A2(new_n1013), .A3(new_n1016), .A4(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n809), .A2(new_n224), .B1(new_n818), .B2(new_n340), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n328), .B(new_n1021), .C1(G159), .C2(new_n875), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n830), .A2(G150), .B1(new_n877), .B2(new_n201), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n827), .A2(G143), .B1(new_n832), .B2(G137), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n823), .A2(new_n218), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1020), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT47), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1010), .B1(new_n1029), .B2(new_n803), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n984), .B2(new_n848), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1007), .A2(new_n1031), .ZN(G387));
  OR2_X1    g0832(.A1(new_n714), .A2(new_n848), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n235), .A2(new_n797), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n1034), .A2(new_n795), .B1(new_n726), .B2(new_n791), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n290), .A2(G50), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  AOI21_X1  g0837(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n726), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1035), .A2(new_n1039), .B1(new_n536), .B2(new_n723), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n787), .B1(new_n1040), .B2(new_n805), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n809), .A2(new_n340), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n826), .A2(new_n838), .B1(new_n817), .B2(new_n290), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(G68), .C2(new_n877), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n829), .A2(new_n443), .B1(new_n831), .B2(new_n867), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n328), .B(new_n1045), .C1(G97), .C2(new_n841), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n338), .A2(new_n823), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n265), .B1(new_n832), .B2(G326), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G322), .A2(new_n827), .B1(new_n875), .B2(G311), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n512), .B2(new_n812), .C1(new_n1017), .C2(new_n829), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT112), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n824), .A2(G283), .B1(new_n1014), .B2(G294), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1049), .B1(new_n480), .B2(new_n818), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1048), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1041), .B1(new_n1061), .B2(new_n803), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1003), .A2(new_n786), .B1(new_n1033), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1003), .A2(new_n779), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n724), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1003), .A2(new_n779), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(G393));
  INV_X1    g0867(.A(new_n1004), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n715), .B1(new_n996), .B2(new_n998), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1064), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n1005), .A3(new_n724), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n804), .B1(new_n226), .B2(new_n212), .C1(new_n246), .C2(new_n795), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n328), .B1(new_n818), .B2(new_n536), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G303), .A2(new_n875), .B1(new_n832), .B2(G322), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n819), .B2(new_n809), .C1(new_n881), .C2(new_n812), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(G116), .C2(new_n824), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n829), .A2(new_n813), .B1(new_n826), .B2(new_n1017), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT52), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n829), .A2(new_n838), .B1(new_n826), .B2(new_n867), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT51), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n218), .A2(new_n809), .B1(new_n812), .B2(new_n290), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n201), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1082), .A2(new_n817), .B1(new_n831), .B2(new_n870), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n823), .A2(new_n340), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n265), .B1(new_n818), .B2(new_n220), .ZN(new_n1085));
  NOR4_X1   g0885(.A1(new_n1081), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1076), .A2(new_n1078), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n803), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n787), .B(new_n1072), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n974), .B2(new_n802), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n786), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1071), .A2(new_n1092), .ZN(G390));
  OAI211_X1 g0893(.A(new_n707), .B(new_n856), .C1(new_n738), .C2(new_n749), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n940), .B1(new_n1094), .B2(new_n942), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n949), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n931), .B2(new_n911), .ZN(new_n1097));
  OAI21_X1  g0897(.A(KEYINPUT113), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n957), .A2(new_n949), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT113), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n683), .A2(new_n597), .A3(new_n644), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n969), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n980), .B1(new_n1102), .B2(new_n747), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n733), .A2(new_n689), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT100), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(new_n735), .A3(new_n734), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n720), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n941), .B1(new_n1108), .B2(new_n856), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1099), .B(new_n1100), .C1(new_n1109), .C2(new_n940), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1098), .A2(new_n1110), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n943), .A2(new_n949), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n948), .B1(new_n957), .B2(KEYINPUT39), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n778), .A2(G330), .A3(new_n856), .A4(new_n939), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1111), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1098), .A2(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n916), .A2(new_n921), .A3(G330), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1113), .A2(new_n800), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n328), .B1(new_n809), .B2(new_n220), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT118), .Z(new_n1123));
  AOI22_X1  g0923(.A1(new_n830), .A2(G116), .B1(new_n877), .B2(G97), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n827), .A2(G283), .B1(new_n832), .B2(G294), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n817), .A2(new_n536), .B1(new_n818), .B2(new_n218), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1126), .A2(new_n1084), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(G128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n829), .A2(new_n863), .B1(new_n826), .B2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT117), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n866), .A2(new_n817), .B1(new_n812), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G159), .B2(new_n824), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n809), .A2(new_n867), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(G125), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n265), .B1(new_n831), .B2(new_n1138), .C1(new_n1082), .C2(new_n818), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT116), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1128), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1141), .A2(new_n803), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n788), .B(new_n1142), .C1(new_n290), .C2(new_n886), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1120), .A2(new_n786), .B1(new_n1121), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT115), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n916), .A2(G330), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n778), .A2(G330), .A3(new_n856), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1146), .A2(new_n921), .B1(new_n1147), .B2(new_n940), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n857), .A2(new_n942), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1094), .A2(new_n1115), .A3(new_n942), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n916), .A2(G330), .A3(new_n856), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1152), .A2(new_n940), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1148), .A2(new_n1150), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1146), .A2(new_n474), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n961), .A2(new_n672), .A3(new_n1155), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1154), .A2(new_n1156), .A3(KEYINPUT114), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT114), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1119), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1152), .A2(new_n940), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1094), .A2(new_n1115), .A3(new_n942), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1147), .A2(new_n940), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n1118), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1161), .A2(new_n1162), .B1(new_n1164), .B2(new_n1149), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n961), .A2(new_n672), .A3(new_n1155), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1116), .B(new_n1167), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1168));
  AND4_X1   g0968(.A1(new_n1145), .A2(new_n1160), .A3(new_n724), .A4(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n725), .B1(new_n1119), .B2(new_n1159), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1145), .B1(new_n1170), .B2(new_n1168), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1144), .B1(new_n1169), .B2(new_n1171), .ZN(G378));
  AOI21_X1  g0972(.A(new_n703), .B1(new_n312), .B2(new_n308), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n322), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1173), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n305), .B(new_n1175), .C1(new_n320), .C2(new_n321), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1177), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT40), .B1(new_n957), .B2(new_n922), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n946), .A2(new_n899), .A3(new_n916), .A4(new_n921), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1181), .B1(new_n1184), .B2(G330), .ZN(new_n1185));
  INV_X1    g0985(.A(G330), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1186), .B(new_n1180), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n960), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1180), .B1(new_n933), .B2(new_n1186), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n947), .A2(new_n958), .A3(new_n959), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1184), .A2(G330), .A3(new_n1181), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1193), .A2(KEYINPUT57), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1168), .A2(new_n1156), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n725), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1188), .A2(new_n1192), .A3(KEYINPUT119), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT119), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1198), .B(new_n960), .C1(new_n1185), .C2(new_n1187), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1195), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1196), .B1(new_n1201), .B2(KEYINPUT120), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT120), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1203), .B(KEYINPUT57), .C1(new_n1200), .C2(new_n1195), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1200), .A2(new_n786), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n788), .B1(new_n1082), .B2(new_n886), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n829), .A2(new_n1129), .B1(new_n817), .B2(new_n863), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G125), .A2(new_n827), .B1(new_n877), .B2(G137), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n809), .B2(new_n1132), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(G150), .C2(new_n824), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT59), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n282), .B(new_n252), .C1(new_n818), .C2(new_n838), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G124), .B2(new_n832), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G58), .A2(new_n841), .B1(new_n832), .B2(G283), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n480), .B2(new_n826), .C1(new_n338), .C2(new_n812), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n328), .A2(new_n252), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1042), .A2(new_n1220), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n829), .A2(new_n536), .B1(new_n817), .B2(new_n226), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(new_n1219), .A2(new_n1025), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT58), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1220), .B(new_n443), .C1(G33), .C2(G41), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1223), .A2(KEYINPUT58), .ZN(new_n1226));
  AND4_X1   g1026(.A1(new_n1217), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1207), .B1(new_n1088), .B2(new_n1227), .C1(new_n1181), .C2(new_n801), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1206), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1205), .A2(new_n1229), .ZN(G375));
  INV_X1    g1030(.A(new_n994), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1159), .B(new_n1231), .C1(new_n1156), .C2(new_n1154), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n940), .A2(new_n800), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n829), .A2(new_n819), .B1(new_n826), .B2(new_n881), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n265), .B(new_n1234), .C1(G77), .C2(new_n841), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G97), .A2(new_n1014), .B1(new_n875), .B2(G116), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G107), .A2(new_n877), .B1(new_n832), .B2(G303), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1235), .A2(new_n1047), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n809), .A2(new_n838), .B1(new_n831), .B2(new_n1129), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n328), .B(new_n1239), .C1(G58), .C2(new_n841), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n826), .A2(new_n863), .B1(new_n817), .B2(new_n1132), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n829), .A2(new_n866), .B1(new_n812), .B2(new_n867), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1240), .B(new_n1243), .C1(new_n443), .C2(new_n823), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1088), .B1(new_n1238), .B2(new_n1244), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n788), .B(new_n1245), .C1(new_n218), .C2(new_n886), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1154), .A2(new_n786), .B1(new_n1233), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1232), .A2(new_n1247), .ZN(G381));
  INV_X1    g1048(.A(KEYINPUT121), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(G375), .B(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1170), .A2(new_n1168), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1251), .A2(new_n1144), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OR4_X1    g1053(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1254));
  OR3_X1    g1054(.A1(new_n1254), .A2(G387), .A3(G381), .ZN(new_n1255));
  OR3_X1    g1055(.A1(new_n1250), .A2(new_n1253), .A3(new_n1255), .ZN(G407));
  NAND2_X1  g1056(.A1(new_n705), .A2(G213), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1252), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G407), .B(G213), .C1(new_n1250), .C2(new_n1259), .ZN(G409));
  INV_X1    g1060(.A(KEYINPUT61), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G378), .B(new_n1229), .C1(new_n1202), .C2(new_n1204), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1200), .A2(new_n1231), .A3(new_n1195), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1193), .A2(new_n786), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1228), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1252), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1258), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT123), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1164), .A2(new_n1149), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1109), .A2(new_n1161), .A3(new_n1115), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1269), .A2(new_n1166), .A3(KEYINPUT60), .A4(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT122), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1165), .A2(KEYINPUT122), .A3(KEYINPUT60), .A4(new_n1166), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n725), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1273), .A2(new_n1274), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1278), .A2(G384), .A3(new_n1247), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1278), .B2(new_n1247), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1268), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1247), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1278), .A2(G384), .A3(new_n1247), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(KEYINPUT123), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1281), .A2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(KEYINPUT125), .A2(G2897), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1257), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1257), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1287), .B2(KEYINPUT125), .ZN(new_n1291));
  INV_X1    g1091(.A(G2897), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1289), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1261), .B1(new_n1267), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(KEYINPUT127), .B(new_n1261), .C1(new_n1267), .C2(new_n1293), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1267), .A2(new_n1287), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT62), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1267), .A2(new_n1300), .A3(new_n1287), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1296), .A2(new_n1297), .A3(new_n1299), .A4(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(G390), .B1(new_n1007), .B2(new_n1031), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1007), .A2(new_n1031), .A3(G390), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  XOR2_X1   g1106(.A(G396), .B(G393), .Z(new_n1307));
  OAI21_X1  g1107(.A(new_n1307), .B1(new_n1303), .B2(KEYINPUT126), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1304), .A2(KEYINPUT126), .A3(new_n1305), .A4(new_n1307), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1302), .A2(new_n1311), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1267), .A2(new_n1287), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1311), .B1(new_n1313), .B2(KEYINPUT63), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1294), .ZN(new_n1315));
  AOI211_X1 g1115(.A(KEYINPUT124), .B(KEYINPUT63), .C1(new_n1267), .C2(new_n1287), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT124), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT63), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1298), .B2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1314), .B(new_n1315), .C1(new_n1316), .C2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1312), .A2(new_n1320), .ZN(G405));
  INV_X1    g1121(.A(G375), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1262), .B1(new_n1322), .B2(new_n1253), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1287), .ZN(new_n1324));
  OAI221_X1 g1124(.A(new_n1262), .B1(new_n1280), .B2(new_n1279), .C1(new_n1322), .C2(new_n1253), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1324), .A2(new_n1311), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1311), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(G402));
endmodule


