

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n364, n365, n366, n367, n368, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792;

  XNOR2_X1 U385 ( .A(n646), .B(KEYINPUT32), .ZN(n788) );
  INV_X1 U386 ( .A(n598), .ZN(n688) );
  AND2_X1 U387 ( .A1(n452), .A2(n451), .ZN(n585) );
  NOR2_X1 U388 ( .A1(n596), .A2(n464), .ZN(n582) );
  AND2_X1 U389 ( .A1(n365), .A2(n427), .ZN(n426) );
  OR2_X1 U390 ( .A1(n758), .A2(G902), .ZN(n479) );
  XNOR2_X1 U391 ( .A(n549), .B(n548), .ZN(n760) );
  XNOR2_X1 U392 ( .A(n364), .B(n546), .ZN(n549) );
  XNOR2_X1 U393 ( .A(n574), .B(n543), .ZN(n364) );
  INV_X1 U394 ( .A(G143), .ZN(n503) );
  NAND2_X4 U395 ( .A1(n426), .A2(n424), .ZN(n400) );
  INV_X1 U396 ( .A(G953), .ZN(n784) );
  AND2_X2 U397 ( .A1(n715), .A2(n716), .ZN(n442) );
  AND2_X2 U398 ( .A1(n446), .A2(n640), .ZN(n379) );
  AND2_X2 U399 ( .A1(n416), .A2(n457), .ZN(n402) );
  XNOR2_X2 U400 ( .A(n554), .B(n495), .ZN(n521) );
  XNOR2_X2 U401 ( .A(n367), .B(KEYINPUT42), .ZN(n792) );
  XNOR2_X2 U402 ( .A(n400), .B(KEYINPUT104), .ZN(n467) );
  XNOR2_X2 U403 ( .A(n777), .B(G101), .ZN(n554) );
  AND2_X1 U404 ( .A1(n423), .A2(n422), .ZN(n421) );
  NAND2_X1 U405 ( .A1(n415), .A2(KEYINPUT0), .ZN(n414) );
  NAND2_X2 U406 ( .A1(n371), .A2(n716), .ZN(n398) );
  INV_X1 U407 ( .A(G146), .ZN(n495) );
  NAND2_X1 U408 ( .A1(n421), .A2(n418), .ZN(n417) );
  NAND2_X1 U409 ( .A1(n402), .A2(n414), .ZN(n622) );
  AND2_X1 U410 ( .A1(n414), .A2(n449), .ZN(n383) );
  XNOR2_X1 U411 ( .A(n538), .B(n539), .ZN(n478) );
  XNOR2_X1 U412 ( .A(n760), .B(n556), .ZN(n666) );
  XNOR2_X1 U413 ( .A(n495), .B(G125), .ZN(n550) );
  NAND2_X1 U414 ( .A1(n672), .A2(n373), .ZN(n365) );
  XNOR2_X2 U415 ( .A(n521), .B(n514), .ZN(n672) );
  XNOR2_X1 U416 ( .A(n366), .B(n475), .ZN(n471) );
  NAND2_X1 U417 ( .A1(n791), .A2(n792), .ZN(n366) );
  NAND2_X1 U418 ( .A1(n713), .A2(n585), .ZN(n367) );
  XNOR2_X2 U419 ( .A(n368), .B(KEYINPUT40), .ZN(n791) );
  NAND2_X1 U420 ( .A1(n605), .A2(n690), .ZN(n368) );
  XNOR2_X2 U421 ( .A(n370), .B(G122), .ZN(n574) );
  XNOR2_X2 U422 ( .A(G113), .B(G104), .ZN(n370) );
  INV_X1 U423 ( .A(n371), .ZN(n592) );
  XNOR2_X2 U424 ( .A(n455), .B(n384), .ZN(n371) );
  NOR2_X1 U425 ( .A1(n612), .A2(n401), .ZN(n613) );
  AND2_X1 U426 ( .A1(n372), .A2(n442), .ZN(n721) );
  INV_X1 U427 ( .A(n720), .ZN(n372) );
  OR2_X2 U428 ( .A1(n650), .A2(KEYINPUT44), .ZN(n381) );
  XNOR2_X2 U429 ( .A(n563), .B(n504), .ZN(n777) );
  AND2_X1 U430 ( .A1(n638), .A2(KEYINPUT64), .ZN(n481) );
  XNOR2_X1 U431 ( .A(n583), .B(n441), .ZN(n619) );
  INV_X1 U432 ( .A(KEYINPUT103), .ZN(n441) );
  AND2_X1 U433 ( .A1(n590), .A2(n589), .ZN(n583) );
  XNOR2_X1 U434 ( .A(n374), .B(n553), .ZN(n555) );
  AND2_X1 U435 ( .A1(n470), .A2(n602), .ZN(n472) );
  INV_X1 U436 ( .A(KEYINPUT89), .ZN(n489) );
  NAND2_X1 U437 ( .A1(n412), .A2(KEYINPUT111), .ZN(n411) );
  INV_X1 U438 ( .A(KEYINPUT45), .ZN(n448) );
  OR2_X1 U439 ( .A1(G237), .A2(G902), .ZN(n557) );
  XNOR2_X1 U440 ( .A(G902), .B(KEYINPUT15), .ZN(n536) );
  OR2_X1 U441 ( .A1(n749), .A2(G902), .ZN(n447) );
  OR2_X1 U442 ( .A1(n672), .A2(n425), .ZN(n424) );
  OR2_X1 U443 ( .A1(n373), .A2(G902), .ZN(n425) );
  XNOR2_X1 U444 ( .A(G137), .B(G116), .ZN(n507) );
  XOR2_X1 U445 ( .A(G119), .B(G113), .Z(n508) );
  XOR2_X1 U446 ( .A(KEYINPUT98), .B(KEYINPUT5), .Z(n506) );
  XNOR2_X1 U447 ( .A(n511), .B(KEYINPUT69), .ZN(n516) );
  XNOR2_X1 U448 ( .A(n550), .B(n477), .ZN(n774) );
  XNOR2_X1 U449 ( .A(KEYINPUT10), .B(G140), .ZN(n477) );
  XNOR2_X1 U450 ( .A(G128), .B(KEYINPUT86), .ZN(n524) );
  XOR2_X1 U451 ( .A(KEYINPUT78), .B(KEYINPUT96), .Z(n526) );
  XOR2_X1 U452 ( .A(G116), .B(G107), .Z(n564) );
  XNOR2_X1 U453 ( .A(n530), .B(n531), .ZN(n561) );
  XNOR2_X1 U454 ( .A(KEYINPUT87), .B(KEYINPUT8), .ZN(n530) );
  XNOR2_X1 U455 ( .A(n562), .B(n392), .ZN(n391) );
  XNOR2_X1 U456 ( .A(G122), .B(KEYINPUT7), .ZN(n392) );
  XOR2_X1 U457 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n562) );
  XNOR2_X1 U458 ( .A(n516), .B(n529), .ZN(n494) );
  INV_X1 U459 ( .A(n579), .ZN(n437) );
  INV_X1 U460 ( .A(n592), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n394), .B(n403), .ZN(n590) );
  INV_X1 U462 ( .A(G478), .ZN(n403) );
  OR2_X1 U463 ( .A1(n754), .A2(G902), .ZN(n394) );
  AND2_X1 U464 ( .A1(n619), .A2(n580), .ZN(n449) );
  XNOR2_X1 U465 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U466 ( .A1(n395), .A2(n433), .ZN(n476) );
  XNOR2_X1 U467 ( .A(n397), .B(n396), .ZN(n395) );
  INV_X1 U468 ( .A(KEYINPUT36), .ZN(n396) );
  INV_X1 U469 ( .A(KEYINPUT46), .ZN(n475) );
  NOR2_X1 U470 ( .A1(n496), .A2(n603), .ZN(n470) );
  NAND2_X1 U471 ( .A1(n382), .A2(n476), .ZN(n473) );
  NAND2_X1 U472 ( .A1(n373), .A2(G902), .ZN(n427) );
  NOR2_X1 U473 ( .A1(G953), .A2(G237), .ZN(n567) );
  INV_X1 U474 ( .A(KEYINPUT16), .ZN(n544) );
  XOR2_X1 U475 ( .A(G131), .B(KEYINPUT11), .Z(n569) );
  XNOR2_X1 U476 ( .A(G143), .B(KEYINPUT12), .ZN(n570) );
  XOR2_X1 U477 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n571) );
  NAND2_X1 U478 ( .A1(n490), .A2(n489), .ZN(n488) );
  XNOR2_X1 U479 ( .A(KEYINPUT95), .B(KEYINPUT79), .ZN(n552) );
  NAND2_X1 U480 ( .A1(G234), .A2(G237), .ZN(n498) );
  INV_X1 U481 ( .A(KEYINPUT30), .ZN(n434) );
  AND2_X1 U482 ( .A1(n411), .A2(n410), .ZN(n409) );
  BUF_X1 U483 ( .A(n464), .Z(n450) );
  XNOR2_X1 U484 ( .A(n595), .B(n594), .ZN(n701) );
  BUF_X1 U485 ( .A(n735), .Z(n782) );
  INV_X1 U486 ( .A(n494), .ZN(n773) );
  NOR2_X1 U487 ( .A1(n597), .A2(n596), .ZN(n404) );
  XNOR2_X1 U488 ( .A(KEYINPUT81), .B(KEYINPUT34), .ZN(n631) );
  NAND2_X1 U489 ( .A1(n463), .A2(KEYINPUT65), .ZN(n462) );
  NAND2_X1 U490 ( .A1(n465), .A2(n450), .ZN(n463) );
  NAND2_X1 U491 ( .A1(n460), .A2(n450), .ZN(n459) );
  NOR2_X1 U492 ( .A1(n433), .A2(KEYINPUT65), .ZN(n460) );
  XNOR2_X1 U493 ( .A(n577), .B(n440), .ZN(n589) );
  XNOR2_X1 U494 ( .A(n578), .B(G475), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n528), .B(n774), .ZN(n535) );
  XNOR2_X1 U496 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U497 ( .A(n566), .B(n565), .ZN(n754) );
  XNOR2_X1 U498 ( .A(n390), .B(n389), .ZN(n566) );
  AND2_X1 U499 ( .A1(n561), .A2(G217), .ZN(n389) );
  XNOR2_X1 U500 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U501 ( .A(n521), .B(n405), .ZN(n749) );
  XNOR2_X1 U502 ( .A(n494), .B(n520), .ZN(n405) );
  XOR2_X1 U503 ( .A(G110), .B(G140), .Z(n497) );
  INV_X1 U504 ( .A(KEYINPUT112), .ZN(n453) );
  AND2_X1 U505 ( .A1(n590), .A2(n393), .ZN(n690) );
  INV_X1 U506 ( .A(n589), .ZN(n393) );
  INV_X1 U507 ( .A(KEYINPUT56), .ZN(n443) );
  INV_X1 U508 ( .A(n476), .ZN(n697) );
  INV_X1 U509 ( .A(n433), .ZN(n465) );
  XNOR2_X1 U510 ( .A(G472), .B(KEYINPUT74), .ZN(n373) );
  XOR2_X1 U511 ( .A(n551), .B(n550), .Z(n374) );
  OR2_X1 U512 ( .A1(n699), .A2(n790), .ZN(n375) );
  XNOR2_X1 U513 ( .A(n541), .B(KEYINPUT21), .ZN(n704) );
  XOR2_X1 U514 ( .A(n508), .B(n507), .Z(n376) );
  XOR2_X1 U515 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n377) );
  AND2_X1 U516 ( .A1(n559), .A2(n401), .ZN(n378) );
  OR2_X2 U517 ( .A1(n703), .A2(n704), .ZN(n412) );
  NOR2_X1 U518 ( .A1(n641), .A2(n433), .ZN(n380) );
  OR2_X1 U519 ( .A1(n720), .A2(n601), .ZN(n382) );
  INV_X1 U520 ( .A(n642), .ZN(n629) );
  XOR2_X1 U521 ( .A(n558), .B(KEYINPUT82), .Z(n384) );
  XOR2_X1 U522 ( .A(KEYINPUT113), .B(KEYINPUT41), .Z(n385) );
  XNOR2_X1 U523 ( .A(n536), .B(KEYINPUT94), .ZN(n386) );
  OR2_X1 U524 ( .A1(n738), .A2(n386), .ZN(n387) );
  XOR2_X1 U525 ( .A(KEYINPUT93), .B(n662), .Z(n759) );
  INV_X1 U526 ( .A(n759), .ZN(n675) );
  NAND2_X1 U527 ( .A1(n383), .A2(n402), .ZN(n620) );
  INV_X1 U528 ( .A(n622), .ZN(n388) );
  NAND2_X1 U529 ( .A1(n388), .A2(n624), .ZN(n625) );
  NAND2_X1 U530 ( .A1(n724), .A2(n388), .ZN(n632) );
  XNOR2_X1 U531 ( .A(n391), .B(n563), .ZN(n390) );
  XNOR2_X2 U532 ( .A(n503), .B(G128), .ZN(n563) );
  INV_X1 U533 ( .A(n590), .ZN(n586) );
  XNOR2_X2 U534 ( .A(n398), .B(KEYINPUT19), .ZN(n584) );
  OR2_X1 U535 ( .A1(n607), .A2(n398), .ZN(n397) );
  INV_X1 U536 ( .A(n400), .ZN(n624) );
  XNOR2_X1 U537 ( .A(n400), .B(n399), .ZN(n642) );
  INV_X1 U538 ( .A(KEYINPUT6), .ZN(n399) );
  NOR2_X1 U539 ( .A1(n707), .A2(n400), .ZN(n708) );
  AND2_X2 U540 ( .A1(n438), .A2(n436), .ZN(n559) );
  NAND2_X1 U541 ( .A1(n666), .A2(n386), .ZN(n455) );
  XNOR2_X1 U542 ( .A(n560), .B(KEYINPUT39), .ZN(n605) );
  XNOR2_X2 U543 ( .A(n592), .B(KEYINPUT38), .ZN(n715) );
  NAND2_X1 U544 ( .A1(n442), .A2(n619), .ZN(n431) );
  OR2_X1 U545 ( .A1(n461), .A2(n458), .ZN(n647) );
  XNOR2_X1 U546 ( .A(n404), .B(KEYINPUT107), .ZN(n607) );
  NAND2_X1 U547 ( .A1(n420), .A2(n419), .ZN(n418) );
  NAND2_X1 U548 ( .A1(n408), .A2(n451), .ZN(n626) );
  NAND2_X1 U549 ( .A1(n409), .A2(n406), .ZN(n542) );
  NAND2_X1 U550 ( .A1(n408), .A2(n407), .ZN(n406) );
  NOR2_X1 U551 ( .A1(n595), .A2(KEYINPUT111), .ZN(n407) );
  INV_X2 U552 ( .A(n412), .ZN(n408) );
  NAND2_X1 U553 ( .A1(n595), .A2(KEYINPUT111), .ZN(n410) );
  XNOR2_X2 U554 ( .A(n479), .B(n478), .ZN(n703) );
  XNOR2_X2 U555 ( .A(n447), .B(n522), .ZN(n595) );
  XNOR2_X1 U556 ( .A(n413), .B(n614), .ZN(n735) );
  NAND2_X1 U557 ( .A1(n655), .A2(n413), .ZN(n739) );
  NOR2_X2 U558 ( .A1(n417), .A2(n375), .ZN(n413) );
  NAND2_X1 U559 ( .A1(n467), .A2(n716), .ZN(n515) );
  INV_X1 U560 ( .A(n584), .ZN(n415) );
  NAND2_X1 U561 ( .A1(n584), .A2(n456), .ZN(n416) );
  NOR2_X1 U562 ( .A1(n473), .A2(n604), .ZN(n419) );
  INV_X1 U563 ( .A(n474), .ZN(n420) );
  NAND2_X1 U564 ( .A1(n473), .A2(n604), .ZN(n422) );
  NAND2_X1 U565 ( .A1(n474), .A2(n604), .ZN(n423) );
  NAND2_X1 U566 ( .A1(n428), .A2(n675), .ZN(n432) );
  XNOR2_X1 U567 ( .A(n673), .B(n674), .ZN(n428) );
  NAND2_X1 U568 ( .A1(n482), .A2(n481), .ZN(n469) );
  XNOR2_X1 U569 ( .A(n515), .B(n434), .ZN(n438) );
  AND2_X1 U570 ( .A1(n429), .A2(n675), .ZN(G66) );
  XNOR2_X1 U571 ( .A(n757), .B(n430), .ZN(n429) );
  INV_X1 U572 ( .A(n758), .ZN(n430) );
  XNOR2_X2 U573 ( .A(n431), .B(n385), .ZN(n713) );
  NAND2_X1 U574 ( .A1(n788), .A2(n683), .ZN(n649) );
  NAND2_X1 U575 ( .A1(n671), .A2(n675), .ZN(n444) );
  XNOR2_X1 U576 ( .A(n432), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U577 ( .A(n376), .B(n509), .ZN(n513) );
  AND2_X1 U578 ( .A1(n484), .A2(n387), .ZN(n492) );
  XNOR2_X1 U579 ( .A(n444), .B(n443), .ZN(G51) );
  BUF_X1 U580 ( .A(n701), .Z(n433) );
  AND2_X1 U581 ( .A1(n542), .A2(n437), .ZN(n436) );
  NAND2_X1 U582 ( .A1(n559), .A2(n715), .ZN(n560) );
  XNOR2_X1 U583 ( .A(n649), .B(KEYINPUT64), .ZN(n651) );
  XNOR2_X1 U584 ( .A(n582), .B(KEYINPUT28), .ZN(n452) );
  INV_X1 U585 ( .A(n467), .ZN(n464) );
  NAND2_X2 U586 ( .A1(n435), .A2(n468), .ZN(n653) );
  AND2_X2 U587 ( .A1(n379), .A2(n652), .ZN(n435) );
  NOR2_X1 U588 ( .A1(n491), .A2(n439), .ZN(n657) );
  AND2_X2 U589 ( .A1(n485), .A2(KEYINPUT89), .ZN(n439) );
  NOR2_X2 U590 ( .A1(n633), .A2(n593), .ZN(n687) );
  NAND2_X1 U591 ( .A1(n471), .A2(n472), .ZN(n474) );
  INV_X1 U592 ( .A(n619), .ZN(n718) );
  XNOR2_X2 U593 ( .A(n445), .B(KEYINPUT33), .ZN(n724) );
  NAND2_X1 U594 ( .A1(n483), .A2(n642), .ZN(n445) );
  NAND2_X1 U595 ( .A1(n454), .A2(n639), .ZN(n446) );
  NAND2_X1 U596 ( .A1(n469), .A2(n480), .ZN(n468) );
  INV_X1 U597 ( .A(n654), .ZN(n655) );
  NAND2_X1 U598 ( .A1(n654), .A2(KEYINPUT89), .ZN(n484) );
  XNOR2_X2 U599 ( .A(n653), .B(n448), .ZN(n654) );
  INV_X1 U600 ( .A(n595), .ZN(n451) );
  XNOR2_X1 U601 ( .A(n378), .B(n453), .ZN(n593) );
  NAND2_X1 U602 ( .A1(n637), .A2(n638), .ZN(n454) );
  INV_X1 U603 ( .A(n630), .ZN(n483) );
  NAND2_X1 U604 ( .A1(n701), .A2(n408), .ZN(n630) );
  NOR2_X1 U605 ( .A1(n618), .A2(KEYINPUT0), .ZN(n456) );
  NAND2_X1 U606 ( .A1(n618), .A2(KEYINPUT0), .ZN(n457) );
  NOR2_X1 U607 ( .A1(n641), .A2(n459), .ZN(n458) );
  NAND2_X1 U608 ( .A1(n466), .A2(n462), .ZN(n461) );
  NAND2_X1 U609 ( .A1(n641), .A2(KEYINPUT65), .ZN(n466) );
  XNOR2_X2 U610 ( .A(n620), .B(KEYINPUT22), .ZN(n641) );
  INV_X1 U611 ( .A(KEYINPUT44), .ZN(n480) );
  NAND2_X1 U612 ( .A1(n648), .A2(KEYINPUT92), .ZN(n482) );
  OR2_X2 U613 ( .A1(n735), .A2(n386), .ZN(n485) );
  NAND2_X1 U614 ( .A1(n487), .A2(n486), .ZN(n493) );
  INV_X1 U615 ( .A(n735), .ZN(n486) );
  NOR2_X1 U616 ( .A1(n654), .A2(n488), .ZN(n487) );
  INV_X1 U617 ( .A(n386), .ZN(n490) );
  NAND2_X1 U618 ( .A1(n493), .A2(n492), .ZN(n491) );
  XNOR2_X1 U619 ( .A(n751), .B(n750), .ZN(n752) );
  NAND2_X1 U620 ( .A1(n663), .A2(n675), .ZN(n665) );
  XNOR2_X1 U621 ( .A(n749), .B(n748), .ZN(n750) );
  XNOR2_X1 U622 ( .A(n554), .B(n555), .ZN(n556) );
  AND2_X1 U623 ( .A1(KEYINPUT47), .A2(n588), .ZN(n496) );
  XNOR2_X1 U624 ( .A(n545), .B(n544), .ZN(n546) );
  INV_X1 U625 ( .A(n607), .ZN(n608) );
  INV_X1 U626 ( .A(KEYINPUT4), .ZN(n504) );
  XNOR2_X1 U627 ( .A(n519), .B(n497), .ZN(n520) );
  XNOR2_X1 U628 ( .A(n661), .B(n660), .ZN(n663) );
  INV_X1 U629 ( .A(KEYINPUT60), .ZN(n664) );
  XNOR2_X1 U630 ( .A(KEYINPUT48), .B(KEYINPUT70), .ZN(n604) );
  NOR2_X1 U631 ( .A1(KEYINPUT84), .A2(KEYINPUT47), .ZN(n603) );
  XNOR2_X1 U632 ( .A(n498), .B(KEYINPUT14), .ZN(n499) );
  NAND2_X1 U633 ( .A1(G952), .A2(n499), .ZN(n700) );
  NOR2_X1 U634 ( .A1(G953), .A2(n700), .ZN(n617) );
  NAND2_X1 U635 ( .A1(G902), .A2(n499), .ZN(n615) );
  NOR2_X1 U636 ( .A1(G900), .A2(n615), .ZN(n500) );
  NAND2_X1 U637 ( .A1(G953), .A2(n500), .ZN(n501) );
  XOR2_X1 U638 ( .A(KEYINPUT106), .B(n501), .Z(n502) );
  NOR2_X1 U639 ( .A1(n617), .A2(n502), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n567), .A2(G210), .ZN(n505) );
  XNOR2_X1 U641 ( .A(n506), .B(n505), .ZN(n509) );
  XNOR2_X1 U642 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n510) );
  XNOR2_X1 U643 ( .A(n510), .B(KEYINPUT73), .ZN(n547) );
  XNOR2_X1 U644 ( .A(G131), .B(G134), .ZN(n511) );
  XNOR2_X1 U645 ( .A(n516), .B(n547), .ZN(n512) );
  XNOR2_X1 U646 ( .A(n513), .B(n512), .ZN(n514) );
  NAND2_X1 U647 ( .A1(G214), .A2(n557), .ZN(n716) );
  XOR2_X1 U648 ( .A(G137), .B(KEYINPUT68), .Z(n529) );
  XOR2_X1 U649 ( .A(G104), .B(G107), .Z(n518) );
  NAND2_X1 U650 ( .A1(G227), .A2(n784), .ZN(n517) );
  XNOR2_X1 U651 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U652 ( .A(KEYINPUT71), .B(G469), .ZN(n522) );
  XNOR2_X1 U653 ( .A(KEYINPUT25), .B(KEYINPUT97), .ZN(n523) );
  XNOR2_X1 U654 ( .A(n523), .B(KEYINPUT77), .ZN(n539) );
  XOR2_X1 U655 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n525) );
  XNOR2_X1 U656 ( .A(n525), .B(n524), .ZN(n527) );
  XOR2_X1 U657 ( .A(G119), .B(G110), .Z(n543) );
  XOR2_X1 U658 ( .A(n543), .B(n529), .Z(n533) );
  NAND2_X1 U659 ( .A1(n784), .A2(G234), .ZN(n531) );
  NAND2_X1 U660 ( .A1(G221), .A2(n561), .ZN(n532) );
  XNOR2_X1 U661 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U662 ( .A(n535), .B(n534), .ZN(n758) );
  NAND2_X1 U663 ( .A1(G234), .A2(n386), .ZN(n537) );
  XNOR2_X1 U664 ( .A(n537), .B(KEYINPUT20), .ZN(n540) );
  NAND2_X1 U665 ( .A1(n540), .A2(G217), .ZN(n538) );
  NAND2_X1 U666 ( .A1(G221), .A2(n540), .ZN(n541) );
  XOR2_X1 U667 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n545) );
  XNOR2_X1 U668 ( .A(n547), .B(n564), .ZN(n548) );
  NAND2_X1 U669 ( .A1(G224), .A2(n784), .ZN(n551) );
  XNOR2_X1 U670 ( .A(n377), .B(n552), .ZN(n553) );
  NAND2_X1 U671 ( .A1(G210), .A2(n557), .ZN(n558) );
  XNOR2_X1 U672 ( .A(G134), .B(n564), .ZN(n565) );
  XNOR2_X1 U673 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n578) );
  NAND2_X1 U674 ( .A1(G214), .A2(n567), .ZN(n568) );
  XNOR2_X1 U675 ( .A(n569), .B(n568), .ZN(n573) );
  XNOR2_X1 U676 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U677 ( .A(n573), .B(n572), .Z(n576) );
  XNOR2_X1 U678 ( .A(n774), .B(n574), .ZN(n575) );
  XNOR2_X1 U679 ( .A(n576), .B(n575), .ZN(n659) );
  NOR2_X1 U680 ( .A1(G902), .A2(n659), .ZN(n577) );
  INV_X1 U681 ( .A(n703), .ZN(n643) );
  NOR2_X1 U682 ( .A1(n579), .A2(n643), .ZN(n581) );
  INV_X1 U683 ( .A(n704), .ZN(n580) );
  NAND2_X1 U684 ( .A1(n581), .A2(n580), .ZN(n596) );
  NAND2_X1 U685 ( .A1(n585), .A2(n584), .ZN(n598) );
  AND2_X1 U686 ( .A1(n589), .A2(n586), .ZN(n692) );
  NOR2_X1 U687 ( .A1(n690), .A2(n692), .ZN(n720) );
  NAND2_X1 U688 ( .A1(KEYINPUT84), .A2(n720), .ZN(n587) );
  NAND2_X1 U689 ( .A1(n688), .A2(n587), .ZN(n588) );
  NOR2_X1 U690 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U691 ( .A(n591), .B(KEYINPUT105), .ZN(n633) );
  XNOR2_X1 U692 ( .A(KEYINPUT85), .B(n687), .ZN(n602) );
  XOR2_X1 U693 ( .A(KEYINPUT1), .B(KEYINPUT66), .Z(n594) );
  NAND2_X1 U694 ( .A1(n690), .A2(n642), .ZN(n597) );
  NOR2_X1 U695 ( .A1(KEYINPUT47), .A2(n598), .ZN(n600) );
  INV_X1 U696 ( .A(KEYINPUT84), .ZN(n599) );
  NOR2_X1 U697 ( .A1(n600), .A2(n599), .ZN(n601) );
  AND2_X1 U698 ( .A1(n605), .A2(n692), .ZN(n699) );
  XOR2_X1 U699 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n606) );
  XNOR2_X1 U700 ( .A(KEYINPUT43), .B(n606), .ZN(n611) );
  NAND2_X1 U701 ( .A1(n608), .A2(n716), .ZN(n609) );
  NOR2_X1 U702 ( .A1(n433), .A2(n609), .ZN(n610) );
  XNOR2_X1 U703 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U704 ( .A(n613), .B(KEYINPUT110), .ZN(n790) );
  INV_X1 U705 ( .A(KEYINPUT90), .ZN(n614) );
  INV_X1 U706 ( .A(G898), .ZN(n768) );
  NAND2_X1 U707 ( .A1(G953), .A2(n768), .ZN(n762) );
  NOR2_X1 U708 ( .A1(n615), .A2(n762), .ZN(n616) );
  NOR2_X1 U709 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U710 ( .A1(n629), .A2(n380), .ZN(n621) );
  NOR2_X1 U711 ( .A1(n703), .A2(n621), .ZN(n676) );
  OR2_X1 U712 ( .A1(n630), .A2(n624), .ZN(n711) );
  NOR2_X1 U713 ( .A1(n711), .A2(n622), .ZN(n623) );
  XOR2_X1 U714 ( .A(KEYINPUT31), .B(n623), .Z(n693) );
  NOR2_X1 U715 ( .A1(n626), .A2(n625), .ZN(n679) );
  NOR2_X1 U716 ( .A1(n693), .A2(n679), .ZN(n627) );
  NOR2_X1 U717 ( .A1(n720), .A2(n627), .ZN(n628) );
  NOR2_X1 U718 ( .A1(n676), .A2(n628), .ZN(n640) );
  INV_X1 U719 ( .A(KEYINPUT91), .ZN(n638) );
  XNOR2_X1 U720 ( .A(n632), .B(n631), .ZN(n635) );
  XOR2_X1 U721 ( .A(n633), .B(KEYINPUT80), .Z(n634) );
  NAND2_X1 U722 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X2 U723 ( .A(n636), .B(KEYINPUT35), .ZN(n787) );
  NAND2_X1 U724 ( .A1(n787), .A2(KEYINPUT44), .ZN(n637) );
  NAND2_X1 U725 ( .A1(n787), .A2(KEYINPUT91), .ZN(n639) );
  NOR2_X1 U726 ( .A1(n641), .A2(n465), .ZN(n645) );
  NOR2_X1 U727 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n647), .A2(n703), .ZN(n683) );
  NOR2_X1 U730 ( .A1(n649), .A2(n787), .ZN(n648) );
  NOR2_X1 U731 ( .A1(n787), .A2(KEYINPUT92), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n651), .A2(n381), .ZN(n652) );
  INV_X1 U733 ( .A(KEYINPUT2), .ZN(n738) );
  NOR2_X1 U734 ( .A1(n738), .A2(n739), .ZN(n656) );
  NOR2_X2 U735 ( .A1(n657), .A2(n656), .ZN(n747) );
  NAND2_X1 U736 ( .A1(n747), .A2(G475), .ZN(n661) );
  XOR2_X1 U737 ( .A(KEYINPUT59), .B(KEYINPUT67), .Z(n658) );
  NOR2_X1 U738 ( .A1(G952), .A2(n784), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n665), .B(n664), .ZN(G60) );
  NAND2_X1 U740 ( .A1(n747), .A2(G210), .ZN(n670) );
  XNOR2_X1 U741 ( .A(KEYINPUT55), .B(KEYINPUT83), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n666), .B(KEYINPUT54), .ZN(n667) );
  XNOR2_X1 U743 ( .A(n670), .B(n669), .ZN(n671) );
  XOR2_X1 U744 ( .A(n672), .B(KEYINPUT62), .Z(n674) );
  NAND2_X1 U745 ( .A1(n747), .A2(G472), .ZN(n673) );
  XOR2_X1 U746 ( .A(G101), .B(n676), .Z(G3) );
  NAND2_X1 U747 ( .A1(n679), .A2(n690), .ZN(n677) );
  XNOR2_X1 U748 ( .A(n677), .B(KEYINPUT114), .ZN(n678) );
  XNOR2_X1 U749 ( .A(G104), .B(n678), .ZN(G6) );
  XOR2_X1 U750 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n681) );
  NAND2_X1 U751 ( .A1(n679), .A2(n692), .ZN(n680) );
  XNOR2_X1 U752 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U753 ( .A(G107), .B(n682), .ZN(G9) );
  BUF_X1 U754 ( .A(n683), .Z(n684) );
  XNOR2_X1 U755 ( .A(G110), .B(n684), .ZN(G12) );
  XOR2_X1 U756 ( .A(G128), .B(KEYINPUT29), .Z(n686) );
  NAND2_X1 U757 ( .A1(n688), .A2(n692), .ZN(n685) );
  XNOR2_X1 U758 ( .A(n686), .B(n685), .ZN(G30) );
  XOR2_X1 U759 ( .A(G143), .B(n687), .Z(G45) );
  NAND2_X1 U760 ( .A1(n688), .A2(n690), .ZN(n689) );
  XNOR2_X1 U761 ( .A(n689), .B(G146), .ZN(G48) );
  NAND2_X1 U762 ( .A1(n693), .A2(n690), .ZN(n691) );
  XNOR2_X1 U763 ( .A(n691), .B(G113), .ZN(G15) );
  XOR2_X1 U764 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n695) );
  NAND2_X1 U765 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U766 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U767 ( .A(G116), .B(n696), .ZN(G18) );
  XNOR2_X1 U768 ( .A(n697), .B(G125), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n698), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U770 ( .A(G134), .B(n699), .Z(G36) );
  NAND2_X1 U771 ( .A1(n713), .A2(n724), .ZN(n733) );
  INV_X1 U772 ( .A(n700), .ZN(n731) );
  NOR2_X1 U773 ( .A1(n433), .A2(n408), .ZN(n702) );
  XOR2_X1 U774 ( .A(KEYINPUT50), .B(n702), .Z(n709) );
  XOR2_X1 U775 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n706) );
  NAND2_X1 U776 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U777 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U778 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U779 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U780 ( .A(KEYINPUT51), .B(n712), .Z(n714) );
  NAND2_X1 U781 ( .A1(n714), .A2(n713), .ZN(n727) );
  NOR2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U784 ( .A(n719), .B(KEYINPUT118), .ZN(n722) );
  NOR2_X1 U785 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U786 ( .A(KEYINPUT119), .B(n723), .ZN(n725) );
  NAND2_X1 U787 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U788 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U789 ( .A(n728), .B(KEYINPUT52), .ZN(n729) );
  XNOR2_X1 U790 ( .A(KEYINPUT120), .B(n729), .ZN(n730) );
  NAND2_X1 U791 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U792 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U793 ( .A(n734), .B(KEYINPUT121), .ZN(n744) );
  XOR2_X1 U794 ( .A(n782), .B(KEYINPUT88), .Z(n736) );
  NAND2_X1 U795 ( .A1(n736), .A2(n655), .ZN(n737) );
  NAND2_X1 U796 ( .A1(n738), .A2(n737), .ZN(n742) );
  NAND2_X1 U797 ( .A1(KEYINPUT88), .A2(n739), .ZN(n740) );
  NAND2_X1 U798 ( .A1(KEYINPUT2), .A2(n740), .ZN(n741) );
  NAND2_X1 U799 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U800 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U801 ( .A1(n745), .A2(G953), .ZN(n746) );
  XNOR2_X1 U802 ( .A(n746), .B(KEYINPUT53), .ZN(G75) );
  BUF_X2 U803 ( .A(n747), .Z(n756) );
  NAND2_X1 U804 ( .A1(n756), .A2(G469), .ZN(n751) );
  XOR2_X1 U805 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n748) );
  NOR2_X1 U806 ( .A1(n759), .A2(n752), .ZN(G54) );
  NAND2_X1 U807 ( .A1(G478), .A2(n756), .ZN(n753) );
  XNOR2_X1 U808 ( .A(n753), .B(n754), .ZN(n755) );
  NOR2_X1 U809 ( .A1(n759), .A2(n755), .ZN(G63) );
  NAND2_X1 U810 ( .A1(G217), .A2(n756), .ZN(n757) );
  XOR2_X1 U811 ( .A(G101), .B(n760), .Z(n761) );
  XNOR2_X1 U812 ( .A(KEYINPUT124), .B(n761), .ZN(n763) );
  NAND2_X1 U813 ( .A1(n763), .A2(n762), .ZN(n772) );
  NAND2_X1 U814 ( .A1(n655), .A2(n784), .ZN(n764) );
  XNOR2_X1 U815 ( .A(n764), .B(KEYINPUT123), .ZN(n770) );
  XOR2_X1 U816 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n766) );
  NAND2_X1 U817 ( .A1(G224), .A2(G953), .ZN(n765) );
  XNOR2_X1 U818 ( .A(n766), .B(n765), .ZN(n767) );
  NOR2_X1 U819 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U820 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U821 ( .A(n772), .B(n771), .ZN(G69) );
  XNOR2_X1 U822 ( .A(n774), .B(n773), .ZN(n775) );
  XNOR2_X1 U823 ( .A(n775), .B(KEYINPUT125), .ZN(n776) );
  XOR2_X1 U824 ( .A(n777), .B(n776), .Z(n781) );
  XOR2_X1 U825 ( .A(G227), .B(n781), .Z(n778) );
  NAND2_X1 U826 ( .A1(n778), .A2(G900), .ZN(n779) );
  XNOR2_X1 U827 ( .A(n779), .B(KEYINPUT126), .ZN(n780) );
  NAND2_X1 U828 ( .A1(n780), .A2(G953), .ZN(n786) );
  XOR2_X1 U829 ( .A(n782), .B(n781), .Z(n783) );
  NAND2_X1 U830 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U831 ( .A1(n786), .A2(n785), .ZN(G72) );
  XOR2_X1 U832 ( .A(n787), .B(G122), .Z(G24) );
  XOR2_X1 U833 ( .A(G119), .B(n788), .Z(n789) );
  XNOR2_X1 U834 ( .A(KEYINPUT127), .B(n789), .ZN(G21) );
  XOR2_X1 U835 ( .A(G140), .B(n790), .Z(G42) );
  XNOR2_X1 U836 ( .A(n791), .B(G131), .ZN(G33) );
  XNOR2_X1 U837 ( .A(n792), .B(G137), .ZN(G39) );
endmodule

